//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n931_, new_n932_, new_n933_, new_n934_, new_n936_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n962_, new_n963_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n975_, new_n976_, new_n977_, new_n979_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n987_, new_n988_;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(new_n216_), .A3(new_n213_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n203_), .A2(new_n204_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .A4(new_n206_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT29), .ZN(new_n222_));
  INV_X1    g021(.A(G204gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT83), .B1(new_n223_), .B2(G197gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT83), .ZN(new_n225_));
  INV_X1    g024(.A(G197gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(G204gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT21), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(G197gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n224_), .A2(new_n227_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n223_), .A2(G197gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n226_), .A2(G204gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT21), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n230_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n228_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n224_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G228gat), .A2(G233gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT82), .Z(new_n241_));
  AND3_X1   g040(.A1(new_n222_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n219_), .A2(new_n218_), .A3(new_n206_), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n214_), .A2(new_n211_), .B1(new_n243_), .B2(new_n217_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT84), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT84), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n221_), .A2(new_n247_), .A3(KEYINPUT29), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n235_), .A2(new_n238_), .A3(KEYINPUT85), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT85), .B1(new_n235_), .B2(new_n238_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n246_), .B(new_n248_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n241_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n242_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G78gat), .B(G106gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT86), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT87), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n259_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n246_), .A2(new_n248_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT85), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n239_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n235_), .A2(new_n238_), .A3(KEYINPUT85), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n241_), .B1(new_n261_), .B2(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(KEYINPUT87), .B(new_n254_), .C1(new_n266_), .C2(new_n242_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n253_), .A2(KEYINPUT86), .A3(new_n255_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n258_), .A2(new_n260_), .A3(new_n267_), .A4(new_n268_), .ZN(new_n269_));
  OR3_X1    g068(.A1(new_n221_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT28), .B1(new_n221_), .B2(KEYINPUT29), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G22gat), .B(G50gat), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n272_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n269_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT88), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT88), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n269_), .A2(new_n279_), .A3(new_n276_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n254_), .B1(new_n266_), .B2(new_n242_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(new_n275_), .A3(new_n256_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT89), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT89), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n281_), .A2(new_n284_), .A3(new_n275_), .A4(new_n256_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n278_), .A2(new_n280_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT96), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G226gat), .A2(G233gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT19), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n292_), .B(new_n293_), .C1(G183gat), .C2(G190gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT80), .ZN(new_n295_));
  INV_X1    g094(.A(G169gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT22), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(G176gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT22), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(KEYINPUT80), .A3(G169gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n297_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n294_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT26), .B(G190gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT78), .B1(new_n305_), .B2(G183gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT25), .B(G183gat), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n304_), .B(new_n306_), .C1(new_n307_), .C2(KEYINPUT78), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n290_), .B(new_n291_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT24), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n312_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT79), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n318_), .A2(KEYINPUT24), .A3(new_n302_), .A4(new_n313_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n303_), .B1(new_n311_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT20), .B1(new_n321_), .B2(new_n239_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n235_), .A2(new_n238_), .ZN(new_n323_));
  INV_X1    g122(.A(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT26), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT26), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G190gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT90), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n304_), .A2(KEYINPUT90), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(new_n331_), .A3(new_n307_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n332_), .A2(new_n319_), .A3(new_n316_), .A4(new_n310_), .ZN(new_n333_));
  XOR2_X1   g132(.A(KEYINPUT22), .B(G169gat), .Z(new_n334_));
  OAI211_X1 g133(.A(new_n294_), .B(new_n302_), .C1(G176gat), .C2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n323_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n289_), .B1(new_n322_), .B2(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G8gat), .B(G36gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n338_), .B(new_n339_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n341_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT20), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n321_), .B2(new_n239_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n289_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n323_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n337_), .A2(new_n347_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT27), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n346_), .A2(KEYINPUT95), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT95), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n342_), .A2(new_n356_), .A3(new_n345_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n263_), .A2(new_n335_), .A3(new_n333_), .A4(new_n264_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n349_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n289_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n322_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n333_), .A2(new_n335_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n239_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n350_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n358_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n287_), .B1(new_n354_), .B2(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n322_), .A2(new_n336_), .A3(new_n289_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n350_), .B1(new_n359_), .B2(new_n349_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n355_), .B(new_n357_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n370_), .A2(KEYINPUT96), .A3(KEYINPUT27), .A4(new_n353_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT27), .ZN(new_n372_));
  INV_X1    g171(.A(new_n353_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n347_), .B1(new_n337_), .B2(new_n352_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n367_), .A2(new_n371_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G227gat), .A2(G233gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(G15gat), .Z(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT30), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n321_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G127gat), .B(G134gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G113gat), .B(G120gat), .Z(new_n384_));
  AOI21_X1  g183(.A(new_n381_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G113gat), .B(G120gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n382_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n382_), .A2(new_n386_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n385_), .B1(new_n390_), .B2(new_n381_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n380_), .B(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G71gat), .B(G99gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G43gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT31), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n393_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n397_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT93), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n388_), .A2(new_n404_), .A3(new_n389_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n389_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT93), .B1(new_n406_), .B2(new_n387_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n407_), .A3(new_n244_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n381_), .B1(new_n406_), .B2(new_n387_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n385_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n221_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n403_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT4), .B1(new_n391_), .B2(new_n221_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n402_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n408_), .A2(new_n411_), .A3(new_n401_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G85gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT0), .B(G57gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n418_), .B(new_n419_), .Z(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n414_), .A2(new_n415_), .A3(new_n420_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n400_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n286_), .A2(new_n376_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n400_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n283_), .A2(new_n285_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n269_), .A2(new_n279_), .A3(new_n276_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n279_), .B1(new_n269_), .B2(new_n276_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n430_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n423_), .A2(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT33), .A4(new_n420_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n408_), .A2(new_n411_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT94), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n401_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(new_n438_), .B2(new_n437_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n401_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n421_), .A3(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n435_), .A2(new_n436_), .A3(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT92), .B1(new_n373_), .B2(new_n374_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n337_), .A2(new_n352_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n346_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT92), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(new_n353_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n347_), .A2(KEYINPUT32), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n445_), .A2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n451_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n429_), .B1(new_n433_), .B2(new_n456_), .ZN(new_n457_));
  AND4_X1   g256(.A1(new_n371_), .A2(new_n425_), .A3(new_n375_), .A4(new_n367_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n278_), .A2(new_n280_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n459_), .B2(new_n430_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n428_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT70), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G190gat), .B(G218gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G134gat), .B(G162gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n465_), .B(KEYINPUT36), .Z(new_n466_));
  INV_X1    g265(.A(G85gat), .ZN(new_n467_));
  INV_X1    g266(.A(G92gat), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n467_), .A2(new_n468_), .A3(KEYINPUT9), .ZN(new_n469_));
  AND2_X1   g268(.A1(G85gat), .A2(G92gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(G85gat), .A2(G92gat), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(KEYINPUT9), .B2(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n474_));
  INV_X1    g273(.A(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT65), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(G99gat), .A3(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT65), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n474_), .A2(new_n484_), .A3(new_n475_), .A4(new_n476_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n473_), .A2(new_n478_), .A3(new_n483_), .A4(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G85gat), .B(G92gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AOI211_X1 g290(.A(KEYINPUT8), .B(new_n487_), .C1(new_n491_), .C2(new_n483_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n494_));
  INV_X1    g293(.A(G99gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n475_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n481_), .B1(G99gat), .B2(G106gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n488_), .B(new_n496_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n493_), .B1(new_n499_), .B2(new_n472_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n486_), .B1(new_n492_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT67), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G29gat), .B(G36gat), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G43gat), .B(G50gat), .Z(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT15), .ZN(new_n511_));
  OAI211_X1 g310(.A(KEYINPUT67), .B(new_n486_), .C1(new_n492_), .C2(new_n500_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n503_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G232gat), .A2(G233gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT34), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT35), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n516_), .B(KEYINPUT69), .Z(new_n517_));
  NOR2_X1   g316(.A1(new_n515_), .A2(KEYINPUT35), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n499_), .A2(new_n472_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT8), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n499_), .A2(new_n493_), .A3(new_n472_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT9), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n487_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n483_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n469_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n478_), .A2(new_n485_), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n520_), .A2(new_n521_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n518_), .B1(new_n527_), .B2(new_n510_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n513_), .A2(new_n517_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n517_), .B1(new_n513_), .B2(new_n528_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n462_), .B(new_n466_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n513_), .A2(new_n528_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n517_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n513_), .A2(new_n517_), .A3(new_n528_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n465_), .A2(KEYINPUT36), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n531_), .A2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n466_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT70), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n461_), .A2(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n542_), .A2(KEYINPUT98), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(KEYINPUT98), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(G127gat), .B(G155gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT16), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G183gat), .B(G211gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G1gat), .B(G8gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT14), .ZN(new_n552_));
  INV_X1    g351(.A(G8gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT72), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT72), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(G8gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n552_), .B1(new_n557_), .B2(G1gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(G15gat), .B(G22gat), .Z(new_n559_));
  OAI21_X1  g358(.A(new_n551_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT72), .B(G8gat), .ZN(new_n561_));
  INV_X1    g360(.A(G1gat), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT14), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n559_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n564_), .A3(new_n550_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT73), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n566_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G57gat), .B(G64gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT11), .ZN(new_n571_));
  XOR2_X1   g370(.A(G71gat), .B(G78gat), .Z(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n570_), .A2(KEYINPUT11), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n571_), .A2(new_n572_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n569_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT74), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n549_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n549_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(KEYINPUT17), .B2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n580_), .A2(KEYINPUT17), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT66), .B1(new_n501_), .B2(new_n577_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n501_), .A2(new_n577_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n520_), .A2(new_n521_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT66), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n571_), .A2(new_n572_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n587_), .A2(new_n588_), .A3(new_n486_), .A4(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n585_), .A2(new_n586_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT64), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n589_), .B(KEYINPUT12), .C1(new_n574_), .C2(new_n573_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n503_), .A2(new_n512_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT12), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n599_), .B1(new_n527_), .B2(new_n590_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n594_), .B1(new_n527_), .B2(new_n590_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G120gat), .B(G148gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT5), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G176gat), .B(G204gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n595_), .A2(new_n602_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT68), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n595_), .A2(new_n602_), .A3(KEYINPUT68), .A4(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n595_), .A2(new_n602_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n606_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(KEYINPUT13), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT13), .B1(new_n611_), .B2(new_n614_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G113gat), .B(G141gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G169gat), .B(G197gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n620_), .B(new_n621_), .Z(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n510_), .B(KEYINPUT15), .Z(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n566_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n507_), .A2(KEYINPUT75), .A3(new_n509_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT75), .B1(new_n507_), .B2(new_n509_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n566_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G229gat), .A2(G233gat), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n625_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT75), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n510_), .A2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n634_), .A2(new_n560_), .A3(new_n565_), .A4(new_n626_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n629_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n630_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT76), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(KEYINPUT76), .A3(new_n637_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n632_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT77), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n623_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT76), .B1(new_n636_), .B2(new_n637_), .ZN(new_n645_));
  AOI211_X1 g444(.A(new_n639_), .B(new_n630_), .C1(new_n629_), .C2(new_n635_), .ZN(new_n646_));
  OAI22_X1  g445(.A1(new_n645_), .A2(new_n646_), .B1(new_n625_), .B2(new_n631_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(KEYINPUT77), .A3(new_n622_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n644_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n619_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n545_), .A2(new_n584_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n424_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G1gat), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT38), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n376_), .B(new_n430_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n426_), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n443_), .A2(new_n449_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n400_), .B1(new_n286_), .B2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n376_), .A2(new_n425_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n433_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n657_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n651_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n584_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT71), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n539_), .A2(new_n537_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(KEYINPUT37), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT37), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n540_), .A2(new_n668_), .A3(new_n537_), .A4(new_n531_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n538_), .A2(new_n665_), .A3(new_n668_), .A4(new_n540_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n664_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n663_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT97), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT97), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n663_), .A2(new_n676_), .A3(new_n673_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n675_), .A2(new_n562_), .A3(new_n424_), .A4(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n655_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n679_), .A2(KEYINPUT99), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(KEYINPUT99), .ZN(new_n681_));
  OAI221_X1 g480(.A(new_n654_), .B1(new_n655_), .B2(new_n678_), .C1(new_n680_), .C2(new_n681_), .ZN(G1324gat));
  XNOR2_X1  g481(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n683_));
  INV_X1    g482(.A(new_n376_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n651_), .A2(new_n584_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n684_), .B(new_n685_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT39), .B1(new_n686_), .B2(G8gat), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n376_), .A2(new_n557_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n675_), .A2(new_n677_), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT100), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n675_), .A2(new_n694_), .A3(new_n677_), .A4(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n683_), .B1(new_n690_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n689_), .ZN(new_n698_));
  AND4_X1   g497(.A1(new_n696_), .A2(new_n687_), .A3(new_n698_), .A4(new_n683_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1325gat));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n400_), .B(new_n685_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G15gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n703_), .A2(new_n705_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n701_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n708_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(KEYINPUT103), .A3(new_n706_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n674_), .A2(G15gat), .A3(new_n429_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT104), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n711_), .A3(new_n713_), .ZN(G1326gat));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n652_), .A2(new_n433_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(G22gat), .ZN(new_n717_));
  INV_X1    g516(.A(G22gat), .ZN(new_n718_));
  AOI211_X1 g517(.A(KEYINPUT42), .B(new_n718_), .C1(new_n652_), .C2(new_n433_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n433_), .A2(new_n718_), .ZN(new_n720_));
  OAI22_X1  g519(.A1(new_n717_), .A2(new_n719_), .B1(new_n674_), .B2(new_n720_), .ZN(G1327gat));
  NOR2_X1   g520(.A1(new_n664_), .A2(new_n541_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n663_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G29gat), .B1(new_n724_), .B2(new_n424_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n651_), .A2(new_n664_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n670_), .A2(new_n671_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n459_), .A2(new_n430_), .A3(new_n658_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n661_), .A2(new_n729_), .A3(new_n429_), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT43), .B(new_n728_), .C1(new_n730_), .C2(new_n428_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n461_), .B2(new_n727_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n726_), .B1(new_n731_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n726_), .B(KEYINPUT44), .C1(new_n731_), .C2(new_n733_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n424_), .A2(G29gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n725_), .B1(new_n738_), .B2(new_n739_), .ZN(G1328gat));
  NOR2_X1   g539(.A1(new_n376_), .A2(G36gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n663_), .A2(new_n722_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n736_), .A2(new_n737_), .A3(new_n684_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(G36gat), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT46), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(KEYINPUT105), .A3(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n747_), .A2(KEYINPUT105), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n747_), .A2(KEYINPUT105), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n746_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1329gat));
  NAND4_X1  g551(.A1(new_n736_), .A2(new_n737_), .A3(G43gat), .A4(new_n400_), .ZN(new_n753_));
  XOR2_X1   g552(.A(KEYINPUT106), .B(G43gat), .Z(new_n754_));
  OAI21_X1  g553(.A(new_n754_), .B1(new_n723_), .B2(new_n429_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  XOR2_X1   g555(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n757_));
  XNOR2_X1  g556(.A(new_n756_), .B(new_n757_), .ZN(G1330gat));
  AOI21_X1  g557(.A(G50gat), .B1(new_n724_), .B2(new_n433_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n433_), .A2(G50gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n738_), .B2(new_n760_), .ZN(G1331gat));
  INV_X1    g560(.A(new_n649_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n618_), .A2(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n461_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n673_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT108), .ZN(new_n766_));
  INV_X1    g565(.A(G57gat), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(new_n424_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n763_), .A2(new_n664_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n545_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n767_), .B1(new_n770_), .B2(new_n424_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n772_));
  OR3_X1    g571(.A1(new_n768_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n768_), .B2(new_n771_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1332gat));
  INV_X1    g574(.A(G64gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n766_), .A2(new_n776_), .A3(new_n684_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n770_), .A2(new_n684_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G64gat), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(KEYINPUT48), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(KEYINPUT48), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(G1333gat));
  INV_X1    g581(.A(G71gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n766_), .A2(new_n783_), .A3(new_n400_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n770_), .A2(new_n400_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(G71gat), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(KEYINPUT49), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(KEYINPUT49), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(G1334gat));
  INV_X1    g588(.A(G78gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n766_), .A2(new_n790_), .A3(new_n433_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n769_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n433_), .B(new_n792_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n793_), .A2(new_n794_), .A3(G78gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n793_), .B2(G78gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n791_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n797_), .B(new_n798_), .ZN(G1335gat));
  NAND2_X1  g598(.A1(new_n763_), .A2(new_n584_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT43), .B1(new_n662_), .B2(new_n728_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n461_), .A2(new_n732_), .A3(new_n727_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n800_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(G85gat), .B1(new_n804_), .B2(new_n425_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n764_), .A2(new_n722_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n467_), .A3(new_n424_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1336gat));
  OAI21_X1  g607(.A(G92gat), .B1(new_n804_), .B2(new_n376_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(new_n468_), .A3(new_n684_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(G1337gat));
  OAI21_X1  g610(.A(G99gat), .B1(new_n804_), .B2(new_n429_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n806_), .A2(new_n474_), .A3(new_n476_), .A4(new_n400_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(KEYINPUT111), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n814_), .B(new_n816_), .ZN(G1338gat));
  INV_X1    g616(.A(new_n800_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n433_), .B(new_n818_), .C1(new_n731_), .C2(new_n733_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n820_));
  OAI21_X1  g619(.A(G106gat), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT112), .B1(new_n803_), .B2(new_n433_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT52), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n803_), .A2(KEYINPUT112), .A3(new_n433_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n820_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .A4(G106gat), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n823_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n806_), .A2(new_n475_), .A3(new_n433_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT53), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n832_), .A3(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1339gat));
  XNOR2_X1  g633(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n629_), .B(new_n637_), .C1(new_n624_), .C2(new_n566_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n636_), .A2(new_n630_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n622_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n647_), .B2(new_n622_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n611_), .B2(new_n614_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n598_), .A2(new_n585_), .A3(new_n591_), .A4(new_n600_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n594_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n598_), .A2(KEYINPUT55), .A3(new_n600_), .A4(new_n601_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n602_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(new_n844_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n613_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(KEYINPUT56), .A3(new_n613_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n611_), .A2(new_n648_), .A3(new_n644_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n841_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n541_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n836_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n611_), .A2(new_n644_), .A3(new_n648_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT57), .B(new_n541_), .C1(new_n858_), .C2(new_n841_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n840_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n847_), .A2(KEYINPUT56), .A3(new_n613_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT56), .B1(new_n847_), .B2(new_n613_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(KEYINPUT58), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  OAI221_X1 g665(.A(new_n860_), .B1(new_n864_), .B2(KEYINPUT58), .C1(new_n861_), .C2(new_n862_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n727_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n856_), .A2(new_n859_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n584_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n617_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n615_), .A3(new_n649_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n873_), .A2(KEYINPUT113), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(KEYINPUT113), .ZN(new_n875_));
  OAI22_X1  g674(.A1(new_n672_), .A2(new_n872_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n616_), .A2(new_n762_), .A3(new_n617_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n875_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n728_), .A2(new_n877_), .A3(new_n664_), .A4(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n870_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n656_), .A2(new_n425_), .A3(new_n429_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n869_), .A2(new_n584_), .B1(new_n876_), .B2(new_n879_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n883_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT116), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n884_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G113gat), .B1(new_n888_), .B2(new_n762_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n881_), .A2(new_n883_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT59), .ZN(new_n891_));
  INV_X1    g690(.A(new_n859_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n856_), .A2(new_n868_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n856_), .A2(KEYINPUT117), .A3(new_n868_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n664_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n880_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n886_), .A2(KEYINPUT59), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n891_), .B1(new_n899_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n762_), .A2(G113gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(KEYINPUT118), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n889_), .B1(new_n903_), .B2(new_n905_), .ZN(G1340gat));
  XNOR2_X1  g705(.A(KEYINPUT119), .B(G120gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n907_), .B1(new_n618_), .B2(KEYINPUT60), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n888_), .B(new_n908_), .C1(KEYINPUT60), .C2(new_n907_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n619_), .B(new_n891_), .C1(new_n899_), .C2(new_n901_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n907_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n909_), .B1(new_n912_), .B2(new_n914_), .ZN(G1341gat));
  OAI21_X1  g714(.A(G127gat), .B1(new_n902_), .B2(new_n584_), .ZN(new_n916_));
  INV_X1    g715(.A(G127gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n888_), .A2(new_n917_), .A3(new_n664_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(G1342gat));
  INV_X1    g718(.A(G134gat), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n728_), .A2(new_n920_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n891_), .B(new_n921_), .C1(new_n899_), .C2(new_n901_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n884_), .A2(new_n887_), .A3(new_n855_), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n923_), .A2(KEYINPUT121), .A3(new_n920_), .ZN(new_n924_));
  AOI21_X1  g723(.A(KEYINPUT121), .B1(new_n923_), .B2(new_n920_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n922_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT122), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n928_), .B(new_n922_), .C1(new_n924_), .C2(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1343gat));
  NOR2_X1   g729(.A1(new_n885_), .A2(new_n400_), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n931_), .A2(new_n376_), .A3(new_n433_), .A4(new_n424_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n649_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(KEYINPUT123), .B(G141gat), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(G1344gat));
  NOR2_X1   g734(.A1(new_n932_), .A2(new_n618_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(new_n204_), .ZN(G1345gat));
  NOR2_X1   g736(.A1(new_n932_), .A2(new_n584_), .ZN(new_n938_));
  XOR2_X1   g737(.A(KEYINPUT61), .B(G155gat), .Z(new_n939_));
  XNOR2_X1  g738(.A(new_n938_), .B(new_n939_), .ZN(G1346gat));
  OAI21_X1  g739(.A(G162gat), .B1(new_n932_), .B2(new_n728_), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n541_), .A2(G162gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n932_), .B2(new_n942_), .ZN(G1347gat));
  NOR2_X1   g742(.A1(new_n376_), .A2(new_n424_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n400_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n433_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n946_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n947_));
  OAI21_X1  g746(.A(G169gat), .B1(new_n947_), .B2(new_n649_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n949_));
  OR2_X1    g748(.A1(new_n948_), .A2(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n948_), .A2(new_n949_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n947_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n762_), .ZN(new_n953_));
  OAI211_X1 g752(.A(new_n950_), .B(new_n951_), .C1(new_n334_), .C2(new_n953_), .ZN(G1348gat));
  AOI21_X1  g753(.A(G176gat), .B1(new_n952_), .B2(new_n619_), .ZN(new_n955_));
  AOI21_X1  g754(.A(KEYINPUT124), .B1(new_n881_), .B2(new_n286_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n885_), .A2(new_n957_), .A3(new_n433_), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n956_), .A2(new_n958_), .A3(new_n945_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n618_), .A2(new_n298_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n955_), .B1(new_n959_), .B2(new_n960_), .ZN(G1349gat));
  AOI21_X1  g760(.A(G183gat), .B1(new_n959_), .B2(new_n664_), .ZN(new_n962_));
  NOR3_X1   g761(.A1(new_n947_), .A2(new_n584_), .A3(new_n307_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n962_), .A2(new_n963_), .ZN(G1350gat));
  NAND4_X1  g763(.A1(new_n952_), .A2(new_n855_), .A3(new_n330_), .A4(new_n331_), .ZN(new_n965_));
  OAI211_X1 g764(.A(new_n727_), .B(new_n946_), .C1(new_n897_), .C2(new_n898_), .ZN(new_n966_));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n967_));
  AND3_X1   g766(.A1(new_n966_), .A2(new_n967_), .A3(G190gat), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n967_), .B1(new_n966_), .B2(G190gat), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n965_), .B1(new_n968_), .B2(new_n969_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n970_), .A2(KEYINPUT126), .ZN(new_n971_));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n972_));
  OAI211_X1 g771(.A(new_n965_), .B(new_n972_), .C1(new_n968_), .C2(new_n969_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n971_), .A2(new_n973_), .ZN(G1351gat));
  AND2_X1   g773(.A1(new_n433_), .A2(new_n944_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n931_), .A2(new_n975_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n976_), .A2(new_n649_), .ZN(new_n977_));
  XNOR2_X1  g776(.A(new_n977_), .B(new_n226_), .ZN(G1352gat));
  NOR2_X1   g777(.A1(new_n976_), .A2(new_n618_), .ZN(new_n979_));
  XNOR2_X1  g778(.A(new_n979_), .B(new_n223_), .ZN(G1353gat));
  INV_X1    g779(.A(new_n976_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n584_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n982_));
  XNOR2_X1  g781(.A(new_n982_), .B(KEYINPUT127), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n981_), .A2(new_n983_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n985_));
  XOR2_X1   g784(.A(new_n984_), .B(new_n985_), .Z(G1354gat));
  OR3_X1    g785(.A1(new_n976_), .A2(G218gat), .A3(new_n541_), .ZN(new_n987_));
  OAI21_X1  g786(.A(G218gat), .B1(new_n976_), .B2(new_n728_), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n987_), .A2(new_n988_), .ZN(G1355gat));
endmodule


