//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_;
  NOR2_X1   g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n205_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(G169gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT76), .ZN(new_n210_));
  INV_X1    g009(.A(G190gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n210_), .B1(new_n211_), .B2(KEYINPUT26), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(KEYINPUT26), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(KEYINPUT75), .A2(G183gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT25), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT26), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(KEYINPUT76), .A3(G190gat), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n214_), .A2(new_n217_), .A3(new_n218_), .A4(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n215_), .B(KEYINPUT25), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n212_), .A2(new_n220_), .A3(new_n213_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT77), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n204_), .A2(KEYINPUT23), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n203_), .A2(G183gat), .A3(G190gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229_));
  INV_X1    g028(.A(G169gat), .ZN(new_n230_));
  INV_X1    g029(.A(G176gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT78), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n228_), .A2(KEYINPUT78), .A3(new_n232_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n209_), .B1(new_n225_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT30), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G71gat), .B(G99gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n244_), .B(KEYINPUT31), .Z(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT80), .B(G15gat), .Z(new_n246_));
  NAND2_X1  g045(.A1(G227gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT79), .B(G43gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  XOR2_X1   g049(.A(G113gat), .B(G120gat), .Z(new_n251_));
  INV_X1    g050(.A(G134gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G127gat), .ZN(new_n253_));
  INV_X1    g052(.A(G127gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G134gat), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n253_), .A2(new_n255_), .A3(KEYINPUT81), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT81), .B1(new_n253_), .B2(new_n255_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n251_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT81), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n254_), .A2(G134gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n252_), .A2(G127gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n253_), .A2(new_n255_), .A3(KEYINPUT81), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G113gat), .B(G120gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n258_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n250_), .B(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n245_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n245_), .A2(new_n269_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G155gat), .B(G162gat), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT83), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n278_));
  NOR2_X1   g077(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n274_), .B(new_n276_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT2), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n285_), .B1(new_n286_), .B2(new_n276_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT84), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n288_), .A2(KEYINPUT84), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n287_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n273_), .B1(new_n282_), .B2(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n273_), .A2(KEYINPUT1), .ZN(new_n293_));
  INV_X1    g092(.A(new_n276_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n283_), .A3(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  OAI211_X1 g096(.A(KEYINPUT99), .B(new_n267_), .C1(new_n292_), .C2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT99), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n276_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT83), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n288_), .B(KEYINPUT84), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n294_), .A2(KEYINPUT3), .B1(new_n284_), .B2(new_n283_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .A4(new_n280_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n273_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n297_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n299_), .B1(new_n306_), .B2(new_n266_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n298_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT100), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n258_), .A2(new_n265_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n309_), .B1(new_n258_), .B2(new_n265_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n306_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT101), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT101), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n306_), .B(new_n316_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n308_), .A2(new_n314_), .A3(new_n315_), .A4(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT102), .ZN(new_n319_));
  INV_X1    g118(.A(new_n317_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n256_), .A2(new_n257_), .A3(new_n251_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n264_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT100), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n310_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n316_), .B1(new_n324_), .B2(new_n306_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT102), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n315_), .A4(new_n308_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n304_), .A2(new_n305_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n297_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT4), .B1(new_n331_), .B2(new_n267_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n308_), .A2(new_n314_), .A3(new_n317_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n332_), .B1(new_n333_), .B2(KEYINPUT4), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n319_), .B(new_n328_), .C1(new_n334_), .C2(new_n315_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G1gat), .B(G29gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G85gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n335_), .A2(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n328_), .A2(new_n319_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n315_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n326_), .B2(new_n308_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n343_), .B1(new_n345_), .B2(new_n332_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n342_), .A2(new_n346_), .A3(new_n339_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n341_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n272_), .A2(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n331_), .A2(KEYINPUT29), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT28), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT85), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n331_), .A2(KEYINPUT29), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT28), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n352_), .A2(new_n353_), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n353_), .B1(new_n352_), .B2(new_n356_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G22gat), .B(G50gat), .Z(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  OR3_X1    g159(.A1(new_n357_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n360_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G197gat), .A2(G204gat), .ZN(new_n363_));
  INV_X1    g162(.A(G197gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT87), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT87), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(G197gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n363_), .B1(new_n368_), .B2(G204gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G211gat), .B(G218gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(KEYINPUT21), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n363_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT87), .B(G197gat), .ZN(new_n374_));
  INV_X1    g173(.A(G204gat), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n373_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(KEYINPUT89), .B(KEYINPUT21), .Z(new_n377_));
  AOI21_X1  g176(.A(new_n371_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT88), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n364_), .B2(G204gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n380_), .B1(new_n374_), .B2(G204gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n366_), .A2(G197gat), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n364_), .A2(KEYINPUT87), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n379_), .B(new_n375_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(KEYINPUT21), .A3(new_n384_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n378_), .A2(KEYINPUT90), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT90), .B1(new_n378_), .B2(new_n385_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n372_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n331_), .A2(KEYINPUT29), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G228gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT86), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT91), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n388_), .B(new_n389_), .C1(KEYINPUT91), .C2(new_n392_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G78gat), .B(G106gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n361_), .A2(new_n362_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(KEYINPUT93), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT93), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n399_), .B1(new_n396_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT94), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n402_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n401_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n361_), .A2(new_n362_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT92), .B1(new_n397_), .B2(new_n399_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n400_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n397_), .A2(KEYINPUT92), .A3(new_n399_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n409_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n408_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G226gat), .A2(G233gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT19), .ZN(new_n417_));
  INV_X1    g216(.A(new_n372_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT90), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n381_), .A2(KEYINPUT21), .A3(new_n384_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n377_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n370_), .B1(new_n369_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n419_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n378_), .A2(KEYINPUT90), .A3(new_n385_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n418_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT26), .B(G190gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT25), .B(G183gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n239_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n429_), .A2(KEYINPUT95), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n233_), .B1(new_n429_), .B2(KEYINPUT95), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n228_), .B(KEYINPUT96), .C1(G183gat), .C2(G190gat), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n432_), .A2(new_n208_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT96), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n206_), .A2(new_n434_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n430_), .A2(new_n431_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT20), .B1(new_n425_), .B2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n388_), .A2(new_n241_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n417_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G8gat), .B(G36gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT18), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G64gat), .B(G92gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n441_), .B(new_n442_), .Z(new_n443_));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n444_), .B1(new_n425_), .B2(new_n436_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n417_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n388_), .A2(new_n241_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n439_), .A2(new_n443_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT105), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n447_), .B1(new_n445_), .B2(new_n450_), .ZN(new_n451_));
  AOI211_X1 g250(.A(KEYINPUT105), .B(new_n444_), .C1(new_n425_), .C2(new_n436_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n417_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n388_), .A2(new_n241_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n430_), .A2(new_n431_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n433_), .A2(new_n435_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n444_), .B1(new_n388_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(new_n446_), .A3(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n453_), .A2(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(KEYINPUT27), .B(new_n449_), .C1(new_n460_), .C2(new_n443_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT97), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n449_), .A2(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n439_), .A2(new_n448_), .A3(KEYINPUT97), .A4(new_n443_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n443_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n448_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n446_), .B1(new_n454_), .B2(new_n458_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n465_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n463_), .A2(new_n464_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT27), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n461_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n415_), .A2(KEYINPUT107), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT107), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n461_), .A2(new_n471_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n474_), .B1(new_n414_), .B2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n350_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n443_), .A2(KEYINPUT32), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n478_), .B1(new_n453_), .B2(new_n459_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n466_), .A2(new_n467_), .ZN(new_n480_));
  AOI221_X4 g279(.A(new_n479_), .B1(new_n478_), .B2(new_n480_), .C1(new_n347_), .C2(new_n341_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n342_), .A2(new_n346_), .A3(KEYINPUT33), .A4(new_n339_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n340_), .B1(new_n333_), .B2(new_n315_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT104), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT104), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n485_), .B(new_n340_), .C1(new_n333_), .C2(new_n315_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n484_), .B(new_n486_), .C1(new_n343_), .C2(new_n334_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n482_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n489_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT103), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT103), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n492_), .B(new_n489_), .C1(new_n335_), .C2(new_n340_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n488_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n443_), .B1(new_n439_), .B2(new_n448_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n462_), .B2(new_n449_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT98), .B1(new_n496_), .B2(new_n464_), .ZN(new_n497_));
  AND4_X1   g296(.A1(KEYINPUT98), .A2(new_n463_), .A3(new_n464_), .A4(new_n468_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n481_), .B1(new_n494_), .B2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT106), .B1(new_n500_), .B2(new_n414_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n480_), .A2(new_n478_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n348_), .B(new_n502_), .C1(new_n460_), .C2(new_n478_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n482_), .A2(new_n487_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n493_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n492_), .B1(new_n347_), .B2(new_n489_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT98), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n469_), .B(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n503_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT106), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(new_n415_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n414_), .A2(new_n472_), .A3(new_n349_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n501_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n272_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n477_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT72), .B(G1gat), .Z(new_n518_));
  INV_X1    g317(.A(G8gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT14), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G1gat), .B(G8gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G29gat), .B(G36gat), .Z(new_n525_));
  XOR2_X1   g324(.A(G43gat), .B(G50gat), .Z(new_n526_));
  XOR2_X1   g325(.A(new_n525_), .B(new_n526_), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n524_), .B(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(G229gat), .A3(G233gat), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n527_), .B(KEYINPUT15), .Z(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n524_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n524_), .A2(new_n527_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT73), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n531_), .A2(new_n532_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n529_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G169gat), .B(G197gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n536_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT74), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n541_), .A2(KEYINPUT74), .A3(new_n543_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n517_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(KEYINPUT70), .A2(KEYINPUT37), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT71), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(G85gat), .B(G92gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT66), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT7), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n558_), .A2(new_n559_), .ZN(new_n561_));
  INV_X1    g360(.A(G99gat), .ZN(new_n562_));
  INV_X1    g361(.A(G106gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n560_), .B1(new_n561_), .B2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n565_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n554_), .B1(new_n557_), .B2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT8), .ZN(new_n568_));
  INV_X1    g367(.A(G85gat), .ZN(new_n569_));
  INV_X1    g368(.A(G92gat), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n569_), .A2(new_n570_), .A3(KEYINPUT9), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n571_), .B1(new_n554_), .B2(KEYINPUT9), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT10), .B(G99gat), .Z(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT64), .B(G106gat), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n572_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(new_n557_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n568_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n530_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT34), .ZN(new_n582_));
  OAI221_X1 g381(.A(new_n580_), .B1(KEYINPUT35), .B2(new_n582_), .C1(new_n527_), .C2(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(KEYINPUT35), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n585_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n585_), .A2(new_n589_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(KEYINPUT70), .A2(KEYINPUT37), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n553_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  OAI221_X1 g394(.A(new_n552_), .B1(KEYINPUT70), .B2(KEYINPUT37), .C1(new_n591_), .C2(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G57gat), .B(G64gat), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT11), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT67), .ZN(new_n600_));
  XOR2_X1   g399(.A(G71gat), .B(G78gat), .Z(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(KEYINPUT11), .B2(new_n598_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n602_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n605_), .B(new_n606_), .Z(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(new_n524_), .Z(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT16), .ZN(new_n611_));
  XOR2_X1   g410(.A(G183gat), .B(G211gat), .Z(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT17), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n613_), .A2(KEYINPUT68), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n609_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n613_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n615_), .B1(KEYINPUT17), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n608_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n597_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT12), .ZN(new_n624_));
  INV_X1    g423(.A(new_n605_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(KEYINPUT68), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n605_), .B1(new_n568_), .B2(new_n578_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n626_), .B1(new_n627_), .B2(KEYINPUT68), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n568_), .A2(new_n605_), .A3(new_n578_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n579_), .A2(new_n625_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n624_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT69), .B1(new_n632_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n629_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n634_), .B1(new_n636_), .B2(new_n627_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n624_), .B2(new_n630_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT69), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n633_), .A4(new_n628_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n635_), .A2(new_n637_), .A3(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT5), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n643_), .B(new_n644_), .Z(new_n645_));
  NAND2_X1  g444(.A1(new_n641_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n645_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n635_), .A2(new_n637_), .A3(new_n640_), .A4(new_n647_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n646_), .A2(KEYINPUT13), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT13), .B1(new_n646_), .B2(new_n648_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n623_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n550_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n348_), .A3(new_n518_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT38), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n517_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n593_), .B(KEYINPUT108), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n652_), .A2(new_n549_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n659_), .A2(new_n620_), .A3(new_n661_), .A4(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G1gat), .B1(new_n663_), .B2(new_n349_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n656_), .A2(new_n657_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n658_), .A2(new_n664_), .A3(new_n665_), .ZN(G1324gat));
  NAND3_X1  g465(.A1(new_n655_), .A2(new_n519_), .A3(new_n475_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n663_), .A2(new_n472_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n668_), .A2(new_n669_), .A3(G8gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n668_), .B2(G8gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n667_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g472(.A(G15gat), .B1(new_n663_), .B2(new_n516_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT41), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n654_), .A2(G15gat), .A3(new_n516_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1326gat));
  OAI21_X1  g476(.A(G22gat), .B1(new_n663_), .B2(new_n415_), .ZN(new_n678_));
  XOR2_X1   g477(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n415_), .A2(G22gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n654_), .B2(new_n681_), .ZN(G1327gat));
  INV_X1    g481(.A(G29gat), .ZN(new_n683_));
  INV_X1    g482(.A(new_n597_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n517_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n491_), .A2(new_n493_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n499_), .A2(new_n687_), .A3(new_n504_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n414_), .B1(new_n688_), .B2(new_n503_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n513_), .B1(new_n689_), .B2(new_n511_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n272_), .B1(new_n690_), .B2(new_n501_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n686_), .B(new_n597_), .C1(new_n691_), .C2(new_n477_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n685_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n662_), .A2(new_n621_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT44), .B1(new_n693_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  AOI211_X1 g496(.A(new_n697_), .B(new_n694_), .C1(new_n685_), .C2(new_n692_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n683_), .B1(new_n699_), .B2(new_n348_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n593_), .A2(new_n621_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n652_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n550_), .A2(new_n703_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n704_), .A2(G29gat), .A3(new_n349_), .ZN(new_n705_));
  OR3_X1    g504(.A1(new_n700_), .A2(new_n701_), .A3(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n701_), .B1(new_n700_), .B2(new_n705_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1328gat));
  NOR3_X1   g507(.A1(new_n704_), .A2(G36gat), .A3(new_n472_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT45), .Z(new_n710_));
  NAND2_X1  g509(.A1(new_n693_), .A2(new_n695_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n697_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n693_), .A2(KEYINPUT44), .A3(new_n695_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n712_), .A2(KEYINPUT111), .A3(new_n475_), .A4(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G36gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT111), .B1(new_n699_), .B2(new_n475_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n710_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT46), .B(new_n710_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  NAND3_X1  g520(.A1(new_n699_), .A2(G43gat), .A3(new_n272_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n704_), .A2(new_n516_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(G43gat), .B2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(G1330gat));
  INV_X1    g525(.A(new_n704_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G50gat), .B1(new_n727_), .B2(new_n414_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n414_), .A2(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n699_), .B2(new_n729_), .ZN(G1331gat));
  NOR4_X1   g529(.A1(new_n517_), .A2(new_n623_), .A3(new_n548_), .A4(new_n651_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G57gat), .B1(new_n731_), .B2(new_n348_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n652_), .A2(new_n549_), .A3(new_n620_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n517_), .A2(new_n660_), .A3(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n349_), .A2(KEYINPUT113), .ZN(new_n735_));
  MUX2_X1   g534(.A(KEYINPUT113), .B(new_n735_), .S(G57gat), .Z(new_n736_));
  AOI21_X1  g535(.A(new_n732_), .B1(new_n734_), .B2(new_n736_), .ZN(G1332gat));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n475_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G64gat), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT48), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n472_), .A2(G64gat), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT114), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n731_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n743_), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n734_), .B2(new_n272_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT49), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n731_), .A2(new_n745_), .A3(new_n272_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1334gat));
  INV_X1    g548(.A(G78gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n734_), .B2(new_n414_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT50), .Z(new_n752_));
  NAND3_X1  g551(.A1(new_n731_), .A2(new_n750_), .A3(new_n414_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1335gat));
  NAND3_X1  g553(.A1(new_n652_), .A2(new_n549_), .A3(new_n621_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n685_), .B2(new_n692_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n349_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n517_), .A2(new_n548_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n651_), .A2(new_n702_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n569_), .A3(new_n348_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n758_), .A2(new_n763_), .ZN(G1336gat));
  OAI21_X1  g563(.A(G92gat), .B1(new_n757_), .B2(new_n472_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(new_n570_), .A3(new_n475_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1337gat));
  AOI21_X1  g566(.A(new_n562_), .B1(new_n756_), .B2(new_n272_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n761_), .A2(new_n516_), .A3(new_n574_), .ZN(new_n769_));
  OAI22_X1  g568(.A1(new_n768_), .A2(new_n769_), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n770_));
  NAND2_X1  g569(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n762_), .A2(new_n414_), .A3(new_n575_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n756_), .A2(new_n414_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(G106gat), .ZN(new_n776_));
  AOI211_X1 g575(.A(KEYINPUT52), .B(new_n563_), .C1(new_n756_), .C2(new_n414_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI211_X1 g578(.A(new_n349_), .B(new_n516_), .C1(new_n473_), .C2(new_n476_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n781_), .A2(KEYINPUT59), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n548_), .A2(new_n648_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n635_), .A2(new_n784_), .A3(new_n640_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n633_), .B1(new_n638_), .B2(new_n628_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n632_), .A2(new_n634_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(KEYINPUT55), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT56), .B1(new_n789_), .B2(new_n645_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  AOI211_X1 g590(.A(new_n791_), .B(new_n647_), .C1(new_n785_), .C2(new_n788_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n783_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n646_), .A2(new_n648_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n534_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n531_), .A2(new_n532_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n540_), .B1(new_n528_), .B2(new_n534_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n537_), .A2(new_n540_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n794_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n593_), .B1(new_n793_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT57), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n648_), .A2(new_n798_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT58), .B(new_n803_), .C1(new_n790_), .C2(new_n792_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n597_), .A3(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(KEYINPUT57), .B2(new_n800_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n802_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n800_), .A2(KEYINPUT57), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(KEYINPUT117), .A3(new_n808_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n620_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n622_), .A2(new_n549_), .A3(new_n651_), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(KEYINPUT54), .Z(new_n816_));
  OAI21_X1  g615(.A(new_n782_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n809_), .B2(new_n802_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n812_), .A2(KEYINPUT116), .A3(new_n808_), .A4(new_n801_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n621_), .A3(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n815_), .B(KEYINPUT54), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n781_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n817_), .B(new_n548_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G113gat), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n821_), .A2(new_n822_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n780_), .ZN(new_n828_));
  OR3_X1    g627(.A1(new_n828_), .A2(G113gat), .A3(new_n549_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n826_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT118), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n826_), .A2(new_n829_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1340gat));
  INV_X1    g633(.A(G120gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n651_), .B2(KEYINPUT60), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n823_), .B(new_n836_), .C1(KEYINPUT60), .C2(new_n835_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n811_), .A2(new_n813_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n621_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n822_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n828_), .A2(KEYINPUT59), .B1(new_n840_), .B2(new_n782_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n652_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n837_), .B1(new_n843_), .B2(new_n835_), .ZN(G1341gat));
  OAI21_X1  g643(.A(new_n254_), .B1(new_n828_), .B2(new_n621_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n845_), .A2(KEYINPUT119), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(KEYINPUT119), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n621_), .A2(new_n254_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n846_), .A2(new_n847_), .B1(new_n841_), .B2(new_n848_), .ZN(G1342gat));
  AOI21_X1  g648(.A(G134gat), .B1(new_n823_), .B2(new_n660_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n597_), .A2(G134gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT120), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n841_), .B2(new_n852_), .ZN(G1343gat));
  NAND4_X1  g652(.A1(new_n516_), .A2(new_n414_), .A3(new_n348_), .A4(new_n472_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT121), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n827_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n548_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n652_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g659(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n856_), .A2(new_n620_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n827_), .A2(new_n855_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n621_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n864_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n862_), .B1(new_n865_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n863_), .A2(new_n864_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n867_), .A2(new_n868_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n861_), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(G1346gat));
  OR3_X1    g673(.A1(new_n866_), .A2(G162gat), .A3(new_n661_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G162gat), .B1(new_n866_), .B2(new_n684_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n350_), .A2(new_n472_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n414_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n839_), .B2(new_n822_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n548_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  AND4_X1   g683(.A1(KEYINPUT124), .A2(new_n883_), .A3(new_n884_), .A4(G169gat), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n230_), .B1(new_n886_), .B2(KEYINPUT62), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n883_), .A2(new_n887_), .B1(KEYINPUT124), .B2(new_n884_), .ZN(new_n888_));
  XOR2_X1   g687(.A(KEYINPUT22), .B(G169gat), .Z(new_n889_));
  OAI22_X1  g688(.A1(new_n885_), .A2(new_n888_), .B1(new_n883_), .B2(new_n889_), .ZN(G1348gat));
  AOI21_X1  g689(.A(G176gat), .B1(new_n882_), .B2(new_n652_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n414_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n879_), .A2(new_n651_), .A3(new_n231_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(G1349gat));
  INV_X1    g693(.A(new_n882_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n895_), .A2(new_n427_), .A3(new_n621_), .ZN(new_n896_));
  INV_X1    g695(.A(G183gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n892_), .A2(new_n620_), .A3(new_n878_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n896_), .B1(new_n897_), .B2(new_n898_), .ZN(G1350gat));
  AND3_X1   g698(.A1(new_n882_), .A2(new_n426_), .A3(new_n660_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n211_), .B1(new_n882_), .B2(new_n597_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902_));
  OR3_X1    g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1351gat));
  NOR4_X1   g704(.A1(new_n272_), .A2(new_n415_), .A3(new_n348_), .A4(new_n472_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n827_), .A2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n549_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(new_n364_), .ZN(G1352gat));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n651_), .ZN(new_n910_));
  XOR2_X1   g709(.A(KEYINPUT126), .B(G204gat), .Z(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1353gat));
  INV_X1    g711(.A(new_n907_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n621_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT127), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n915_), .B(new_n917_), .ZN(G1354gat));
  OR3_X1    g717(.A1(new_n907_), .A2(G218gat), .A3(new_n661_), .ZN(new_n919_));
  OAI21_X1  g718(.A(G218gat), .B1(new_n907_), .B2(new_n684_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1355gat));
endmodule


