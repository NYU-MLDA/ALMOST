//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n945_, new_n946_, new_n948_,
    new_n949_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n959_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n982_, new_n983_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n997_, new_n998_,
    new_n1000_, new_n1001_, new_n1002_, new_n1004_, new_n1005_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  XOR2_X1   g001(.A(G190gat), .B(G218gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT36), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT71), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n208_), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT9), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G85gat), .B(G92gat), .Z(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT9), .ZN(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT10), .B(G99gat), .Z(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n216_), .B(new_n218_), .C1(G106gat), .C2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NOR3_X1   g022(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n225_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT8), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(new_n217_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT65), .B1(new_n209_), .B2(new_n211_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n233_), .A3(new_n225_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n227_), .B1(new_n234_), .B2(new_n217_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n228_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  AOI211_X1 g036(.A(KEYINPUT66), .B(new_n227_), .C1(new_n234_), .C2(new_n217_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n221_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G29gat), .B(G36gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G43gat), .B(G50gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT15), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT69), .ZN(new_n245_));
  INV_X1    g044(.A(new_n239_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT35), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G232gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT34), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n246_), .A2(new_n242_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n247_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n245_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n253_), .B1(new_n245_), .B2(new_n251_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n207_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n245_), .A2(new_n251_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n252_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT36), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n205_), .A2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n261_), .B(KEYINPUT70), .Z(new_n262_));
  NAND3_X1  g061(.A1(new_n259_), .A2(new_n254_), .A3(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n202_), .B1(new_n257_), .B2(new_n263_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n259_), .A2(new_n254_), .A3(new_n262_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n206_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n266_), .B1(new_n259_), .B2(new_n254_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n264_), .B1(new_n268_), .B2(new_n202_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G57gat), .B(G64gat), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n270_), .A2(KEYINPUT11), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(KEYINPUT11), .ZN(new_n272_));
  XOR2_X1   g071(.A(G71gat), .B(G78gat), .Z(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n272_), .A2(new_n273_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G231gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G15gat), .B(G22gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G1gat), .A2(G8gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT14), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G1gat), .B(G8gat), .Z(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n282_), .A2(KEYINPUT72), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n285_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n287_), .B1(new_n285_), .B2(new_n288_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n278_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT17), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G127gat), .B(G155gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT16), .ZN(new_n296_));
  XOR2_X1   g095(.A(G183gat), .B(G211gat), .Z(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n293_), .A2(new_n294_), .A3(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(KEYINPUT17), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n293_), .A2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n303_), .A2(KEYINPUT73), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(KEYINPUT73), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT74), .B1(new_n269_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n207_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(new_n259_), .B2(new_n254_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT37), .B1(new_n265_), .B2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n206_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(new_n263_), .A3(new_n202_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n314_));
  INV_X1    g113(.A(new_n306_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT13), .ZN(new_n317_));
  XOR2_X1   g116(.A(G120gat), .B(G148gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(G176gat), .B(G204gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n276_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n239_), .A2(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n221_), .B(new_n276_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(KEYINPUT12), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT12), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n239_), .A2(new_n327_), .A3(new_n323_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G230gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT64), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n331_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n322_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n331_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n322_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n337_), .A2(new_n333_), .A3(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n317_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n332_), .A2(new_n334_), .A3(new_n322_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n338_), .B1(new_n337_), .B2(new_n333_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(KEYINPUT13), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT68), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT68), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n307_), .A2(new_n316_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355_));
  XOR2_X1   g154(.A(G141gat), .B(G148gat), .Z(new_n356_));
  INV_X1    g155(.A(G155gat), .ZN(new_n357_));
  INV_X1    g156(.A(G162gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT82), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(G155gat), .A3(G162gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT1), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n364_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT83), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n359_), .B(new_n365_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  AOI211_X1 g167(.A(KEYINPUT83), .B(new_n364_), .C1(new_n361_), .C2(new_n363_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n356_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372_));
  NOR2_X1   g171(.A1(G141gat), .A2(G148gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n372_), .B1(new_n373_), .B2(KEYINPUT84), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT84), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n375_), .A2(G141gat), .A3(G148gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n371_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G141gat), .ZN(new_n378_));
  INV_X1    g177(.A(G148gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT2), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT2), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(G141gat), .A3(G148gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n373_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n380_), .A2(new_n382_), .B1(new_n383_), .B2(KEYINPUT3), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n373_), .A2(KEYINPUT84), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n375_), .B1(G141gat), .B2(G148gat), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n385_), .A2(KEYINPUT85), .A3(new_n386_), .A4(new_n372_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n377_), .A2(new_n384_), .A3(new_n387_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n361_), .A2(new_n363_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n355_), .B1(new_n370_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G211gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT88), .B1(new_n393_), .B2(G218gat), .ZN(new_n394_));
  INV_X1    g193(.A(G218gat), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n395_), .A2(G211gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(G197gat), .ZN(new_n398_));
  INV_X1    g197(.A(G204gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G197gat), .A2(G204gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(KEYINPUT21), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT21), .ZN(new_n403_));
  AND2_X1   g202(.A1(G197gat), .A2(G204gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(G197gat), .A2(G204gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n397_), .A2(new_n402_), .A3(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n404_), .A2(new_n405_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n408_), .B(KEYINPUT21), .C1(new_n396_), .C2(new_n394_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n412_));
  OAI21_X1  g211(.A(G228gat), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n413_), .B(KEYINPUT89), .Z(new_n414_));
  OR3_X1    g213(.A1(new_n392_), .A2(new_n410_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(KEYINPUT89), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(new_n392_), .B2(new_n410_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n354_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT83), .B1(new_n389_), .B2(new_n364_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n365_), .A2(new_n359_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n366_), .A2(new_n367_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n424_), .A2(new_n356_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n420_), .B1(new_n425_), .B2(new_n355_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n355_), .A3(new_n420_), .ZN(new_n428_));
  XOR2_X1   g227(.A(G22gat), .B(G50gat), .Z(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n429_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n370_), .A2(new_n391_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n432_), .A2(KEYINPUT29), .A3(new_n419_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n433_), .B2(new_n426_), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n418_), .A2(KEYINPUT90), .B1(new_n430_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n417_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n392_), .A2(new_n410_), .A3(new_n414_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n353_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n415_), .A2(new_n354_), .A3(new_n417_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n438_), .A2(new_n439_), .A3(new_n430_), .A4(new_n434_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT91), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n430_), .A2(new_n434_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT91), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n442_), .A2(new_n444_), .A3(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(G8gat), .B(G36gat), .Z(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT18), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G64gat), .B(G92gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n454_));
  INV_X1    g253(.A(G176gat), .ZN(new_n455_));
  INV_X1    g254(.A(G169gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT22), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT22), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(G169gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT92), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n457_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n460_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n455_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  AND3_X1   g262(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(G183gat), .ZN(new_n467_));
  INV_X1    g266(.A(G190gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n466_), .A2(new_n469_), .B1(G169gat), .B2(G176gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n463_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G183gat), .A2(G190gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT23), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT26), .B(G190gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT25), .B(G183gat), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n476_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n456_), .A2(new_n455_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G169gat), .A2(G176gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(KEYINPUT24), .A3(new_n481_), .ZN(new_n482_));
  OR3_X1    g281(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n471_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n407_), .A2(new_n409_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n454_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G226gat), .A2(G233gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT19), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n467_), .A2(KEYINPUT78), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT78), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(G183gat), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n492_), .A2(new_n494_), .A3(new_n468_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT79), .B1(new_n495_), .B2(new_n476_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n492_), .A2(new_n494_), .A3(new_n468_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT79), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n466_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(new_n456_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n496_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT25), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n504_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n477_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(new_n484_), .A3(new_n466_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n410_), .A3(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n488_), .A2(new_n491_), .A3(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT97), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n410_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n463_), .A2(new_n470_), .B1(new_n479_), .B2(new_n484_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n454_), .B1(new_n513_), .B2(new_n410_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n512_), .B1(new_n515_), .B2(KEYINPUT96), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n491_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n453_), .B1(new_n511_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT20), .B1(new_n513_), .B2(new_n410_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n503_), .A2(new_n410_), .A3(new_n508_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n490_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n466_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n498_), .B1(new_n466_), .B2(new_n497_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n524_), .A2(new_n525_), .A3(new_n501_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n466_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n506_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n492_), .A2(new_n494_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n528_), .B1(new_n529_), .B2(new_n504_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n527_), .B1(new_n530_), .B2(new_n477_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n487_), .B1(new_n526_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n514_), .A2(new_n532_), .A3(new_n491_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n523_), .A2(new_n452_), .A3(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n534_), .A2(KEYINPUT27), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT93), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n523_), .A2(new_n533_), .A3(KEYINPUT93), .A4(new_n452_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n533_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n491_), .B1(new_n488_), .B2(new_n509_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n453_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n538_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT27), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n520_), .A2(new_n535_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n448_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G71gat), .B(G99gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(G43gat), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n503_), .A2(new_n508_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n547_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G227gat), .A2(G233gat), .ZN(new_n551_));
  INV_X1    g350(.A(G15gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT30), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT81), .ZN(new_n556_));
  INV_X1    g355(.A(new_n554_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n548_), .A2(new_n549_), .A3(new_n557_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n555_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n556_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G127gat), .B(G134gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G113gat), .B(G120gat), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(KEYINPUT80), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT80), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n562_), .A2(new_n563_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT31), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n560_), .A2(new_n561_), .A3(new_n570_), .ZN(new_n571_));
  OR4_X1    g370(.A1(new_n556_), .A2(new_n555_), .A3(new_n558_), .A4(new_n570_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n370_), .A2(new_n391_), .B1(new_n568_), .B2(new_n566_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n564_), .A2(new_n565_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n575_), .B1(new_n425_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G225gat), .A2(G233gat), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT4), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n578_), .B1(new_n575_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT94), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n370_), .A2(new_n391_), .A3(new_n576_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n569_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n583_), .B(KEYINPUT4), .C1(new_n425_), .C2(new_n584_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n581_), .A2(new_n582_), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n582_), .B1(new_n581_), .B2(new_n585_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n579_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G1gat), .B(G29gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G57gat), .B(G85gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n588_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n593_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT98), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT98), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n598_), .B(new_n595_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n574_), .A2(new_n594_), .A3(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n545_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n442_), .A2(new_n444_), .A3(new_n447_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n603_), .A2(new_n544_), .A3(new_n594_), .A4(new_n600_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n581_), .A2(new_n585_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT94), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n581_), .A2(new_n585_), .A3(new_n582_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n598_), .B1(new_n608_), .B2(new_n595_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n599_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n594_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(KEYINPUT32), .B(new_n452_), .C1(new_n511_), .C2(new_n519_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n452_), .A2(KEYINPUT32), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n523_), .A2(new_n533_), .A3(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n578_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n575_), .B2(new_n580_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n585_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n583_), .B(new_n616_), .C1(new_n425_), .C2(new_n584_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n593_), .A3(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n620_), .A2(new_n537_), .A3(new_n538_), .A4(new_n541_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n622_), .B2(new_n596_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n608_), .A2(KEYINPUT33), .A3(new_n595_), .ZN(new_n624_));
  AOI22_X1  g423(.A1(new_n611_), .A2(new_n615_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n604_), .B1(new_n625_), .B2(new_n603_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n602_), .B1(new_n626_), .B2(new_n573_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n242_), .B(KEYINPUT76), .Z(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n242_), .B(KEYINPUT76), .ZN(new_n630_));
  INV_X1    g429(.A(new_n291_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n630_), .B1(new_n631_), .B2(new_n289_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(G229gat), .A3(G233gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n243_), .B1(new_n631_), .B2(new_n289_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT77), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n629_), .A2(new_n635_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n634_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G113gat), .B(G141gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G169gat), .B(G197gat), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n640_), .B(new_n641_), .Z(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n634_), .A2(new_n638_), .A3(new_n642_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n627_), .A2(new_n647_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n307_), .A2(new_n349_), .A3(KEYINPUT75), .A4(new_n316_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n611_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(G1gat), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n352_), .A2(new_n648_), .A3(new_n649_), .A4(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT99), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n649_), .A2(new_n648_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n352_), .A4(new_n651_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n653_), .A2(new_n656_), .A3(KEYINPUT38), .ZN(new_n657_));
  INV_X1    g456(.A(new_n268_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n612_), .A2(new_n614_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n600_), .B2(new_n594_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n624_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT33), .B1(new_n608_), .B2(new_n595_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n661_), .A2(new_n662_), .A3(new_n621_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n448_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n574_), .B1(new_n664_), .B2(new_n604_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n658_), .B1(new_n665_), .B2(new_n602_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n340_), .A2(new_n343_), .A3(new_n646_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT100), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n340_), .A2(new_n343_), .A3(new_n669_), .A4(new_n646_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n302_), .A3(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n666_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n611_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G1gat), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n657_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT38), .B1(new_n653_), .B2(new_n656_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT102), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n678_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n680_), .A2(new_n681_), .A3(new_n676_), .A4(new_n657_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(G1324gat));
  NOR2_X1   g482(.A1(new_n544_), .A2(G8gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n654_), .A2(new_n352_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT103), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n654_), .A2(new_n687_), .A3(new_n352_), .A4(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(G8gat), .ZN(new_n690_));
  INV_X1    g489(.A(new_n544_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n672_), .B2(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT39), .Z(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n689_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n689_), .B2(new_n693_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1325gat));
  NAND2_X1  g496(.A1(new_n654_), .A2(new_n352_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(new_n552_), .A3(new_n574_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n701_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n552_), .B1(new_n672_), .B2(new_n574_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n705_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n702_), .A2(new_n703_), .A3(new_n706_), .A4(new_n707_), .ZN(G1326gat));
  INV_X1    g507(.A(G22gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n672_), .B2(new_n603_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT42), .Z(new_n711_));
  NAND2_X1  g510(.A1(new_n603_), .A2(new_n709_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n698_), .B2(new_n712_), .ZN(G1327gat));
  NAND2_X1  g512(.A1(new_n306_), .A2(new_n268_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n714_), .A2(new_n344_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n648_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G29gat), .B1(new_n717_), .B2(new_n611_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n269_), .B(new_n719_), .C1(new_n665_), .C2(new_n602_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n611_), .A2(new_n615_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n623_), .A2(new_n624_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n603_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n604_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n573_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n602_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n313_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n719_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n720_), .B1(new_n727_), .B2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n668_), .A2(new_n306_), .A3(new_n670_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n668_), .A2(KEYINPUT106), .A3(new_n306_), .A4(new_n670_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n731_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT44), .B1(new_n737_), .B2(KEYINPUT108), .ZN(new_n740_));
  INV_X1    g539(.A(new_n730_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n741_), .B1(new_n627_), .B2(new_n313_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n742_), .A2(new_n720_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n739_), .B1(new_n740_), .B2(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n611_), .A2(G29gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n718_), .B1(new_n746_), .B2(new_n747_), .ZN(G1328gat));
  NAND2_X1  g547(.A1(new_n737_), .A2(KEYINPUT108), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(new_n738_), .A3(new_n745_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n743_), .A2(KEYINPUT44), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n691_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G36gat), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n691_), .A2(KEYINPUT109), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n691_), .A2(KEYINPUT109), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(G36gat), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OR3_X1    g557(.A1(new_n716_), .A2(KEYINPUT110), .A3(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT110), .B1(new_n716_), .B2(new_n758_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(KEYINPUT45), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n760_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n753_), .A2(KEYINPUT46), .A3(new_n761_), .A4(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n757_), .B1(new_n746_), .B2(new_n691_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n761_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n765_), .A2(new_n769_), .ZN(G1329gat));
  AND2_X1   g569(.A1(new_n574_), .A2(G43gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n738_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n731_), .A2(new_n744_), .A3(new_n736_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n751_), .B(new_n771_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT111), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n750_), .A2(new_n776_), .A3(new_n751_), .A4(new_n771_), .ZN(new_n777_));
  XOR2_X1   g576(.A(KEYINPUT112), .B(G43gat), .Z(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(new_n716_), .B2(new_n573_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT47), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n775_), .A2(new_n777_), .A3(new_n782_), .A4(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1330gat));
  AOI21_X1  g583(.A(G50gat), .B1(new_n717_), .B2(new_n603_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n603_), .A2(G50gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n746_), .B2(new_n786_), .ZN(G1331gat));
  NOR2_X1   g586(.A1(new_n627_), .A2(new_n646_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n788_), .A2(new_n307_), .A3(new_n316_), .A4(new_n344_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(new_n650_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n304_), .A2(new_n305_), .A3(new_n647_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n666_), .A2(new_n349_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(G57gat), .B1(new_n650_), .B2(KEYINPUT113), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(KEYINPUT113), .B2(G57gat), .ZN(new_n795_));
  OAI22_X1  g594(.A1(new_n790_), .A2(G57gat), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT114), .ZN(G1332gat));
  INV_X1    g596(.A(new_n756_), .ZN(new_n798_));
  OAI21_X1  g597(.A(G64gat), .B1(new_n793_), .B2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT48), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(G64gat), .ZN(new_n801_));
  XOR2_X1   g600(.A(new_n801_), .B(KEYINPUT115), .Z(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n789_), .B2(new_n802_), .ZN(G1333gat));
  OR3_X1    g602(.A1(new_n789_), .A2(G71gat), .A3(new_n573_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n792_), .A2(new_n574_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT116), .B(KEYINPUT49), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n805_), .A2(G71gat), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n805_), .B2(G71gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(G1334gat));
  OAI21_X1  g608(.A(G78gat), .B1(new_n793_), .B2(new_n448_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT50), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n448_), .A2(G78gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n789_), .B2(new_n812_), .ZN(G1335gat));
  NOR3_X1   g612(.A1(new_n315_), .A2(new_n345_), .A3(new_n646_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n731_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(G85gat), .B1(new_n816_), .B2(new_n650_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n349_), .A2(new_n714_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n788_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(new_n213_), .A3(new_n611_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n821_), .ZN(G1336gat));
  OAI21_X1  g621(.A(G92gat), .B1(new_n816_), .B2(new_n798_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n214_), .A3(new_n691_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(G1337gat));
  NOR3_X1   g624(.A1(new_n819_), .A2(new_n220_), .A3(new_n573_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n815_), .A2(new_n574_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(G99gat), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT51), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n828_), .B(new_n830_), .ZN(G1338gat));
  INV_X1    g630(.A(G106gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n820_), .A2(new_n832_), .A3(new_n603_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n815_), .A2(new_n603_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(G106gat), .ZN(new_n836_));
  AOI211_X1 g635(.A(KEYINPUT52), .B(new_n832_), .C1(new_n815_), .C2(new_n603_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n833_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT53), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n840_), .B(new_n833_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(G1339gat));
  NOR2_X1   g641(.A1(new_n791_), .A2(new_n344_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n313_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n844_), .A2(KEYINPUT54), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(KEYINPUT54), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n326_), .A2(new_n336_), .A3(new_n328_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n337_), .B1(KEYINPUT55), .B2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n329_), .A2(KEYINPUT55), .A3(new_n331_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT56), .B(new_n338_), .C1(new_n849_), .C2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n338_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n855_), .A2(new_n853_), .A3(new_n856_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n861_));
  INV_X1    g660(.A(new_n637_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n629_), .A2(new_n635_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n643_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n629_), .B2(new_n632_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT118), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n865_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n643_), .A4(new_n863_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(new_n869_), .A3(new_n645_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n861_), .B1(new_n871_), .B2(new_n341_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n339_), .A2(new_n870_), .A3(KEYINPUT119), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n860_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n874_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT58), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n878_), .A2(new_n269_), .A3(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n341_), .A2(new_n646_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n848_), .A2(KEYINPUT55), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n332_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n850_), .ZN(new_n886_));
  AOI21_X1  g685(.A(KEYINPUT56), .B1(new_n886_), .B2(new_n338_), .ZN(new_n887_));
  AOI211_X1 g686(.A(new_n856_), .B(new_n322_), .C1(new_n885_), .C2(new_n850_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n883_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n870_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT57), .B1(new_n892_), .B2(new_n658_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894_));
  AOI211_X1 g693(.A(new_n894_), .B(new_n268_), .C1(new_n889_), .C2(new_n891_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n881_), .A2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n847_), .B1(new_n897_), .B2(new_n303_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n545_), .A2(new_n650_), .A3(new_n573_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT59), .B1(new_n898_), .B2(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n900_), .A2(KEYINPUT59), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n315_), .B1(new_n881_), .B2(new_n896_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n847_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G113gat), .B1(new_n905_), .B2(new_n647_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n269_), .B1(new_n879_), .B2(KEYINPUT58), .ZN(new_n907_));
  AOI211_X1 g706(.A(new_n877_), .B(new_n874_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n882_), .B1(new_n857_), .B2(new_n852_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n658_), .B1(new_n910_), .B2(new_n890_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n894_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n892_), .A2(KEYINPUT57), .A3(new_n658_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n303_), .B1(new_n909_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n847_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n900_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n647_), .A2(G113gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n906_), .B1(new_n918_), .B2(new_n919_), .ZN(G1340gat));
  INV_X1    g719(.A(new_n349_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n904_), .B(new_n921_), .C1(new_n917_), .C2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(KEYINPUT121), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n901_), .A2(new_n925_), .A3(new_n921_), .A4(new_n904_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n924_), .A2(G120gat), .A3(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(G120gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n928_), .B1(new_n345_), .B2(KEYINPUT60), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n917_), .B(new_n929_), .C1(KEYINPUT60), .C2(new_n928_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n927_), .A2(new_n930_), .ZN(G1341gat));
  INV_X1    g730(.A(G127gat), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n932_), .B1(new_n918_), .B2(new_n306_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(KEYINPUT122), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n935_), .B(new_n932_), .C1(new_n918_), .C2(new_n306_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n905_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n303_), .A2(new_n932_), .ZN(new_n938_));
  AOI22_X1  g737(.A1(new_n934_), .A2(new_n936_), .B1(new_n937_), .B2(new_n938_), .ZN(G1342gat));
  OAI21_X1  g738(.A(G134gat), .B1(new_n905_), .B2(new_n313_), .ZN(new_n940_));
  OR2_X1    g739(.A1(new_n658_), .A2(G134gat), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n918_), .B2(new_n941_), .ZN(G1343gat));
  NOR3_X1   g741(.A1(new_n756_), .A2(new_n448_), .A3(new_n650_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n302_), .B1(new_n881_), .B2(new_n896_), .ZN(new_n944_));
  OAI211_X1 g743(.A(new_n573_), .B(new_n943_), .C1(new_n944_), .C2(new_n847_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n647_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(new_n378_), .ZN(G1344gat));
  NOR2_X1   g746(.A1(new_n945_), .A2(new_n349_), .ZN(new_n948_));
  XOR2_X1   g747(.A(KEYINPUT123), .B(G148gat), .Z(new_n949_));
  XNOR2_X1  g748(.A(new_n948_), .B(new_n949_), .ZN(G1345gat));
  OAI21_X1  g749(.A(KEYINPUT124), .B1(new_n945_), .B2(new_n306_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n574_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n953_));
  NAND4_X1  g752(.A1(new_n952_), .A2(new_n953_), .A3(new_n315_), .A4(new_n943_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(KEYINPUT61), .B(G155gat), .ZN(new_n955_));
  AND3_X1   g754(.A1(new_n951_), .A2(new_n954_), .A3(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n955_), .B1(new_n951_), .B2(new_n954_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1346gat));
  OAI21_X1  g757(.A(G162gat), .B1(new_n945_), .B2(new_n313_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n268_), .A2(new_n358_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n945_), .B2(new_n960_), .ZN(G1347gat));
  NAND2_X1  g760(.A1(new_n897_), .A2(new_n306_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(new_n916_), .ZN(new_n963_));
  NOR3_X1   g762(.A1(new_n798_), .A2(new_n603_), .A3(new_n601_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n963_), .A2(new_n646_), .A3(new_n964_), .ZN(new_n965_));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n966_));
  AND3_X1   g765(.A1(new_n965_), .A2(new_n966_), .A3(G169gat), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n963_), .A2(new_n964_), .ZN(new_n968_));
  INV_X1    g767(.A(new_n968_), .ZN(new_n969_));
  OAI211_X1 g768(.A(new_n969_), .B(new_n646_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n966_), .B1(new_n965_), .B2(G169gat), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n967_), .B1(new_n970_), .B2(new_n971_), .ZN(G1348gat));
  NAND2_X1  g771(.A1(new_n915_), .A2(new_n916_), .ZN(new_n973_));
  AND2_X1   g772(.A1(new_n973_), .A2(new_n964_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n349_), .A2(new_n455_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n974_), .A2(new_n975_), .ZN(new_n976_));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n976_), .A2(new_n977_), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n974_), .A2(KEYINPUT125), .A3(new_n975_), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n455_), .B1(new_n968_), .B2(new_n345_), .ZN(new_n980_));
  AND3_X1   g779(.A1(new_n978_), .A2(new_n979_), .A3(new_n980_), .ZN(G1349gat));
  NOR3_X1   g780(.A1(new_n968_), .A2(new_n303_), .A3(new_n478_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n974_), .A2(new_n315_), .ZN(new_n983_));
  AOI21_X1  g782(.A(new_n982_), .B1(new_n529_), .B2(new_n983_), .ZN(G1350gat));
  NAND3_X1  g783(.A1(new_n969_), .A2(new_n268_), .A3(new_n477_), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n963_), .A2(new_n269_), .A3(new_n964_), .ZN(new_n986_));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n987_));
  AND3_X1   g786(.A1(new_n986_), .A2(new_n987_), .A3(G190gat), .ZN(new_n988_));
  AOI21_X1  g787(.A(new_n987_), .B1(new_n986_), .B2(G190gat), .ZN(new_n989_));
  OAI21_X1  g788(.A(new_n985_), .B1(new_n988_), .B2(new_n989_), .ZN(G1351gat));
  NOR3_X1   g789(.A1(new_n798_), .A2(new_n448_), .A3(new_n611_), .ZN(new_n991_));
  NAND3_X1  g790(.A1(new_n952_), .A2(new_n646_), .A3(new_n991_), .ZN(new_n992_));
  AND2_X1   g791(.A1(new_n398_), .A2(KEYINPUT127), .ZN(new_n993_));
  NOR2_X1   g792(.A1(new_n992_), .A2(new_n993_), .ZN(new_n994_));
  XOR2_X1   g793(.A(KEYINPUT127), .B(G197gat), .Z(new_n995_));
  AOI21_X1  g794(.A(new_n994_), .B1(new_n992_), .B2(new_n995_), .ZN(G1352gat));
  NAND2_X1  g795(.A1(new_n952_), .A2(new_n991_), .ZN(new_n997_));
  NOR2_X1   g796(.A1(new_n997_), .A2(new_n349_), .ZN(new_n998_));
  XNOR2_X1  g797(.A(new_n998_), .B(new_n399_), .ZN(G1353gat));
  NAND3_X1  g798(.A1(new_n952_), .A2(new_n302_), .A3(new_n991_), .ZN(new_n1000_));
  OAI21_X1  g799(.A(new_n1000_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1001_));
  XOR2_X1   g800(.A(KEYINPUT63), .B(G211gat), .Z(new_n1002_));
  OAI21_X1  g801(.A(new_n1001_), .B1(new_n1000_), .B2(new_n1002_), .ZN(G1354gat));
  OAI21_X1  g802(.A(G218gat), .B1(new_n997_), .B2(new_n313_), .ZN(new_n1004_));
  NAND2_X1  g803(.A1(new_n268_), .A2(new_n395_), .ZN(new_n1005_));
  OAI21_X1  g804(.A(new_n1004_), .B1(new_n997_), .B2(new_n1005_), .ZN(G1355gat));
endmodule


