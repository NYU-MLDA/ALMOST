//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n961_, new_n962_, new_n964_, new_n965_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n979_, new_n980_, new_n981_;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n202_));
  INV_X1    g001(.A(G183gat), .ZN(new_n203_));
  INV_X1    g002(.A(G190gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n204_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209_));
  INV_X1    g008(.A(G176gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT26), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT75), .B1(new_n217_), .B2(G190gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT26), .B(G190gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n216_), .B(new_n218_), .C1(new_n219_), .C2(KEYINPUT75), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(new_n212_), .A3(new_n210_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n205_), .A2(new_n207_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n212_), .A2(new_n210_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(KEYINPUT24), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT76), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n221_), .B1(G169gat), .B2(G176gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(KEYINPUT76), .A3(new_n226_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n215_), .B1(new_n225_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G71gat), .B(G99gat), .ZN(new_n235_));
  INV_X1    g034(.A(G43gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n234_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT77), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n239_), .A2(new_n240_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n239_), .A2(new_n240_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n242_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n238_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250_));
  INV_X1    g049(.A(G15gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT30), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT31), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n249_), .B(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT86), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT85), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n215_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n208_), .A2(KEYINPUT85), .A3(new_n214_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n219_), .A2(new_n216_), .B1(new_n231_), .B2(new_n226_), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n259_), .A2(new_n260_), .B1(new_n224_), .B2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G211gat), .B(G218gat), .Z(new_n263_));
  INV_X1    g062(.A(G197gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(G204gat), .ZN(new_n265_));
  INV_X1    g064(.A(G204gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(G197gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n263_), .A2(KEYINPUT21), .A3(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n264_), .A2(KEYINPUT82), .A3(G204gat), .ZN(new_n270_));
  OAI211_X1 g069(.A(KEYINPUT21), .B(new_n270_), .C1(new_n268_), .C2(KEYINPUT82), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G211gat), .B(G218gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(new_n268_), .B2(KEYINPUT21), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n269_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n257_), .B1(new_n262_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT20), .ZN(new_n277_));
  INV_X1    g076(.A(new_n215_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n216_), .A2(new_n218_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT75), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n217_), .A2(G190gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n204_), .A2(KEYINPUT26), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n280_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n223_), .B1(new_n279_), .B2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n230_), .A2(new_n232_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n278_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n277_), .B1(new_n286_), .B2(new_n275_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n261_), .A2(new_n224_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n260_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT85), .B1(new_n208_), .B2(new_n214_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n263_), .A2(KEYINPUT21), .A3(new_n268_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n271_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n292_), .B1(new_n293_), .B2(new_n273_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n291_), .A2(KEYINPUT86), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G226gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT19), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT84), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n276_), .A2(new_n287_), .A3(new_n295_), .A4(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n288_), .A2(new_n215_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n294_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(new_n286_), .B2(new_n275_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n234_), .A2(KEYINPUT88), .A3(new_n294_), .ZN(new_n304_));
  AOI211_X1 g103(.A(new_n277_), .B(new_n301_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n297_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n299_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G8gat), .B(G36gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT18), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G64gat), .B(G92gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT27), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n277_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT89), .B1(new_n291_), .B2(new_n294_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT89), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n262_), .A2(new_n316_), .A3(new_n275_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n314_), .A2(new_n306_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n311_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n276_), .A2(new_n287_), .A3(new_n295_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT87), .ZN(new_n322_));
  INV_X1    g121(.A(new_n298_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n322_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n319_), .B(new_n320_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT94), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n321_), .A2(new_n323_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT87), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT94), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(new_n319_), .A4(new_n320_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n313_), .B1(new_n327_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT93), .ZN(new_n335_));
  INV_X1    g134(.A(G141gat), .ZN(new_n336_));
  INV_X1    g135(.A(G148gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT80), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n336_), .B(new_n337_), .C1(new_n338_), .C2(KEYINPUT3), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n340_), .B(KEYINPUT80), .C1(G141gat), .C2(G148gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346_));
  NAND3_X1  g145(.A1(KEYINPUT78), .A2(G141gat), .A3(G148gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n343_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT2), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n342_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT81), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n354_), .A2(new_n359_), .A3(new_n355_), .A4(new_n356_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n351_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n345_), .A2(new_n347_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n356_), .B(KEYINPUT1), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n354_), .A2(new_n355_), .ZN(new_n365_));
  OAI221_X1 g164(.A(new_n363_), .B1(G141gat), .B2(G148gat), .C1(new_n364_), .C2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n248_), .A2(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n244_), .A2(new_n361_), .A3(new_n366_), .A4(new_n247_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(KEYINPUT4), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n248_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT90), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n370_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n368_), .A2(new_n369_), .A3(new_n373_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT91), .B(G85gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT0), .B(G57gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n375_), .A2(new_n376_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n335_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n375_), .A2(new_n376_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n381_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n388_), .A2(new_n382_), .A3(KEYINPUT93), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT83), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n294_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT29), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n393_), .B1(new_n361_), .B2(new_n366_), .ZN(new_n394_));
  OAI21_X1  g193(.A(G78gat), .B1(new_n394_), .B2(new_n275_), .ZN(new_n395_));
  INV_X1    g194(.A(G78gat), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n339_), .A2(new_n341_), .B1(new_n349_), .B2(KEYINPUT2), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n397_), .A2(new_n348_), .B1(new_n357_), .B2(KEYINPUT81), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n364_), .A2(new_n365_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n362_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n398_), .A2(new_n360_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n396_), .B(new_n294_), .C1(new_n401_), .C2(new_n393_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n395_), .A2(new_n402_), .A3(G106gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(G106gat), .B1(new_n395_), .B2(new_n402_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n392_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n395_), .A2(new_n402_), .ZN(new_n406_));
  INV_X1    g205(.A(G106gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n395_), .A2(new_n402_), .A3(G106gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n392_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  OR3_X1    g210(.A1(new_n367_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT28), .B1(new_n367_), .B2(KEYINPUT29), .ZN(new_n413_));
  XOR2_X1   g212(.A(G22gat), .B(G50gat), .Z(new_n414_));
  AND3_X1   g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n405_), .A2(new_n411_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(new_n405_), .B2(new_n411_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n385_), .B(new_n389_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n319_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n311_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT27), .B1(new_n422_), .B2(new_n326_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n334_), .A2(new_n420_), .A3(new_n423_), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n418_), .A2(new_n419_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n383_), .A2(KEYINPUT33), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n370_), .A2(new_n373_), .A3(new_n372_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n368_), .A2(new_n369_), .A3(new_n374_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n387_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT33), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n382_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n422_), .A2(new_n326_), .A3(new_n426_), .A4(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT92), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n324_), .A2(new_n325_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT32), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n319_), .B1(new_n435_), .B2(new_n311_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n433_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n311_), .A2(new_n435_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n382_), .A2(new_n388_), .B1(new_n307_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n303_), .A2(new_n304_), .ZN(new_n440_));
  AND4_X1   g239(.A1(KEYINPUT20), .A2(new_n440_), .A3(new_n318_), .A4(new_n306_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n441_), .A2(new_n438_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(new_n331_), .A3(KEYINPUT92), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n437_), .A2(new_n439_), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n425_), .B1(new_n432_), .B2(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(KEYINPUT95), .B(new_n256_), .C1(new_n424_), .C2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n385_), .A2(new_n389_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n448_), .A2(new_n256_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n334_), .A2(new_n423_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n425_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n446_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n420_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n327_), .A2(new_n333_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n313_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n423_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n444_), .A2(new_n432_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n451_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT95), .B1(new_n462_), .B2(new_n256_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n453_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G113gat), .B(G141gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G169gat), .B(G197gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  NAND2_X1  g266(.A1(G229gat), .A2(G233gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G29gat), .B(G36gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G43gat), .B(G50gat), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n471_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G1gat), .B(G8gat), .Z(new_n475_));
  OR2_X1    g274(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G22gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n476_), .A2(G22gat), .A3(new_n477_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G1gat), .ZN(new_n483_));
  INV_X1    g282(.A(G8gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n475_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n482_), .A2(new_n475_), .A3(new_n485_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n474_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n488_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n472_), .A2(new_n473_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n490_), .A2(new_n486_), .A3(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n469_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(KEYINPUT15), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT15), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n474_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n494_), .B(new_n496_), .C1(new_n490_), .C2(new_n486_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n487_), .A2(new_n474_), .A3(new_n488_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n468_), .A3(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n493_), .A2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n467_), .B1(new_n500_), .B2(KEYINPUT74), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT74), .ZN(new_n502_));
  INV_X1    g301(.A(new_n467_), .ZN(new_n503_));
  AOI211_X1 g302(.A(new_n502_), .B(new_n503_), .C1(new_n493_), .C2(new_n499_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n464_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT67), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT8), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT66), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n510_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT6), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT7), .ZN(new_n520_));
  INV_X1    g319(.A(G99gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n407_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(KEYINPUT66), .A3(new_n511_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n514_), .A2(new_n519_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(G85gat), .ZN(new_n525_));
  INV_X1    g324(.A(G92gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n509_), .B1(new_n524_), .B2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n529_), .A2(KEYINPUT8), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n516_), .A2(new_n518_), .A3(KEYINPUT64), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT64), .B1(new_n516_), .B2(new_n518_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n522_), .A2(new_n511_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n533_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n508_), .B1(new_n531_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT64), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n519_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n516_), .A2(new_n518_), .A3(KEYINPUT64), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n538_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n532_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n537_), .A2(new_n510_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n529_), .B1(new_n546_), .B2(new_n523_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n545_), .B(KEYINPUT67), .C1(new_n547_), .C2(new_n509_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n540_), .A2(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n407_), .A3(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n527_), .A2(KEYINPUT9), .A3(new_n528_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n528_), .A2(KEYINPUT9), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT65), .B1(new_n536_), .B2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT65), .ZN(new_n558_));
  NOR4_X1   g357(.A1(new_n557_), .A2(new_n534_), .A3(new_n535_), .A4(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n549_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G57gat), .B(G64gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT11), .ZN(new_n563_));
  XOR2_X1   g362(.A(G71gat), .B(G78gat), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n562_), .A2(KEYINPUT11), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n563_), .A2(new_n564_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT12), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n561_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n524_), .A2(new_n530_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n574_), .A2(KEYINPUT8), .B1(new_n544_), .B2(new_n532_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n542_), .A2(new_n543_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n558_), .B1(new_n576_), .B2(new_n557_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n536_), .A2(new_n555_), .A3(KEYINPUT65), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n569_), .B1(new_n575_), .B2(new_n579_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n575_), .A2(new_n579_), .A3(new_n569_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT12), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n580_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n572_), .A2(new_n573_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n573_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n567_), .A2(new_n568_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n545_), .B1(new_n547_), .B2(new_n509_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n586_), .B1(new_n560_), .B2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n585_), .B1(new_n581_), .B2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G120gat), .B(G148gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G176gat), .B(G204gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n590_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n590_), .A2(new_n596_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n584_), .A2(new_n589_), .A3(new_n596_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(KEYINPUT13), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT69), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G134gat), .B(G162gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT36), .Z(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT34), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT35), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT70), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n612_), .A2(KEYINPUT35), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n612_), .A2(KEYINPUT70), .A3(KEYINPUT35), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n575_), .A2(new_n579_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n620_), .B2(new_n474_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n579_), .B1(new_n540_), .B2(new_n548_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n494_), .A2(new_n496_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n616_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n621_), .B(new_n615_), .C1(new_n624_), .C2(new_n623_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT72), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n610_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(new_n627_), .A3(KEYINPUT72), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n608_), .A2(KEYINPUT36), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n628_), .A2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT37), .B1(new_n632_), .B2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n609_), .B(KEYINPUT71), .Z(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n634_), .B(KEYINPUT37), .C1(new_n628_), .C2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n487_), .A2(new_n488_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(new_n586_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(G231gat), .A2(G233gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT17), .ZN(new_n645_));
  XOR2_X1   g444(.A(G127gat), .B(G155gat), .Z(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT16), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G183gat), .B(G211gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  OR3_X1    g448(.A1(new_n644_), .A2(new_n645_), .A3(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(KEYINPUT17), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n644_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n640_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n605_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n507_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n483_), .A3(new_n448_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n634_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n631_), .B2(new_n630_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT96), .Z(new_n662_));
  NOR2_X1   g461(.A1(new_n464_), .A2(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n603_), .A2(new_n653_), .A3(new_n506_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G1gat), .B1(new_n665_), .B2(new_n447_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n659_), .A2(new_n666_), .ZN(new_n667_));
  MUX2_X1   g466(.A(new_n659_), .B(new_n667_), .S(KEYINPUT38), .Z(G1324gat));
  OAI21_X1  g467(.A(G8gat), .B1(new_n665_), .B2(new_n450_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT39), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n450_), .A2(G8gat), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  OR3_X1    g472(.A1(new_n657_), .A2(KEYINPUT97), .A3(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT97), .B1(new_n657_), .B2(new_n673_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n669_), .A2(new_n670_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n671_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n671_), .A2(new_n676_), .A3(KEYINPUT40), .A4(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1325gat));
  NAND3_X1  g481(.A1(new_n658_), .A2(new_n251_), .A3(new_n255_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT98), .ZN(new_n684_));
  OAI21_X1  g483(.A(G15gat), .B1(new_n665_), .B2(new_n256_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT41), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n685_), .A2(KEYINPUT41), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n686_), .A3(new_n687_), .ZN(G1326gat));
  INV_X1    g487(.A(new_n665_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n425_), .B(KEYINPUT99), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n479_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT42), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n658_), .A2(new_n479_), .A3(new_n690_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n661_), .A2(new_n653_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n603_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n507_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n448_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT101), .B1(new_n635_), .B2(new_n639_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n702_), .B(new_n638_), .C1(new_n661_), .C2(KEYINPUT37), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n704_), .B1(new_n453_), .B2(new_n463_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT95), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n420_), .A2(new_n423_), .ZN(new_n707_));
  AOI22_X1  g506(.A1(new_n707_), .A2(new_n457_), .B1(new_n460_), .B2(new_n451_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n706_), .B1(new_n708_), .B2(new_n255_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(new_n452_), .A3(new_n446_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n640_), .A2(KEYINPUT43), .ZN(new_n711_));
  AOI22_X1  g510(.A1(new_n705_), .A2(KEYINPUT43), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n599_), .A2(new_n602_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n653_), .A3(new_n505_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT100), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n700_), .B1(new_n712_), .B2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n714_), .B(KEYINPUT100), .Z(new_n717_));
  AND2_X1   g516(.A1(new_n710_), .A2(new_n711_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n710_), .B2(new_n704_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n717_), .B(KEYINPUT44), .C1(new_n718_), .C2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n716_), .A2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n448_), .A2(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n699_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  INV_X1    g523(.A(new_n450_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n716_), .A2(new_n721_), .A3(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G36gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n728_));
  NOR2_X1   g527(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n450_), .A2(G36gat), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n697_), .B2(new_n733_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n507_), .A2(new_n696_), .A3(new_n730_), .A4(new_n732_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n729_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n727_), .A2(new_n728_), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n728_), .B1(new_n727_), .B2(new_n736_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1329gat));
  NOR2_X1   g538(.A1(new_n256_), .A2(new_n236_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n716_), .A2(new_n721_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT104), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n716_), .A2(new_n721_), .A3(new_n743_), .A4(new_n740_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n236_), .B1(new_n697_), .B2(new_n256_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n742_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT47), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n742_), .A2(new_n748_), .A3(new_n744_), .A4(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1330gat));
  AOI21_X1  g549(.A(G50gat), .B1(new_n698_), .B2(new_n690_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n425_), .A2(G50gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n722_), .B2(new_n752_), .ZN(G1331gat));
  NOR2_X1   g552(.A1(new_n655_), .A2(new_n713_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT105), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n464_), .A2(new_n505_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(G57gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(new_n758_), .A3(new_n448_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n604_), .A2(new_n653_), .A3(new_n505_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n663_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G57gat), .B1(new_n761_), .B2(new_n447_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n762_), .ZN(G1332gat));
  INV_X1    g562(.A(G64gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n757_), .A2(new_n764_), .A3(new_n725_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G64gat), .B1(new_n761_), .B2(new_n450_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(KEYINPUT48), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(KEYINPUT48), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n765_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT106), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n765_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1333gat));
  OAI21_X1  g572(.A(G71gat), .B1(new_n761_), .B2(new_n256_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT49), .ZN(new_n775_));
  INV_X1    g574(.A(G71gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n757_), .A2(new_n776_), .A3(new_n255_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1334gat));
  NAND3_X1  g577(.A1(new_n663_), .A2(new_n690_), .A3(new_n760_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(G78gat), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT50), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n757_), .A2(new_n396_), .A3(new_n690_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1335gat));
  NOR3_X1   g582(.A1(new_n713_), .A2(new_n654_), .A3(new_n505_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n718_), .B2(new_n720_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n785_), .A2(new_n525_), .A3(new_n447_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n604_), .A2(new_n695_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n756_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n756_), .A2(KEYINPUT107), .A3(new_n787_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT108), .B(new_n525_), .C1(new_n792_), .C2(new_n447_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n447_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(G85gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n786_), .B1(new_n793_), .B2(new_n796_), .ZN(G1336gat));
  NOR2_X1   g596(.A1(new_n450_), .A2(new_n526_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT110), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n785_), .A2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(KEYINPUT109), .B(new_n526_), .C1(new_n792_), .C2(new_n450_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT109), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n450_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(G92gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n800_), .B1(new_n801_), .B2(new_n804_), .ZN(G1337gat));
  OAI211_X1 g604(.A(new_n255_), .B(new_n784_), .C1(new_n718_), .C2(new_n720_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n806_), .A2(new_n807_), .A3(G99gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n806_), .B2(G99gat), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n255_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n810_));
  OAI22_X1  g609(.A1(new_n808_), .A2(new_n809_), .B1(new_n792_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT51), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n813_));
  OAI221_X1 g612(.A(new_n813_), .B1(new_n792_), .B2(new_n810_), .C1(new_n809_), .C2(new_n808_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1338gat));
  OAI211_X1 g614(.A(new_n425_), .B(new_n784_), .C1(new_n718_), .C2(new_n720_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n816_), .A2(new_n817_), .A3(G106gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n816_), .B2(G106gat), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n425_), .A2(new_n407_), .ZN(new_n820_));
  OAI22_X1  g619(.A1(new_n818_), .A2(new_n819_), .B1(new_n792_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT53), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n823_));
  OAI221_X1 g622(.A(new_n823_), .B1(new_n792_), .B2(new_n820_), .C1(new_n819_), .C2(new_n818_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(G1339gat));
  NAND4_X1  g624(.A1(new_n713_), .A2(new_n654_), .A3(new_n640_), .A4(new_n506_), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(KEYINPUT54), .Z(new_n827_));
  INV_X1    g626(.A(new_n640_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n560_), .A2(new_n587_), .A3(new_n586_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n588_), .B1(KEYINPUT12), .B2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n570_), .B1(new_n549_), .B2(new_n560_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n585_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n585_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(KEYINPUT55), .B2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n572_), .A2(new_n583_), .A3(KEYINPUT55), .A4(new_n573_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n595_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT56), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n573_), .B1(new_n572_), .B2(new_n583_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n584_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n596_), .B1(new_n841_), .B2(new_n835_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n497_), .A2(new_n498_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n845_), .A2(KEYINPUT114), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(KEYINPUT114), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n468_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n489_), .A2(new_n492_), .A3(new_n469_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n503_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n493_), .A2(new_n499_), .A3(new_n467_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n850_), .A2(new_n601_), .A3(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n838_), .A2(new_n844_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(KEYINPUT116), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(KEYINPUT116), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n838_), .A2(new_n856_), .A3(new_n844_), .A4(new_n852_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n828_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n837_), .A2(new_n860_), .A3(KEYINPUT56), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n843_), .B1(new_n842_), .B2(KEYINPUT113), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n505_), .A2(new_n601_), .A3(KEYINPUT112), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT112), .B1(new_n505_), .B2(new_n601_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n861_), .A2(new_n862_), .A3(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n597_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n628_), .A2(new_n629_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n869_), .A2(new_n631_), .A3(new_n609_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT57), .B1(new_n870_), .B2(new_n660_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n859_), .B1(new_n868_), .B2(new_n872_), .ZN(new_n873_));
  AOI211_X1 g672(.A(KEYINPUT117), .B(new_n871_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n661_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(KEYINPUT115), .ZN(new_n877_));
  INV_X1    g676(.A(new_n661_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n868_), .A2(KEYINPUT115), .A3(new_n878_), .ZN(new_n879_));
  OAI221_X1 g678(.A(new_n858_), .B1(new_n873_), .B2(new_n874_), .C1(new_n877_), .C2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n827_), .B1(new_n880_), .B2(new_n653_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n725_), .A2(new_n425_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(new_n448_), .A3(new_n255_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(G113gat), .B1(new_n884_), .B2(new_n505_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n877_), .A2(new_n879_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n858_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n653_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n826_), .B(KEYINPUT54), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n883_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT59), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894_));
  AOI211_X1 g693(.A(new_n894_), .B(new_n883_), .C1(new_n889_), .C2(new_n890_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n886_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n891_), .A2(KEYINPUT59), .A3(new_n892_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n897_), .A2(KEYINPUT118), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n899_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n505_), .A2(G113gat), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n885_), .B1(new_n900_), .B2(new_n901_), .ZN(G1340gat));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n903_));
  AOI21_X1  g702(.A(G120gat), .B1(new_n603_), .B2(new_n903_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(KEYINPUT119), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n903_), .B2(G120gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n891_), .A2(new_n892_), .A3(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT120), .ZN(new_n908_));
  INV_X1    g707(.A(G120gat), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n604_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(G1341gat));
  AOI21_X1  g710(.A(G127gat), .B1(new_n884_), .B2(new_n654_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n654_), .A2(G127gat), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n900_), .B2(new_n913_), .ZN(G1342gat));
  AOI21_X1  g713(.A(G134gat), .B1(new_n884_), .B2(new_n662_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n828_), .A2(G134gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n900_), .B2(new_n916_), .ZN(G1343gat));
  NOR4_X1   g716(.A1(new_n725_), .A2(new_n447_), .A3(new_n255_), .A4(new_n451_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n891_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n506_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(new_n336_), .ZN(G1344gat));
  NOR2_X1   g720(.A1(new_n919_), .A2(new_n604_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(new_n337_), .ZN(G1345gat));
  XNOR2_X1  g722(.A(KEYINPUT61), .B(G155gat), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n891_), .A2(new_n654_), .A3(new_n918_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT121), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n926_), .A2(KEYINPUT121), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n925_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n930_));
  OR2_X1    g729(.A1(new_n926_), .A2(KEYINPUT121), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n931_), .A2(new_n927_), .A3(new_n924_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1346gat));
  NAND4_X1  g732(.A1(new_n891_), .A2(G162gat), .A3(new_n704_), .A4(new_n918_), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n891_), .A2(new_n662_), .A3(new_n918_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n935_), .B2(G162gat), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  OAI211_X1 g737(.A(KEYINPUT122), .B(new_n934_), .C1(new_n935_), .C2(G162gat), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1347gat));
  NAND2_X1  g739(.A1(new_n725_), .A2(new_n449_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n690_), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n891_), .A2(new_n209_), .A3(new_n505_), .A4(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(KEYINPUT62), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(G169gat), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n891_), .A2(new_n942_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n946_), .A2(KEYINPUT62), .A3(new_n506_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n212_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n945_), .B1(new_n948_), .B2(new_n944_), .ZN(G1348gat));
  OAI21_X1  g748(.A(new_n210_), .B1(new_n946_), .B2(new_n713_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  OAI211_X1 g751(.A(KEYINPUT123), .B(new_n210_), .C1(new_n946_), .C2(new_n713_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n954_), .B1(new_n881_), .B2(new_n425_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n941_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n891_), .A2(KEYINPUT124), .A3(new_n451_), .ZN(new_n957_));
  AND3_X1   g756(.A1(new_n955_), .A2(new_n956_), .A3(new_n957_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n604_), .A2(new_n210_), .ZN(new_n959_));
  AOI22_X1  g758(.A1(new_n952_), .A2(new_n953_), .B1(new_n958_), .B2(new_n959_), .ZN(G1349gat));
  NOR3_X1   g759(.A1(new_n946_), .A2(new_n216_), .A3(new_n653_), .ZN(new_n961_));
  NAND4_X1  g760(.A1(new_n955_), .A2(new_n654_), .A3(new_n956_), .A4(new_n957_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n961_), .B1(new_n962_), .B2(new_n203_), .ZN(G1350gat));
  OAI21_X1  g762(.A(G190gat), .B1(new_n946_), .B2(new_n640_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n662_), .A2(new_n219_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n964_), .B1(new_n946_), .B2(new_n965_), .ZN(G1351gat));
  NAND3_X1  g765(.A1(new_n725_), .A2(new_n256_), .A3(new_n454_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n881_), .A2(new_n967_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(new_n505_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g769(.A1(new_n968_), .A2(new_n605_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n266_), .A2(KEYINPUT125), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n971_), .B(new_n972_), .ZN(G1353gat));
  AOI21_X1  g772(.A(new_n653_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(KEYINPUT126), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n968_), .A2(new_n975_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n977_));
  XOR2_X1   g776(.A(new_n976_), .B(new_n977_), .Z(G1354gat));
  INV_X1    g777(.A(G218gat), .ZN(new_n979_));
  NAND3_X1  g778(.A1(new_n968_), .A2(new_n979_), .A3(new_n662_), .ZN(new_n980_));
  NOR3_X1   g779(.A1(new_n881_), .A2(new_n640_), .A3(new_n967_), .ZN(new_n981_));
  OAI21_X1  g780(.A(new_n980_), .B1(new_n981_), .B2(new_n979_), .ZN(G1355gat));
endmodule


