//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT73), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n202_), .A2(KEYINPUT73), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n202_), .A2(KEYINPUT73), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(new_n208_), .A3(new_n204_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211_));
  INV_X1    g010(.A(G1gat), .ZN(new_n212_));
  INV_X1    g011(.A(G8gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G1gat), .B(G8gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n210_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT80), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n210_), .B(KEYINPUT15), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n217_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G229gat), .A2(G233gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n210_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n217_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n220_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT81), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n223_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n225_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G141gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G169gat), .B(G197gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT83), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT83), .B1(new_n232_), .B2(new_n235_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n232_), .A2(KEYINPUT82), .ZN(new_n241_));
  INV_X1    g040(.A(new_n235_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n232_), .B2(KEYINPUT82), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G230gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G99gat), .A2(G106gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT6), .ZN(new_n251_));
  INV_X1    g050(.A(G99gat), .ZN(new_n252_));
  INV_X1    g051(.A(G106gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(KEYINPUT68), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT7), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT7), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n256_), .A2(new_n252_), .A3(new_n253_), .A4(KEYINPUT68), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n251_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(G92gat), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n259_), .A2(G85gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(G85gat), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT69), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT8), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT10), .B(G99gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT66), .B(G85gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT9), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n259_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n268_), .B1(KEYINPUT9), .B2(G85gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n270_), .B(KEYINPUT67), .Z(new_n271_));
  OAI221_X1 g070(.A(new_n251_), .B1(G106gat), .B2(new_n265_), .C1(new_n269_), .C2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n264_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G57gat), .B(G64gat), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(KEYINPUT11), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT11), .ZN(new_n276_));
  XOR2_X1   g075(.A(G71gat), .B(G78gat), .Z(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n276_), .A2(new_n277_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n273_), .A2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n282_), .A2(KEYINPUT12), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n264_), .A2(new_n272_), .A3(new_n280_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(KEYINPUT12), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n249_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n249_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G120gat), .B(G148gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(G176gat), .B(G204gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n289_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT13), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n296_), .A2(KEYINPUT71), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(KEYINPUT71), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n295_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n295_), .A2(new_n298_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT72), .ZN(new_n302_));
  OR3_X1    g101(.A1(new_n299_), .A2(new_n300_), .A3(KEYINPUT72), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G231gat), .A2(G233gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n217_), .B(new_n305_), .Z(new_n306_));
  OR2_X1    g105(.A1(new_n306_), .A2(new_n280_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n280_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT77), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G127gat), .B(G155gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT16), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G183gat), .B(G211gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n314_), .B(KEYINPUT17), .Z(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT78), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n309_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n307_), .A2(KEYINPUT75), .A3(new_n308_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n314_), .A2(KEYINPUT17), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n321_), .B(KEYINPUT76), .Z(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT79), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n221_), .A2(new_n273_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G232gat), .A2(G233gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT34), .ZN(new_n330_));
  OAI221_X1 g129(.A(new_n328_), .B1(KEYINPUT35), .B2(new_n330_), .C1(new_n226_), .C2(new_n273_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(KEYINPUT35), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G190gat), .B(G218gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G134gat), .B(G162gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n336_), .A2(KEYINPUT36), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n333_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n336_), .B(KEYINPUT36), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n333_), .A2(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT26), .ZN(new_n343_));
  OR3_X1    g142(.A1(new_n343_), .A2(KEYINPUT84), .A3(G190gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT25), .B(G183gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT84), .B1(new_n343_), .B2(G190gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(G190gat), .B1(KEYINPUT85), .B2(KEYINPUT26), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(KEYINPUT85), .B2(KEYINPUT26), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT23), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(G183gat), .A3(G190gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT86), .B1(G169gat), .B2(G176gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NOR3_X1   g158(.A1(KEYINPUT86), .A2(G169gat), .A3(G176gat), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(KEYINPUT24), .A3(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n361_), .A2(KEYINPUT24), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n350_), .A2(new_n357_), .A3(new_n363_), .A4(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(new_n352_), .B2(new_n356_), .ZN(new_n367_));
  INV_X1    g166(.A(G169gat), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n368_), .A2(KEYINPUT22), .ZN(new_n369_));
  INV_X1    g168(.A(G176gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(KEYINPUT22), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n362_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT88), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n367_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(KEYINPUT88), .A3(new_n362_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n365_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G15gat), .B(G43gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT89), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT30), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n378_), .B(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G227gat), .A2(G233gat), .ZN(new_n383_));
  INV_X1    g182(.A(G71gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n382_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G127gat), .B(G134gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT90), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G113gat), .B(G120gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT31), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(new_n252_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n386_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G22gat), .B(G50gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G155gat), .A2(G162gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT92), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT92), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n403_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(G141gat), .A2(G148gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT2), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n409_), .B1(G141gat), .B2(G148gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G141gat), .A2(G148gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n411_), .A2(KEYINPUT2), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n408_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT93), .B1(new_n405_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(KEYINPUT2), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(G141gat), .A3(G148gat), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n415_), .A2(new_n416_), .B1(new_n407_), .B2(new_n406_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n402_), .A2(new_n404_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT93), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n400_), .B1(new_n414_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n406_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n411_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n396_), .B1(new_n398_), .B2(KEYINPUT1), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n424_), .A2(KEYINPUT91), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n396_), .A2(KEYINPUT1), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n424_), .B2(KEYINPUT91), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n423_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT94), .B1(new_n421_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n420_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n419_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n399_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n428_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT94), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n429_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT28), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n437_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n395_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(new_n439_), .A3(new_n394_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n444_), .A3(KEYINPUT99), .ZN(new_n445_));
  AND2_X1   g244(.A1(KEYINPUT95), .A2(G197gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(KEYINPUT95), .A2(G197gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(G204gat), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OR2_X1    g247(.A1(G197gat), .A2(G204gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT21), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OR3_X1    g251(.A1(new_n446_), .A2(new_n447_), .A3(G204gat), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n451_), .B1(G197gat), .B2(G204gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G211gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n456_), .A2(G218gat), .ZN(new_n457_));
  INV_X1    g256(.A(G218gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n458_), .A2(G211gat), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT96), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(G211gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(G218gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT96), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n452_), .A2(new_n455_), .A3(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n460_), .A2(KEYINPUT21), .A3(new_n464_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT97), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n448_), .A2(new_n468_), .A3(new_n449_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT98), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n471_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT98), .ZN(new_n474_));
  NOR4_X1   g273(.A1(new_n473_), .A2(new_n467_), .A3(new_n469_), .A4(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n466_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n414_), .A2(new_n420_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n428_), .B1(new_n477_), .B2(new_n399_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n476_), .B1(new_n438_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(G228gat), .A3(G233gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G228gat), .A2(G233gat), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n481_), .B(new_n476_), .C1(new_n436_), .C2(new_n438_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G78gat), .B(G106gat), .Z(new_n484_));
  AND2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n483_), .A2(new_n484_), .ZN(new_n486_));
  OR3_X1    g285(.A1(new_n445_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n483_), .B(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n442_), .A2(new_n444_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT99), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n488_), .A2(new_n491_), .A3(new_n445_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G8gat), .B(G36gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT18), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G64gat), .B(G92gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n496_), .B(new_n497_), .Z(new_n498_));
  AND2_X1   g297(.A1(new_n498_), .A2(KEYINPUT32), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n365_), .A2(new_n377_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT20), .B1(new_n476_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G226gat), .A2(G233gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT19), .ZN(new_n503_));
  INV_X1    g302(.A(new_n466_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n450_), .A2(KEYINPUT97), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n463_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n505_), .A2(new_n508_), .A3(new_n471_), .A4(KEYINPUT21), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n474_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n470_), .A2(KEYINPUT98), .A3(new_n471_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n504_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n366_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n373_), .B1(new_n357_), .B2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT26), .B(G190gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n345_), .A2(new_n515_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n356_), .B2(new_n352_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n363_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n514_), .A2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n512_), .A2(new_n520_), .ZN(new_n521_));
  NOR3_X1   g320(.A1(new_n501_), .A2(new_n503_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n503_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT20), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n524_), .B1(new_n512_), .B2(new_n520_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n476_), .A2(new_n500_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n523_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n499_), .B1(new_n522_), .B2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n503_), .B1(new_n501_), .B2(new_n521_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n525_), .A2(new_n523_), .A3(new_n526_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n528_), .B1(new_n531_), .B2(new_n499_), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n388_), .B(new_n389_), .Z(new_n533_));
  NAND3_X1  g332(.A1(new_n429_), .A2(new_n435_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT101), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n535_), .B1(new_n478_), .B2(new_n390_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n429_), .A2(new_n435_), .A3(new_n533_), .A4(new_n535_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT4), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT4), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n429_), .A2(new_n435_), .A3(new_n533_), .A4(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G225gat), .A2(G233gat), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n540_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n539_), .A2(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(G1gat), .B(G29gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(G57gat), .B(G85gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n539_), .B2(new_n543_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n547_), .A2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n532_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n498_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n525_), .A2(new_n523_), .A3(new_n526_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n524_), .B1(new_n512_), .B2(new_n378_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n520_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n476_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n523_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n559_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n529_), .A2(new_n498_), .A3(new_n530_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(KEYINPUT100), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT100), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n531_), .A2(new_n568_), .A3(new_n559_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n540_), .A2(KEYINPUT103), .A3(new_n543_), .A4(new_n542_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT103), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n541_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n542_), .A2(new_n543_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n554_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n576_), .B1(new_n539_), .B2(new_n544_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n571_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n547_), .B2(new_n556_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n548_), .A2(new_n576_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n545_), .B1(new_n539_), .B2(KEYINPUT4), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n581_), .A2(KEYINPUT33), .A3(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n570_), .B(new_n578_), .C1(new_n580_), .C2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n558_), .B1(new_n584_), .B2(KEYINPUT104), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n557_), .A2(KEYINPUT33), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n547_), .A2(new_n579_), .A3(new_n556_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT104), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(new_n570_), .A4(new_n578_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n494_), .B1(new_n585_), .B2(new_n590_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n549_), .A2(new_n554_), .B1(new_n547_), .B2(new_n556_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n487_), .A2(new_n492_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT105), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n566_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n566_), .A2(new_n594_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n559_), .B1(new_n522_), .B2(new_n527_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n595_), .A2(KEYINPUT27), .A3(new_n596_), .A4(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT27), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n567_), .A2(new_n599_), .A3(new_n569_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n593_), .A2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n393_), .B1(new_n591_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n592_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(new_n393_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n601_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n493_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n342_), .B1(new_n603_), .B2(new_n607_), .ZN(new_n608_));
  AND4_X1   g407(.A1(new_n246_), .A2(new_n304_), .A3(new_n327_), .A4(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n609_), .A2(new_n604_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n212_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n245_), .B1(new_n603_), .B2(new_n607_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n341_), .B(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n326_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n304_), .A2(new_n612_), .A3(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT106), .Z(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n212_), .A3(new_n604_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT38), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n611_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n620_), .B2(new_n619_), .ZN(G1324gat));
  AOI21_X1  g421(.A(new_n213_), .B1(new_n609_), .B2(new_n601_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT39), .Z(new_n624_));
  NAND3_X1  g423(.A1(new_n618_), .A2(new_n213_), .A3(new_n601_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g426(.A(new_n393_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n609_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(G15gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT41), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n617_), .A2(G15gat), .A3(new_n393_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1326gat));
  NAND2_X1  g432(.A1(new_n609_), .A2(new_n494_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(G22gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT42), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n493_), .A2(G22gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n636_), .B1(new_n617_), .B2(new_n637_), .ZN(G1327gat));
  NAND2_X1  g437(.A1(new_n302_), .A2(new_n303_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT108), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(new_n327_), .B2(new_n341_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n326_), .A2(KEYINPUT108), .A3(new_n342_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n639_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n612_), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n644_), .A2(G29gat), .A3(new_n592_), .ZN(new_n645_));
  AND4_X1   g444(.A1(new_n246_), .A2(new_n302_), .A3(new_n303_), .A4(new_n326_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n341_), .B(new_n613_), .ZN(new_n647_));
  AOI211_X1 g446(.A(KEYINPUT43), .B(new_n647_), .C1(new_n603_), .C2(new_n607_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n570_), .A2(new_n578_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n583_), .A2(new_n580_), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT104), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n558_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n590_), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n602_), .B1(new_n654_), .B2(new_n493_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n607_), .B1(new_n655_), .B2(new_n628_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n649_), .B1(new_n656_), .B2(new_n615_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n646_), .B1(new_n648_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n646_), .B(KEYINPUT44), .C1(new_n648_), .C2(new_n657_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n604_), .A3(new_n661_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n662_), .A2(KEYINPUT107), .A3(G29gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT107), .B1(new_n662_), .B2(G29gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n645_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT109), .Z(G1328gat));
  XNOR2_X1  g465(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT111), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n660_), .A2(new_n601_), .A3(new_n661_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(KEYINPUT110), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n660_), .A2(new_n671_), .A3(new_n601_), .A4(new_n661_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G36gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n668_), .B1(new_n670_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n669_), .A2(KEYINPUT110), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n675_), .A2(KEYINPUT111), .A3(G36gat), .A4(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n606_), .A2(G36gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n643_), .A2(new_n612_), .A3(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT45), .Z(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n667_), .B1(new_n677_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n667_), .ZN(new_n683_));
  AOI211_X1 g482(.A(new_n680_), .B(new_n683_), .C1(new_n674_), .C2(new_n676_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1329gat));
  NAND4_X1  g484(.A1(new_n660_), .A2(G43gat), .A3(new_n628_), .A4(new_n661_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n644_), .A2(new_n393_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(G43gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n688_), .B2(KEYINPUT113), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(KEYINPUT113), .B2(new_n686_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g490(.A1(new_n660_), .A2(G50gat), .A3(new_n494_), .A4(new_n661_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n644_), .A2(new_n493_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(G50gat), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT114), .ZN(G1331gat));
  NAND2_X1  g494(.A1(new_n656_), .A2(new_n245_), .ZN(new_n696_));
  NOR4_X1   g495(.A1(new_n304_), .A2(new_n696_), .A3(new_n326_), .A4(new_n615_), .ZN(new_n697_));
  INV_X1    g496(.A(G57gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n604_), .ZN(new_n699_));
  AND4_X1   g498(.A1(new_n245_), .A2(new_n608_), .A3(new_n639_), .A4(new_n327_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(new_n604_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n699_), .B1(new_n701_), .B2(new_n698_), .ZN(G1332gat));
  INV_X1    g501(.A(G64gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n700_), .B2(new_n601_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT48), .Z(new_n705_));
  NAND2_X1  g504(.A1(new_n601_), .A2(new_n703_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT115), .Z(new_n707_));
  NAND2_X1  g506(.A1(new_n697_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(G1333gat));
  AOI21_X1  g508(.A(new_n384_), .B1(new_n700_), .B2(new_n628_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT49), .Z(new_n711_));
  NAND3_X1  g510(.A1(new_n697_), .A2(new_n384_), .A3(new_n628_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT116), .Z(G1334gat));
  INV_X1    g513(.A(G78gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n700_), .B2(new_n494_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT50), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n697_), .A2(new_n715_), .A3(new_n494_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1335gat));
  AOI211_X1 g518(.A(new_n696_), .B(new_n304_), .C1(new_n642_), .C2(new_n641_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G85gat), .B1(new_n720_), .B2(new_n604_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n648_), .A2(new_n657_), .ZN(new_n722_));
  NOR4_X1   g521(.A1(new_n722_), .A2(new_n246_), .A3(new_n304_), .A4(new_n327_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n592_), .A2(new_n266_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT117), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n721_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT118), .ZN(G1336gat));
  AOI21_X1  g526(.A(G92gat), .B1(new_n720_), .B2(new_n601_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n601_), .A2(G92gat), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT119), .Z(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n723_), .B2(new_n730_), .ZN(G1337gat));
  AOI21_X1  g530(.A(new_n252_), .B1(new_n723_), .B2(new_n628_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n393_), .A2(new_n265_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n720_), .B2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g534(.A1(new_n720_), .A2(new_n253_), .A3(new_n494_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n723_), .A2(new_n494_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(G106gat), .ZN(new_n739_));
  AOI211_X1 g538(.A(KEYINPUT52), .B(new_n253_), .C1(new_n723_), .C2(new_n494_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g541(.A1(new_n601_), .A2(new_n592_), .A3(new_n393_), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n289_), .A2(new_n294_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n240_), .B2(new_n244_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n283_), .A2(new_n285_), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT120), .B(KEYINPUT55), .C1(new_n746_), .C2(new_n249_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT120), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n286_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT122), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n283_), .A2(new_n249_), .A3(new_n285_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT121), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n751_), .A2(new_n752_), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n752_), .B1(new_n751_), .B2(new_n755_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n294_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT56), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n751_), .A2(new_n755_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT122), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n751_), .A2(new_n752_), .A3(new_n755_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(KEYINPUT56), .A3(new_n294_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n745_), .B1(new_n760_), .B2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n236_), .B(new_n237_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n230_), .A2(new_n223_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n220_), .A2(new_n222_), .A3(new_n231_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n242_), .A3(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n295_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n341_), .B1(new_n766_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n744_), .B(new_n770_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n760_), .B2(new_n765_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n647_), .B1(new_n776_), .B2(KEYINPUT58), .ZN(new_n777_));
  INV_X1    g576(.A(new_n775_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n758_), .A2(new_n759_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT56), .B1(new_n764_), .B2(new_n294_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n773_), .A2(new_n774_), .B1(new_n777_), .B2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT57), .B(new_n341_), .C1(new_n766_), .C2(new_n772_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n327_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n616_), .A2(new_n245_), .A3(new_n301_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n493_), .B(new_n743_), .C1(new_n786_), .C2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(G113gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n246_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n790_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n773_), .A2(new_n774_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n777_), .A2(new_n783_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n785_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n326_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n787_), .B(KEYINPUT54), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n801_), .A2(KEYINPUT59), .A3(new_n493_), .A4(new_n743_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n245_), .B1(new_n795_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n793_), .B1(new_n803_), .B2(new_n792_), .ZN(G1340gat));
  INV_X1    g603(.A(G120gat), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n304_), .B2(KEYINPUT60), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n791_), .B(new_n806_), .C1(KEYINPUT60), .C2(new_n805_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n304_), .B1(new_n795_), .B2(new_n802_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n805_), .ZN(G1341gat));
  INV_X1    g608(.A(G127gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n791_), .A2(new_n810_), .A3(new_n327_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n326_), .B1(new_n795_), .B2(new_n802_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n810_), .ZN(G1342gat));
  INV_X1    g612(.A(G134gat), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n791_), .A2(new_n814_), .A3(new_n342_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n647_), .B1(new_n795_), .B2(new_n802_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(new_n814_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT123), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT123), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n819_), .B(new_n815_), .C1(new_n816_), .C2(new_n814_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(G1343gat));
  NOR3_X1   g620(.A1(new_n493_), .A2(new_n592_), .A3(new_n628_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n801_), .A2(new_n606_), .A3(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(new_n245_), .ZN(new_n824_));
  XOR2_X1   g623(.A(new_n824_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n304_), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g626(.A1(new_n823_), .A2(new_n326_), .ZN(new_n828_));
  XOR2_X1   g627(.A(KEYINPUT61), .B(G155gat), .Z(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(G1346gat));
  OAI21_X1  g629(.A(G162gat), .B1(new_n823_), .B2(new_n647_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n341_), .A2(G162gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n823_), .B2(new_n832_), .ZN(G1347gat));
  NOR2_X1   g632(.A1(new_n786_), .A2(new_n789_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n494_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n605_), .A2(new_n601_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n838_), .A2(new_n371_), .A3(new_n369_), .A4(new_n246_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n246_), .A2(new_n836_), .ZN(new_n840_));
  XOR2_X1   g639(.A(new_n840_), .B(KEYINPUT124), .Z(new_n841_));
  NAND3_X1  g640(.A1(new_n801_), .A2(new_n493_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT125), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n368_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT62), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(KEYINPUT125), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n839_), .B1(new_n848_), .B2(new_n849_), .ZN(G1348gat));
  NOR2_X1   g649(.A1(new_n837_), .A2(new_n304_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(new_n370_), .ZN(G1349gat));
  NOR2_X1   g651(.A1(new_n837_), .A2(new_n326_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n853_), .B(new_n345_), .C1(KEYINPUT126), .C2(G183gat), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT126), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(G183gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n853_), .B2(new_n856_), .ZN(G1350gat));
  OAI21_X1  g656(.A(G190gat), .B1(new_n837_), .B2(new_n647_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n342_), .A2(new_n515_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n837_), .B2(new_n859_), .ZN(G1351gat));
  NOR4_X1   g659(.A1(new_n834_), .A2(new_n593_), .A3(new_n606_), .A4(new_n628_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n246_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n639_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g664(.A1(new_n861_), .A2(new_n327_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT63), .B(G211gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n866_), .B2(new_n869_), .ZN(G1354gat));
  NAND2_X1  g669(.A1(new_n861_), .A2(new_n342_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT127), .B(G218gat), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n647_), .A2(new_n872_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n871_), .A2(new_n872_), .B1(new_n861_), .B2(new_n873_), .ZN(G1355gat));
endmodule


