//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n204_));
  OR3_X1    g003(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT8), .ZN(new_n211_));
  OR3_X1    g010(.A1(new_n210_), .A2(KEYINPUT66), .A3(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT65), .B(KEYINPUT9), .Z(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n214_));
  AOI22_X1  g013(.A1(new_n213_), .A2(new_n209_), .B1(new_n207_), .B2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT10), .B(G99gat), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G106gat), .Z(new_n217_));
  OAI211_X1 g016(.A(new_n215_), .B(new_n203_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n210_), .B1(KEYINPUT66), .B2(new_n211_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n212_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G57gat), .B(G64gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(KEYINPUT11), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G71gat), .B(G78gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(KEYINPUT11), .ZN(new_n225_));
  XOR2_X1   g024(.A(new_n224_), .B(new_n225_), .Z(new_n226_));
  AND2_X1   g025(.A1(new_n220_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT12), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n229_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n227_), .B2(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n220_), .A2(new_n226_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NOR3_X1   g034(.A1(new_n231_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G230gat), .ZN(new_n237_));
  INV_X1    g036(.A(G233gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n239_), .B1(new_n235_), .B2(new_n227_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G120gat), .B(G148gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G204gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT5), .B(G176gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n243_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n241_), .A2(new_n242_), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n247_), .B(KEYINPUT68), .Z(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n252_), .A2(KEYINPUT13), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(KEYINPUT13), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT69), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G15gat), .B(G22gat), .ZN(new_n260_));
  INV_X1    g059(.A(G1gat), .ZN(new_n261_));
  INV_X1    g060(.A(G8gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT14), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G1gat), .B(G8gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n264_), .B(new_n265_), .Z(new_n266_));
  XNOR2_X1  g065(.A(G29gat), .B(G36gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G43gat), .B(G50gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  XNOR2_X1  g068(.A(new_n266_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT72), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G229gat), .A2(G233gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n269_), .B(KEYINPUT15), .Z(new_n274_));
  INV_X1    g073(.A(new_n266_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n269_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n273_), .B1(new_n266_), .B2(new_n277_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n271_), .A2(new_n273_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G113gat), .B(G141gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G169gat), .ZN(new_n281_));
  INV_X1    g080(.A(G197gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n279_), .B(new_n283_), .Z(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n259_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G232gat), .A2(G233gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT34), .ZN(new_n288_));
  OAI22_X1  g087(.A1(new_n220_), .A2(new_n269_), .B1(KEYINPUT35), .B2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n220_), .B2(new_n274_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(KEYINPUT35), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n291_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G190gat), .B(G218gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G134gat), .B(G162gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NOR3_X1   g096(.A1(new_n294_), .A2(KEYINPUT36), .A3(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(KEYINPUT36), .Z(new_n299_));
  AND2_X1   g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(KEYINPUT70), .A3(KEYINPUT37), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT37), .B1(new_n301_), .B2(KEYINPUT70), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G127gat), .B(G155gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT16), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(G183gat), .ZN(new_n309_));
  INV_X1    g108(.A(G211gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n226_), .B(new_n275_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G231gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(new_n314_), .B2(KEYINPUT71), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n311_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n315_), .B1(KEYINPUT17), .B2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(KEYINPUT17), .B2(new_n315_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n306_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321_));
  INV_X1    g120(.A(G183gat), .ZN(new_n322_));
  INV_X1    g121(.A(G190gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n323_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(G176gat), .B1(KEYINPUT73), .B2(KEYINPUT22), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(G169gat), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n324_), .A2(new_n325_), .A3(KEYINPUT74), .A4(new_n326_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n324_), .A2(new_n326_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT25), .B(G183gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT26), .B(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(G169gat), .ZN(new_n338_));
  INV_X1    g137(.A(G176gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(KEYINPUT24), .A3(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n340_), .A2(KEYINPUT24), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n334_), .A2(new_n337_), .A3(new_n342_), .A4(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n333_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT30), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT75), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G71gat), .B(G99gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n346_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G15gat), .B(G43gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT77), .ZN(new_n354_));
  XOR2_X1   g153(.A(G127gat), .B(G134gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(G113gat), .B(G120gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT31), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n354_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT77), .B1(new_n353_), .B2(new_n360_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n358_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n366_));
  INV_X1    g165(.A(G155gat), .ZN(new_n367_));
  INV_X1    g166(.A(G162gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT1), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT78), .B1(G155gat), .B2(G162gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n369_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT79), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n369_), .A2(new_n371_), .A3(new_n375_), .A4(new_n372_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT80), .B1(new_n370_), .B2(KEYINPUT1), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT1), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n378_), .A2(new_n379_), .A3(G155gat), .A4(G162gat), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n374_), .A2(new_n376_), .A3(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G141gat), .B(G148gat), .Z(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n369_), .A2(new_n372_), .A3(new_n370_), .ZN(new_n385_));
  INV_X1    g184(.A(G141gat), .ZN(new_n386_));
  INV_X1    g185(.A(G148gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(KEYINPUT3), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(G141gat), .B2(G148gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n391_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n385_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n384_), .A2(new_n398_), .A3(new_n357_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n357_), .B1(new_n384_), .B2(new_n398_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT4), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT93), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n384_), .A2(new_n398_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n357_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n402_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G225gat), .A2(G233gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT92), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n384_), .A2(new_n398_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n409_), .A2(KEYINPUT93), .A3(new_n404_), .A4(new_n357_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n401_), .A2(new_n406_), .A3(new_n408_), .A4(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT0), .ZN(new_n413_));
  INV_X1    g212(.A(G57gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(G85gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n407_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT94), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  OAI211_X1 g218(.A(KEYINPUT94), .B(new_n407_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n411_), .A2(new_n416_), .A3(new_n419_), .A4(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n419_), .A2(new_n420_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n416_), .B1(new_n422_), .B2(new_n411_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n409_), .A2(KEYINPUT29), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G22gat), .B(G50gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT82), .B(KEYINPUT28), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n425_), .B(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(G204gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G197gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n282_), .A2(G204gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n433_), .A2(KEYINPUT21), .ZN(new_n434_));
  XOR2_X1   g233(.A(G211gat), .B(G218gat), .Z(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OR3_X1    g235(.A1(new_n282_), .A2(KEYINPUT84), .A3(G204gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n431_), .A2(KEYINPUT84), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n432_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT21), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n433_), .A2(KEYINPUT21), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n436_), .A2(new_n440_), .B1(new_n435_), .B2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n409_), .B2(KEYINPUT29), .ZN(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT83), .B(G233gat), .Z(new_n444_));
  AND2_X1   g243(.A1(new_n444_), .A2(G228gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n445_), .B(KEYINPUT85), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n448_), .B1(new_n443_), .B2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G78gat), .B(G106gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n429_), .B1(new_n452_), .B2(KEYINPUT86), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n450_), .B(new_n451_), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n453_), .B(new_n454_), .Z(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n333_), .A2(new_n344_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n457_), .B1(new_n458_), .B2(new_n442_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n344_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n338_), .A2(KEYINPUT22), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT22), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G169gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n463_), .A3(new_n339_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT87), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n341_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n465_), .B1(new_n464_), .B2(new_n341_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n327_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(KEYINPUT88), .B(new_n327_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n460_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n459_), .B1(new_n472_), .B2(new_n442_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G226gat), .A2(G233gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT19), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n442_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n436_), .A2(new_n440_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n441_), .A2(new_n435_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI211_X1 g278(.A(new_n457_), .B(new_n475_), .C1(new_n479_), .C2(new_n345_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n473_), .A2(new_n475_), .B1(new_n476_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G64gat), .B(G92gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G8gat), .B(G36gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT90), .B1(new_n481_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n473_), .A2(new_n475_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n476_), .A2(new_n480_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n489_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT90), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n481_), .A2(new_n493_), .A3(new_n487_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  OR3_X1    g294(.A1(new_n492_), .A2(KEYINPUT27), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n481_), .A2(new_n487_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT101), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n479_), .A2(new_n345_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n442_), .A2(new_n344_), .A3(new_n468_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n475_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT99), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(KEYINPUT99), .A3(new_n475_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n505_), .B(new_n506_), .C1(new_n475_), .C2(new_n473_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n486_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n498_), .A2(KEYINPUT27), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n496_), .A2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n456_), .A2(new_n510_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n365_), .A2(new_n421_), .A3(new_n424_), .A4(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n424_), .A2(new_n421_), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n510_), .A2(new_n455_), .A3(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT91), .B1(new_n492_), .B2(new_n495_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n421_), .A2(KEYINPUT95), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT33), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n421_), .A2(KEYINPUT95), .A3(KEYINPUT33), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n399_), .A2(new_n400_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n416_), .B1(new_n408_), .B2(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n401_), .A2(new_n406_), .A3(new_n407_), .A4(new_n410_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT20), .B1(new_n479_), .B2(new_n345_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n467_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n464_), .A2(new_n465_), .A3(new_n341_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT88), .B1(new_n528_), .B2(new_n327_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n471_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n344_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n525_), .B1(new_n531_), .B2(new_n479_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n475_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n490_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n486_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(new_n497_), .A3(KEYINPUT90), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT91), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n494_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n515_), .A2(new_n520_), .A3(new_n524_), .A4(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT96), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n518_), .A2(new_n519_), .B1(new_n523_), .B2(new_n522_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT96), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n541_), .A2(new_n542_), .A3(new_n538_), .A4(new_n515_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n487_), .A2(KEYINPUT32), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n507_), .A2(KEYINPUT100), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT100), .B1(new_n507_), .B2(new_n544_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  OR3_X1    g346(.A1(new_n534_), .A2(KEYINPUT97), .A3(new_n544_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT97), .B1(new_n534_), .B2(new_n544_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n421_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n548_), .B(new_n549_), .C1(new_n550_), .C2(new_n423_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n540_), .A2(new_n543_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n514_), .B1(new_n554_), .B2(new_n455_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n512_), .B1(new_n555_), .B2(new_n365_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n286_), .A2(new_n320_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT102), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n513_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n424_), .A2(KEYINPUT102), .A3(new_n421_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n558_), .A2(new_n261_), .A3(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT38), .ZN(new_n564_));
  INV_X1    g363(.A(new_n301_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n556_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT103), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n286_), .A2(new_n318_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n513_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n564_), .B1(new_n570_), .B2(new_n261_), .ZN(G1324gat));
  NAND2_X1  g370(.A1(new_n567_), .A2(new_n568_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n510_), .ZN(new_n573_));
  OAI21_X1  g372(.A(G8gat), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT39), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n558_), .A2(new_n262_), .A3(new_n510_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g377(.A(new_n365_), .ZN(new_n579_));
  OAI21_X1  g378(.A(G15gat), .B1(new_n572_), .B2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT41), .Z(new_n581_));
  INV_X1    g380(.A(G15gat), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n558_), .A2(new_n582_), .A3(new_n365_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(G1326gat));
  OAI21_X1  g383(.A(G22gat), .B1(new_n572_), .B2(new_n455_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT42), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n455_), .A2(G22gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT104), .Z(new_n588_));
  NAND2_X1  g387(.A1(new_n558_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(G1327gat));
  NAND3_X1  g389(.A1(new_n259_), .A2(new_n318_), .A3(new_n285_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n557_), .A2(new_n565_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT110), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n592_), .A2(KEYINPUT110), .A3(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(G29gat), .B1(new_n599_), .B2(new_n513_), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT105), .B(new_n512_), .C1(new_n555_), .C2(new_n365_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT106), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n304_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(KEYINPUT106), .A3(new_n302_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n601_), .A2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n552_), .B1(new_n539_), .B2(KEYINPUT96), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n456_), .B1(new_n608_), .B2(new_n543_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n579_), .B1(new_n609_), .B2(new_n514_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT105), .B1(new_n610_), .B2(new_n512_), .ZN(new_n611_));
  OAI21_X1  g410(.A(KEYINPUT43), .B1(new_n607_), .B2(new_n611_), .ZN(new_n612_));
  AOI211_X1 g411(.A(KEYINPUT43), .B(new_n305_), .C1(new_n610_), .C2(new_n512_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n591_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT109), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n615_), .A2(new_n616_), .A3(KEYINPUT44), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n616_), .B1(new_n615_), .B2(KEYINPUT44), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT105), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n556_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n601_), .A3(new_n606_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n613_), .B1(new_n622_), .B2(KEYINPUT43), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT107), .B1(new_n623_), .B2(new_n591_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n612_), .A2(new_n614_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT107), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n626_), .A3(new_n592_), .ZN(new_n627_));
  XOR2_X1   g426(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n628_));
  NAND3_X1  g427(.A1(new_n624_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n619_), .A2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n562_), .A2(G29gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n600_), .B1(new_n630_), .B2(new_n631_), .ZN(G1328gat));
  NOR2_X1   g431(.A1(new_n573_), .A2(G36gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n596_), .A2(new_n597_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT112), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT112), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n596_), .A2(new_n636_), .A3(new_n597_), .A4(new_n633_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(KEYINPUT45), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT45), .B1(new_n635_), .B2(new_n637_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n629_), .B(new_n510_), .C1(new_n618_), .C2(new_n617_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(KEYINPUT111), .A3(G36gat), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT111), .B1(new_n642_), .B2(G36gat), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n641_), .B(KEYINPUT46), .C1(new_n644_), .C2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n635_), .A2(new_n637_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT45), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(new_n638_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n645_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n651_), .B2(new_n643_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n646_), .B1(new_n652_), .B2(new_n653_), .ZN(G1329gat));
  NAND4_X1  g453(.A1(new_n619_), .A2(G43gat), .A3(new_n365_), .A4(new_n629_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n598_), .A2(new_n579_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(G43gat), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g457(.A1(new_n598_), .A2(G50gat), .A3(new_n455_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n629_), .B(new_n456_), .C1(new_n618_), .C2(new_n617_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(KEYINPUT114), .A3(G50gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT114), .B1(new_n660_), .B2(G50gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT115), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT115), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n665_), .B(new_n659_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1331gat));
  INV_X1    g466(.A(new_n259_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(new_n284_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n669_), .A2(new_n557_), .A3(new_n320_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n414_), .A3(new_n562_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n669_), .A2(new_n318_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n567_), .A3(new_n513_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n674_), .B2(new_n414_), .ZN(G1332gat));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n567_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G64gat), .B1(new_n676_), .B2(new_n573_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT48), .ZN(new_n678_));
  INV_X1    g477(.A(G64gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n670_), .A2(new_n679_), .A3(new_n510_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1333gat));
  OAI21_X1  g480(.A(G71gat), .B1(new_n676_), .B2(new_n579_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT49), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n579_), .A2(G71gat), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT116), .Z(new_n685_));
  NAND2_X1  g484(.A1(new_n670_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(G1334gat));
  OAI21_X1  g486(.A(G78gat), .B1(new_n676_), .B2(new_n455_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT50), .ZN(new_n689_));
  INV_X1    g488(.A(G78gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n670_), .A2(new_n690_), .A3(new_n456_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1335gat));
  INV_X1    g491(.A(new_n318_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n669_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n593_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(G85gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n697_), .A3(new_n562_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n694_), .A2(new_n625_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT117), .Z(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(new_n513_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n698_), .B1(new_n701_), .B2(new_n697_), .ZN(G1336gat));
  AOI21_X1  g501(.A(G92gat), .B1(new_n696_), .B2(new_n510_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n510_), .A2(G92gat), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT118), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n703_), .B1(new_n700_), .B2(new_n705_), .ZN(G1337gat));
  NOR3_X1   g505(.A1(new_n695_), .A2(new_n216_), .A3(new_n579_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n699_), .A2(new_n365_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(G99gat), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g509(.A(G106gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n699_), .B2(new_n456_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT52), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n455_), .A2(new_n217_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n695_), .B2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g516(.A1(new_n365_), .A2(new_n511_), .A3(new_n562_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT55), .B1(new_n236_), .B2(new_n240_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(new_n241_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n250_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT56), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n279_), .A2(new_n283_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n271_), .A2(new_n272_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n272_), .B1(new_n266_), .B2(new_n277_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n283_), .B1(new_n276_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n724_), .A2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n243_), .B2(new_n247_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n723_), .A2(KEYINPUT58), .A3(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT120), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT58), .B1(new_n723_), .B2(new_n730_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n302_), .B2(new_n604_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  OR2_X1    g535(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n285_), .B(new_n248_), .C1(new_n721_), .C2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n721_), .A2(new_n737_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n252_), .ZN(new_n740_));
  OAI22_X1  g539(.A1(new_n738_), .A2(new_n739_), .B1(new_n740_), .B2(new_n729_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n565_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT57), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n736_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n318_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n319_), .B(new_n284_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT54), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(KEYINPUT121), .A3(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT121), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n746_), .B(KEYINPUT54), .Z(new_n750_));
  AOI21_X1  g549(.A(new_n693_), .B1(new_n736_), .B2(new_n743_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n718_), .B1(new_n748_), .B2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G113gat), .B1(new_n753_), .B2(new_n285_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n753_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n745_), .A2(new_n747_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n718_), .A2(KEYINPUT59), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n755_), .A2(KEYINPUT59), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n285_), .A2(G113gat), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT122), .Z(new_n760_));
  AOI21_X1  g559(.A(new_n754_), .B1(new_n758_), .B2(new_n760_), .ZN(G1340gat));
  INV_X1    g560(.A(G120gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n259_), .B2(KEYINPUT60), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n753_), .B(new_n763_), .C1(KEYINPUT60), .C2(new_n762_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n756_), .A2(new_n757_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT59), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n668_), .B(new_n765_), .C1(new_n753_), .C2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n768_), .B2(new_n762_), .ZN(G1341gat));
  INV_X1    g568(.A(G127gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n753_), .A2(new_n770_), .A3(new_n693_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n693_), .B(new_n765_), .C1(new_n753_), .C2(new_n766_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n771_), .B1(new_n773_), .B2(new_n770_), .ZN(G1342gat));
  AOI211_X1 g573(.A(new_n565_), .B(new_n718_), .C1(new_n748_), .C2(new_n752_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT123), .B1(new_n775_), .B2(G134gat), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT123), .ZN(new_n777_));
  INV_X1    g576(.A(G134gat), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n777_), .B(new_n778_), .C1(new_n755_), .C2(new_n565_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n305_), .A2(new_n778_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n776_), .A2(new_n779_), .B1(new_n758_), .B2(new_n780_), .ZN(G1343gat));
  AND2_X1   g580(.A1(new_n748_), .A2(new_n752_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n510_), .A2(new_n455_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n562_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n782_), .A2(new_n365_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n285_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(G141gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n386_), .A3(new_n285_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1344gat));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n668_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G148gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n785_), .A2(new_n387_), .A3(new_n668_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1345gat));
  NAND2_X1  g592(.A1(new_n785_), .A2(new_n693_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(KEYINPUT61), .B(G155gat), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n795_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n785_), .A2(new_n693_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1346gat));
  NAND2_X1  g598(.A1(new_n785_), .A2(new_n301_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n368_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n800_), .A2(new_n368_), .B1(new_n785_), .B2(new_n801_), .ZN(G1347gat));
  NOR3_X1   g601(.A1(new_n579_), .A2(new_n573_), .A3(new_n562_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n756_), .A2(new_n455_), .A3(new_n285_), .A4(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT124), .B1(new_n804_), .B2(G169gat), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT62), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n804_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n461_), .A2(new_n463_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n805_), .A2(new_n806_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n812_), .ZN(G1348gat));
  NOR2_X1   g612(.A1(new_n782_), .A2(new_n456_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n668_), .A2(G176gat), .A3(new_n803_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n756_), .A2(new_n455_), .A3(new_n803_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n816_), .A2(new_n259_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n814_), .A2(new_n815_), .B1(new_n817_), .B2(new_n339_), .ZN(G1349gat));
  NAND2_X1  g617(.A1(new_n756_), .A2(new_n455_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n803_), .A2(new_n693_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n819_), .A2(new_n335_), .A3(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n814_), .A2(new_n693_), .A3(new_n803_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n322_), .ZN(G1350gat));
  OAI21_X1  g622(.A(G190gat), .B1(new_n816_), .B2(new_n305_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n301_), .A2(new_n336_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n816_), .B2(new_n825_), .ZN(G1351gat));
  NAND2_X1  g625(.A1(new_n748_), .A2(new_n752_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n573_), .A2(new_n513_), .A3(new_n455_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n827_), .A2(new_n579_), .A3(new_n285_), .A4(new_n828_), .ZN(new_n829_));
  XOR2_X1   g628(.A(KEYINPUT125), .B(G197gat), .Z(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1352gat));
  NOR2_X1   g630(.A1(new_n782_), .A2(new_n365_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n430_), .A2(KEYINPUT126), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n832_), .A2(new_n668_), .A3(new_n828_), .A4(new_n833_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n832_), .A2(new_n668_), .A3(new_n828_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT126), .B(G204gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n835_), .B2(new_n836_), .ZN(G1353gat));
  NAND4_X1  g636(.A1(new_n827_), .A2(new_n579_), .A3(new_n693_), .A4(new_n828_), .ZN(new_n838_));
  AND2_X1   g637(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n840_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT127), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n838_), .A2(KEYINPUT127), .A3(new_n840_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n841_), .B1(new_n844_), .B2(new_n845_), .ZN(G1354gat));
  NAND3_X1  g645(.A1(new_n832_), .A2(new_n306_), .A3(new_n828_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G218gat), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n565_), .A2(G218gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n832_), .A2(new_n828_), .A3(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(G1355gat));
endmodule


