//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n909_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_;
  XOR2_X1   g000(.A(G127gat), .B(G155gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G183gat), .B(G211gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT17), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n206_), .A2(KEYINPUT17), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G57gat), .B(G64gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT11), .ZN(new_n210_));
  XOR2_X1   g009(.A(G71gat), .B(G78gat), .Z(new_n211_));
  OR2_X1    g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n209_), .A2(KEYINPUT11), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n211_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(G231gat), .A2(G233gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT77), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219_));
  INV_X1    g018(.A(G1gat), .ZN(new_n220_));
  INV_X1    g019(.A(G8gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT14), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G1gat), .B(G8gat), .ZN(new_n224_));
  XOR2_X1   g023(.A(new_n223_), .B(new_n224_), .Z(new_n225_));
  XNOR2_X1  g024(.A(new_n218_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT80), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n225_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n218_), .B(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(KEYINPUT80), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n207_), .B(new_n208_), .C1(new_n228_), .C2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT81), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n207_), .B(KEYINPUT79), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n226_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n232_), .A2(new_n233_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G230gat), .A2(G233gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT64), .Z(new_n241_));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G99gat), .A2(G106gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT6), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT6), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(G99gat), .A3(G106gat), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT7), .ZN(new_n248_));
  INV_X1    g047(.A(G99gat), .ZN(new_n249_));
  INV_X1    g048(.A(G106gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n242_), .B1(new_n247_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n244_), .A2(new_n246_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n255_), .A2(KEYINPUT68), .A3(new_n252_), .A4(new_n251_), .ZN(new_n256_));
  INV_X1    g055(.A(G85gat), .ZN(new_n257_));
  INV_X1    g056(.A(G92gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G85gat), .A2(G92gat), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n259_), .A2(KEYINPUT8), .A3(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n254_), .A2(new_n256_), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT69), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n254_), .A2(new_n264_), .A3(new_n256_), .A4(new_n261_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT8), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n255_), .A2(new_n252_), .A3(new_n251_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n259_), .A2(new_n260_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n266_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n263_), .A2(new_n265_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n257_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n258_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n272_), .B1(new_n276_), .B2(KEYINPUT9), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT9), .ZN(new_n278_));
  AND2_X1   g077(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  OAI211_X1 g080(.A(KEYINPUT67), .B(new_n278_), .C1(new_n281_), .C2(new_n258_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n260_), .B1(new_n259_), .B2(KEYINPUT9), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n277_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(KEYINPUT65), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT65), .ZN(new_n289_));
  INV_X1    g088(.A(new_n287_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n289_), .B1(new_n290_), .B2(new_n285_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n247_), .B1(new_n292_), .B2(new_n250_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n284_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n271_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n215_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT70), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n271_), .A2(new_n295_), .A3(new_n215_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n241_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(new_n301_), .B2(new_n299_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT12), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n269_), .B1(new_n262_), .B2(KEYINPUT69), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n294_), .B1(new_n305_), .B2(new_n265_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n304_), .B1(new_n306_), .B2(new_n215_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n298_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n296_), .A2(new_n304_), .A3(new_n297_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n241_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G120gat), .B(G148gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(G176gat), .B(G204gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  OR3_X1    g115(.A1(new_n303_), .A2(new_n310_), .A3(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n316_), .B1(new_n303_), .B2(new_n310_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n317_), .A2(KEYINPUT13), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT13), .B1(new_n317_), .B2(new_n318_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G113gat), .B(G141gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT84), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G169gat), .B(G197gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G29gat), .B(G36gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G43gat), .B(G50gat), .Z(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G43gat), .B(G50gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n330_), .A2(new_n334_), .A3(new_n332_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(new_n225_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G229gat), .A2(G233gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n342_), .A2(KEYINPUT82), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT82), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n338_), .A2(new_n225_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n340_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT15), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n330_), .A2(new_n334_), .A3(new_n332_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n334_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n349_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n336_), .A2(KEYINPUT15), .A3(new_n337_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(KEYINPUT83), .A3(new_n229_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT83), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n353_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n356_), .B1(new_n357_), .B2(new_n225_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n348_), .B1(new_n355_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n326_), .B1(new_n346_), .B2(new_n359_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n346_), .A2(new_n359_), .A3(new_n326_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT85), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NOR4_X1   g162(.A1(new_n346_), .A2(new_n359_), .A3(KEYINPUT85), .A4(new_n326_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n360_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n239_), .A2(new_n321_), .A3(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT102), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G227gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(G71gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(new_n249_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G15gat), .B(G43gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT88), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n371_), .B(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT23), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT23), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(G183gat), .A3(G190gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(G183gat), .B2(G190gat), .ZN(new_n380_));
  NOR2_X1   g179(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(G169gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT86), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT86), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n386_), .B1(G169gat), .B2(G176gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT24), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n385_), .A2(new_n387_), .A3(KEYINPUT24), .A4(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT25), .B(G183gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT26), .B(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n390_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n378_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT87), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n376_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n375_), .A2(KEYINPUT87), .A3(KEYINPUT23), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n397_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n383_), .B1(new_n396_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT89), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n374_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n404_), .B(new_n405_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n407_), .B2(new_n374_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G127gat), .B(G134gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G113gat), .B(G120gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n411_), .B(KEYINPUT31), .Z(new_n412_));
  OR2_X1    g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n374_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n406_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n412_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT92), .ZN(new_n423_));
  INV_X1    g222(.A(G204gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n423_), .B1(new_n424_), .B2(G197gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(G197gat), .ZN(new_n426_));
  INV_X1    g225(.A(G197gat), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n429_), .A2(KEYINPUT21), .ZN(new_n430_));
  XOR2_X1   g229(.A(G211gat), .B(G218gat), .Z(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(G204gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n426_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n431_), .B1(KEYINPUT21), .B2(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n431_), .A2(KEYINPUT21), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n430_), .A2(new_n434_), .B1(new_n435_), .B2(new_n429_), .ZN(new_n436_));
  INV_X1    g235(.A(G176gat), .ZN(new_n437_));
  INV_X1    g236(.A(G169gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT22), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT22), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(G169gat), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n439_), .A2(new_n441_), .A3(KEYINPUT97), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT97), .B1(new_n439_), .B2(new_n441_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n437_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G183gat), .A2(G190gat), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n444_), .B(new_n391_), .C1(new_n401_), .C2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n390_), .A2(new_n395_), .A3(new_n392_), .A4(new_n379_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n436_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT20), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT101), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(KEYINPUT101), .A3(KEYINPUT20), .ZN(new_n452_));
  INV_X1    g251(.A(new_n436_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n402_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n451_), .A2(new_n452_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G226gat), .A2(G233gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT19), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n446_), .A2(new_n447_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n460_), .B2(new_n453_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n457_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n436_), .B(new_n383_), .C1(new_n396_), .C2(new_n401_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n422_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n457_), .B1(new_n453_), .B2(new_n402_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(KEYINPUT20), .A3(new_n448_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n461_), .A2(new_n463_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n422_), .B(new_n467_), .C1(new_n468_), .C2(new_n462_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT27), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n465_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n422_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n466_), .A2(new_n448_), .A3(KEYINPUT20), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n462_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT27), .B1(new_n469_), .B2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G1gat), .B(G29gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(G85gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT0), .B(G57gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G225gat), .A2(G233gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  OR2_X1    g282(.A1(G155gat), .A2(G162gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G155gat), .A2(G162gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(KEYINPUT90), .A2(G155gat), .A3(G162gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G141gat), .A2(G148gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT3), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G141gat), .A2(G148gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT91), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n492_), .B(new_n493_), .C1(new_n496_), .C2(KEYINPUT2), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n496_), .A2(KEYINPUT2), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n484_), .B(new_n489_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(KEYINPUT90), .A2(G155gat), .A3(G162gat), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT90), .B1(G155gat), .B2(G162gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT1), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT1), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n487_), .A2(new_n503_), .A3(new_n488_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n504_), .A3(new_n484_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G141gat), .B(G148gat), .Z(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n499_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n411_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n483_), .B1(new_n510_), .B2(KEYINPUT4), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n499_), .A2(new_n507_), .A3(new_n411_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n411_), .B1(new_n499_), .B2(new_n507_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT99), .B1(new_n515_), .B2(KEYINPUT4), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n499_), .A2(new_n507_), .A3(new_n411_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n510_), .A2(KEYINPUT99), .A3(KEYINPUT4), .A4(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT100), .B(new_n512_), .C1(new_n516_), .C2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n482_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n510_), .A2(KEYINPUT4), .A3(new_n517_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT99), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n511_), .B1(new_n525_), .B2(new_n518_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(KEYINPUT100), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n481_), .B1(new_n522_), .B2(new_n527_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n526_), .A2(KEYINPUT100), .B1(new_n515_), .B2(new_n482_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n512_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT100), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n481_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n528_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT29), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n499_), .B2(new_n507_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n538_), .A2(new_n436_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G228gat), .A2(G233gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(G228gat), .B(G233gat), .C1(new_n538_), .C2(new_n436_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G78gat), .B(G106gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT28), .B1(new_n508_), .B2(KEYINPUT29), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT28), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n499_), .A2(new_n507_), .A3(new_n548_), .A4(new_n537_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G22gat), .B(G50gat), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n547_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n545_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n541_), .A2(new_n542_), .A3(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n546_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n544_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT96), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n553_), .A2(new_n555_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n543_), .A2(new_n545_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT95), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT96), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n559_), .A2(new_n561_), .A3(new_n562_), .A4(new_n546_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT94), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n543_), .A2(KEYINPUT94), .A3(new_n545_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n555_), .A2(KEYINPUT93), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n541_), .A2(new_n568_), .A3(new_n542_), .A4(new_n554_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .A4(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n553_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n558_), .A2(new_n563_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  AND4_X1   g371(.A1(new_n417_), .A2(new_n477_), .A3(new_n536_), .A4(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n558_), .A2(new_n563_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n571_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(new_n536_), .A3(new_n477_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n482_), .B1(new_n510_), .B2(KEYINPUT4), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n578_), .B1(new_n525_), .B2(new_n518_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n515_), .A2(new_n483_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n481_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n469_), .B(new_n475_), .C1(new_n579_), .C2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT33), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n582_), .B1(new_n534_), .B2(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n529_), .A2(new_n532_), .A3(KEYINPUT33), .A4(new_n533_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n422_), .A2(KEYINPUT32), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n473_), .A2(new_n474_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n458_), .A2(new_n464_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n587_), .B1(new_n588_), .B2(new_n586_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n584_), .A2(new_n585_), .B1(new_n535_), .B2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n577_), .B1(new_n590_), .B2(new_n576_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n417_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n573_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n271_), .A2(new_n338_), .A3(new_n295_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT76), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n598_), .B(new_n599_), .C1(new_n357_), .C2(new_n306_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT74), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n597_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT35), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT76), .B1(new_n296_), .B2(new_n354_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n605_), .A2(KEYINPUT74), .A3(new_n598_), .A4(new_n596_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n602_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT75), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n609_), .A2(KEYINPUT36), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n607_), .A2(new_n612_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT36), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n612_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n593_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n367_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G1gat), .B1(new_n622_), .B2(new_n536_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n619_), .A2(KEYINPUT37), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT36), .B1(new_n607_), .B2(new_n612_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n606_), .A2(new_n604_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT75), .B1(new_n626_), .B2(new_n602_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n625_), .B1(new_n627_), .B2(new_n612_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT37), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n614_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n624_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n239_), .A2(new_n321_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n365_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n632_), .A2(new_n633_), .A3(new_n593_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n220_), .A3(new_n535_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT38), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n636_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n623_), .A2(new_n637_), .A3(new_n638_), .ZN(G1324gat));
  AND2_X1   g438(.A1(new_n469_), .A2(new_n475_), .ZN(new_n640_));
  OAI22_X1  g439(.A1(new_n640_), .A2(KEYINPUT27), .B1(new_n465_), .B2(new_n470_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n634_), .A2(new_n221_), .A3(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G8gat), .B1(new_n622_), .B2(new_n477_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(KEYINPUT39), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(KEYINPUT39), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n642_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT40), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI211_X1 g447(.A(KEYINPUT40), .B(new_n642_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1325gat));
  OAI21_X1  g449(.A(G15gat), .B1(new_n622_), .B2(new_n592_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT41), .Z(new_n652_));
  INV_X1    g451(.A(G15gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n634_), .A2(new_n653_), .A3(new_n417_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(G1326gat));
  NOR2_X1   g454(.A1(new_n572_), .A2(G22gat), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT103), .Z(new_n657_));
  NAND2_X1  g456(.A1(new_n634_), .A2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G22gat), .B1(new_n622_), .B2(new_n572_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(KEYINPUT42), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(KEYINPUT42), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(KEYINPUT104), .B(new_n658_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1327gat));
  INV_X1    g465(.A(new_n321_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n239_), .A2(new_n667_), .A3(new_n619_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n593_), .A2(new_n633_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n671_), .A2(G29gat), .A3(new_n536_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n624_), .A2(new_n674_), .A3(new_n630_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n593_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n534_), .A2(new_n583_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n582_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n585_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n535_), .A2(new_n589_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n576_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n572_), .A2(new_n641_), .A3(new_n535_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n592_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n573_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n628_), .A2(new_n629_), .A3(new_n614_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n629_), .B1(new_n628_), .B2(new_n614_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n686_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT105), .B1(new_n624_), .B2(new_n630_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n685_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n676_), .B1(new_n691_), .B2(KEYINPUT43), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n237_), .A2(new_n238_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(new_n365_), .A3(new_n321_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n673_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n239_), .A2(new_n667_), .A3(new_n633_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n688_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n624_), .A2(KEYINPUT105), .A3(new_n630_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n674_), .B1(new_n700_), .B2(new_n685_), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT106), .B(new_n697_), .C1(new_n701_), .C2(new_n676_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n695_), .A2(new_n696_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n691_), .A2(KEYINPUT43), .ZN(new_n704_));
  INV_X1    g503(.A(new_n676_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n694_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT44), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n703_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708_), .B2(new_n536_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT107), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT107), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n672_), .B1(new_n710_), .B2(new_n711_), .ZN(G1328gat));
  INV_X1    g511(.A(G36gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n670_), .A2(new_n713_), .A3(new_n641_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n477_), .B1(new_n706_), .B2(KEYINPUT44), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n703_), .A2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n719_), .B2(G36gat), .ZN(new_n720_));
  AOI211_X1 g519(.A(KEYINPUT108), .B(new_n713_), .C1(new_n703_), .C2(new_n718_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n716_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(KEYINPUT46), .B(new_n716_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1329gat));
  OAI21_X1  g525(.A(G43gat), .B1(new_n708_), .B2(new_n592_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n671_), .A2(G43gat), .A3(new_n592_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n730_), .B(new_n732_), .ZN(G1330gat));
  AOI21_X1  g532(.A(G50gat), .B1(new_n670_), .B2(new_n576_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n708_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n576_), .A2(G50gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(G1331gat));
  NAND4_X1  g536(.A1(new_n621_), .A2(new_n633_), .A3(new_n667_), .A4(new_n239_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT111), .Z(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(G57gat), .A3(new_n535_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n739_), .A2(KEYINPUT112), .A3(G57gat), .A4(new_n535_), .ZN(new_n743_));
  INV_X1    g542(.A(G57gat), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n593_), .A2(new_n321_), .A3(new_n365_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n631_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n746_), .A2(new_n238_), .A3(new_n237_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n748_), .B2(new_n536_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n742_), .A2(new_n743_), .A3(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n742_), .A2(KEYINPUT113), .A3(new_n743_), .A4(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1332gat));
  INV_X1    g553(.A(G64gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n739_), .B2(new_n641_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT48), .Z(new_n757_));
  INV_X1    g556(.A(new_n748_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n755_), .A3(new_n641_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1333gat));
  AOI21_X1  g559(.A(new_n369_), .B1(new_n739_), .B2(new_n417_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT49), .Z(new_n762_));
  NAND3_X1  g561(.A1(new_n758_), .A2(new_n369_), .A3(new_n417_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1334gat));
  INV_X1    g563(.A(G78gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n739_), .B2(new_n576_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT50), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n758_), .A2(new_n765_), .A3(new_n576_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1335gat));
  NAND2_X1  g568(.A1(new_n704_), .A2(new_n705_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n239_), .A2(new_n321_), .A3(new_n365_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n772_), .A2(new_n536_), .A3(new_n281_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n745_), .A2(new_n693_), .A3(new_n620_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT114), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n535_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n773_), .B1(new_n776_), .B2(new_n257_), .ZN(G1336gat));
  NOR3_X1   g576(.A1(new_n772_), .A2(new_n258_), .A3(new_n477_), .ZN(new_n778_));
  AOI21_X1  g577(.A(G92gat), .B1(new_n775_), .B2(new_n641_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n779_), .A2(KEYINPUT115), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(KEYINPUT115), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n778_), .B1(new_n780_), .B2(new_n781_), .ZN(G1337gat));
  AND2_X1   g581(.A1(new_n417_), .A2(new_n292_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n770_), .A2(new_n417_), .A3(new_n771_), .ZN(new_n784_));
  AOI22_X1  g583(.A1(new_n775_), .A2(new_n783_), .B1(G99gat), .B2(new_n784_), .ZN(new_n785_));
  XOR2_X1   g584(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n786_));
  XNOR2_X1  g585(.A(new_n785_), .B(new_n786_), .ZN(G1338gat));
  XNOR2_X1  g586(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n770_), .A2(new_n576_), .A3(new_n771_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(G106gat), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n790_), .A2(KEYINPUT52), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(KEYINPUT52), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n775_), .A2(new_n250_), .A3(new_n576_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n788_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n794_), .B(new_n788_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1339gat));
  XNOR2_X1  g597(.A(new_n361_), .B(new_n362_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n355_), .A2(new_n358_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(new_n347_), .A3(new_n341_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n325_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n799_), .A2(new_n317_), .A3(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n308_), .A2(new_n241_), .A3(new_n309_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n308_), .A2(KEYINPUT118), .A3(new_n241_), .A4(new_n309_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n310_), .A2(new_n811_), .ZN(new_n812_));
  AOI211_X1 g611(.A(KEYINPUT55), .B(new_n241_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n809_), .B(new_n810_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n316_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  INV_X1    g615(.A(new_n241_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n300_), .A2(KEYINPUT12), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n306_), .A2(new_n215_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n309_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n817_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT55), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n310_), .A2(new_n811_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n810_), .B1(new_n825_), .B2(new_n809_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n815_), .A2(new_n816_), .A3(new_n826_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n823_), .A2(new_n824_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n315_), .B1(new_n828_), .B2(new_n810_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n825_), .A2(new_n809_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT119), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT56), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT58), .B(new_n804_), .C1(new_n827_), .C2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n804_), .B1(new_n827_), .B2(new_n832_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n631_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n365_), .A2(new_n317_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n816_), .B1(new_n815_), .B2(new_n826_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n829_), .A2(new_n831_), .A3(KEYINPUT56), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n799_), .A2(new_n803_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n318_), .B2(new_n317_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n619_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n833_), .A2(new_n836_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT57), .B(new_n619_), .C1(new_n840_), .C2(new_n842_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n239_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n747_), .A2(new_n848_), .A3(new_n633_), .A4(new_n321_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT54), .B1(new_n632_), .B2(new_n365_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n847_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n576_), .A2(new_n641_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n417_), .A3(new_n535_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(G113gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n365_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n855_), .A2(new_n858_), .A3(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n859_), .B(new_n860_), .C1(new_n852_), .C2(new_n854_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n633_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n857_), .B1(new_n864_), .B2(new_n856_), .ZN(G1340gat));
  INV_X1    g664(.A(G120gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n321_), .B2(KEYINPUT60), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n855_), .B(new_n867_), .C1(KEYINPUT60), .C2(new_n866_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n321_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n866_), .ZN(G1341gat));
  INV_X1    g669(.A(G127gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n855_), .A2(new_n871_), .A3(new_n239_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n693_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n871_), .ZN(G1342gat));
  INV_X1    g673(.A(G134gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n855_), .A2(new_n875_), .A3(new_n620_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n631_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n875_), .ZN(G1343gat));
  NAND4_X1  g677(.A1(new_n592_), .A2(new_n576_), .A3(new_n535_), .A4(new_n477_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n852_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n365_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT121), .B(G141gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1344gat));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n667_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g684(.A1(new_n880_), .A2(new_n239_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT61), .B(G155gat), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1346gat));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n852_), .A2(new_n619_), .A3(new_n879_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(G162gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n700_), .A2(G162gat), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n852_), .A2(new_n879_), .A3(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n889_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n893_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n895_), .B(KEYINPUT122), .C1(G162gat), .C2(new_n890_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1347gat));
  NOR4_X1   g696(.A1(new_n592_), .A2(new_n576_), .A3(new_n477_), .A4(new_n535_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n852_), .A2(new_n899_), .ZN(new_n900_));
  AOI211_X1 g699(.A(KEYINPUT62), .B(new_n438_), .C1(new_n900_), .C2(new_n365_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n365_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(G169gat), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n900_), .B(new_n365_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n901_), .B1(new_n904_), .B2(new_n905_), .ZN(G1348gat));
  NAND2_X1  g705(.A1(new_n900_), .A2(new_n667_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g707(.A1(new_n900_), .A2(new_n239_), .ZN(new_n909_));
  MUX2_X1   g708(.A(new_n393_), .B(G183gat), .S(new_n909_), .Z(G1350gat));
  NOR3_X1   g709(.A1(new_n852_), .A2(new_n631_), .A3(new_n899_), .ZN(new_n911_));
  INV_X1    g710(.A(G190gat), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n620_), .A2(new_n394_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n852_), .A2(new_n899_), .A3(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(KEYINPUT123), .B1(new_n913_), .B2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n915_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n917_), .B(new_n918_), .C1(new_n912_), .C2(new_n911_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n916_), .A2(new_n919_), .ZN(G1351gat));
  NOR4_X1   g719(.A1(new_n417_), .A2(new_n477_), .A3(new_n572_), .A4(new_n535_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n843_), .A2(new_n844_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n834_), .A2(new_n835_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n924_), .A2(new_n746_), .A3(new_n833_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n925_), .A3(new_n846_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n693_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n849_), .A2(new_n850_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n922_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n365_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT124), .B(G197gat), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n930_), .B(new_n931_), .ZN(G1352gat));
  NAND2_X1  g731(.A1(new_n929_), .A2(new_n667_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g733(.A1(new_n929_), .A2(new_n239_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AND2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n935_), .B2(new_n936_), .ZN(G1354gat));
  NAND2_X1  g738(.A1(new_n746_), .A2(G218gat), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(KEYINPUT126), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n929_), .A2(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(G218gat), .ZN(new_n943_));
  OAI211_X1 g742(.A(new_n620_), .B(new_n921_), .C1(new_n847_), .C2(new_n851_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n944_), .B2(KEYINPUT125), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n946_), .B1(new_n929_), .B2(new_n620_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n942_), .B1(new_n945_), .B2(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(KEYINPUT127), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n950_));
  OAI211_X1 g749(.A(new_n950_), .B(new_n942_), .C1(new_n945_), .C2(new_n947_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n949_), .A2(new_n951_), .ZN(G1355gat));
endmodule


