//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT84), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G113gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G120gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT4), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT85), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT1), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n208_), .B(new_n209_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n207_), .B(KEYINPUT3), .Z(new_n216_));
  XOR2_X1   g015(.A(new_n209_), .B(KEYINPUT2), .Z(new_n217_));
  OAI221_X1 g016(.A(new_n212_), .B1(G155gat), .B2(G162gat), .C1(new_n216_), .C2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n205_), .A2(new_n206_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT94), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G225gat), .A2(G233gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G120gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n204_), .B(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n219_), .A2(KEYINPUT93), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n219_), .A2(KEYINPUT93), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n205_), .B1(KEYINPUT93), .B2(new_n219_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(KEYINPUT4), .A3(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n222_), .A2(new_n224_), .A3(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT95), .B(G85gat), .Z(new_n233_));
  XNOR2_X1  g032(.A(G1gat), .B(G29gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT0), .B(G57gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n235_), .B(new_n236_), .Z(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n229_), .A2(new_n230_), .ZN(new_n239_));
  OR3_X1    g038(.A1(new_n239_), .A2(KEYINPUT96), .A3(new_n224_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT96), .B1(new_n239_), .B2(new_n224_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n232_), .A2(new_n238_), .A3(new_n240_), .A4(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT97), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(KEYINPUT33), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n222_), .A2(new_n223_), .A3(new_n231_), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n239_), .B(KEYINPUT98), .Z(new_n247_));
  OAI211_X1 g046(.A(new_n237_), .B(new_n246_), .C1(new_n247_), .C2(new_n223_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n242_), .A2(new_n244_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT25), .B(G183gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT26), .B(G190gat), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n253_), .B1(G169gat), .B2(G176gat), .ZN(new_n254_));
  NOR3_X1   g053(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n252_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G183gat), .ZN(new_n257_));
  INV_X1    g056(.A(G190gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT23), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT80), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT23), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(G183gat), .A3(G190gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n260_), .B1(new_n264_), .B2(KEYINPUT80), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n256_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT91), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(G169gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(G183gat), .A2(G190gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n270_), .B1(new_n264_), .B2(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(G197gat), .B(G204gat), .Z(new_n275_));
  OAI21_X1  g074(.A(new_n274_), .B1(new_n275_), .B2(KEYINPUT21), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(KEYINPUT21), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G226gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT19), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT20), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n265_), .B1(G183gat), .B2(G190gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n270_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n256_), .A2(new_n263_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n278_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n283_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n279_), .A2(new_n282_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT92), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n285_), .A2(new_n286_), .A3(new_n278_), .ZN(new_n293_));
  OAI211_X1 g092(.A(KEYINPUT20), .B(new_n293_), .C1(new_n273_), .C2(new_n278_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n281_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n279_), .A2(KEYINPUT92), .A3(new_n282_), .A4(new_n289_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G8gat), .B(G36gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT18), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(G64gat), .ZN(new_n300_));
  INV_X1    g099(.A(G92gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n297_), .B(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n245_), .A2(new_n248_), .A3(new_n249_), .A4(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n232_), .A2(new_n241_), .A3(new_n240_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n237_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n242_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n278_), .A2(new_n272_), .A3(new_n266_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n289_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n281_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(new_n294_), .B2(new_n281_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n302_), .A2(KEYINPUT32), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n297_), .A2(new_n312_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n307_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n304_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G50gat), .ZN(new_n317_));
  OR3_X1    g116(.A1(new_n219_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n318_));
  INV_X1    g117(.A(G22gat), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT28), .B1(new_n219_), .B2(KEYINPUT29), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n319_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n317_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n323_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(G50gat), .A3(new_n321_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n328_), .B1(new_n327_), .B2(KEYINPUT90), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n332_));
  NAND2_X1  g131(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(G228gat), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n332_), .A2(new_n288_), .A3(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n337_), .B(KEYINPUT87), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT88), .B(KEYINPUT29), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n219_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT89), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n278_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n336_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n339_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n331_), .A2(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n330_), .B(new_n329_), .C1(new_n347_), .C2(new_n339_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n316_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT99), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n287_), .B(KEYINPUT30), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G15gat), .B(G43gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n354_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(KEYINPUT82), .Z(new_n362_));
  NOR2_X1   g161(.A1(new_n354_), .A2(new_n360_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT81), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n226_), .B(KEYINPUT31), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT83), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n365_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT99), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n316_), .A2(new_n369_), .A3(new_n351_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n353_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n368_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n351_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n349_), .A2(new_n368_), .A3(new_n350_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n307_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n303_), .A2(KEYINPUT27), .ZN(new_n377_));
  INV_X1    g176(.A(new_n302_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n311_), .A2(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(KEYINPUT27), .B(new_n379_), .C1(new_n297_), .C2(new_n378_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n375_), .A2(new_n376_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n371_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G230gat), .A2(G233gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(G71gat), .B(G78gat), .Z(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G57gat), .B(G64gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT11), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n388_), .A2(KEYINPUT11), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n386_), .A2(KEYINPUT11), .A3(new_n388_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(G99gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT10), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(G99gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G106gat), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n398_), .A2(KEYINPUT64), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT64), .B1(new_n398_), .B2(new_n399_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT9), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n301_), .A2(G85gat), .ZN(new_n404_));
  INV_X1    g203(.A(G85gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G92gat), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n403_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n403_), .A2(G85gat), .A3(G92gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT65), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT65), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G85gat), .B(G92gat), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n411_), .B(new_n408_), .C1(new_n412_), .C2(new_n403_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G99gat), .A2(G106gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT6), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(G99gat), .A3(G106gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n402_), .A2(new_n414_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT66), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT7), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n421_), .B(new_n422_), .C1(G99gat), .C2(G106gat), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n394_), .B(new_n399_), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI211_X1 g224(.A(KEYINPUT8), .B(new_n412_), .C1(new_n425_), .C2(new_n419_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n412_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT68), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT67), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT67), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT68), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n416_), .A2(new_n418_), .A3(new_n429_), .A4(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n425_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n416_), .A2(new_n418_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n427_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n426_), .B1(new_n435_), .B2(KEYINPUT8), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n393_), .B1(new_n420_), .B2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n402_), .A2(new_n414_), .A3(new_n419_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n393_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT8), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n429_), .A2(new_n431_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n419_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(new_n432_), .A3(new_n425_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n440_), .B1(new_n443_), .B2(new_n427_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n438_), .B(new_n439_), .C1(new_n444_), .C2(new_n426_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n385_), .B1(new_n437_), .B2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n437_), .A2(KEYINPUT12), .A3(new_n445_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n438_), .B1(new_n444_), .B2(new_n426_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT12), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n393_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n446_), .B1(new_n451_), .B2(new_n385_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G120gat), .B(G148gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT5), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(G176gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n455_), .B(G204gat), .Z(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n452_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(KEYINPUT69), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n452_), .A2(new_n457_), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n460_), .B(new_n461_), .Z(new_n462_));
  XOR2_X1   g261(.A(new_n462_), .B(KEYINPUT13), .Z(new_n463_));
  XNOR2_X1  g262(.A(G29gat), .B(G36gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT70), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(G43gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(G50gat), .ZN(new_n467_));
  INV_X1    g266(.A(G43gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n465_), .B(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n317_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT15), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT73), .B(G15gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(new_n319_), .ZN(new_n475_));
  INV_X1    g274(.A(G1gat), .ZN(new_n476_));
  INV_X1    g275(.A(G8gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT14), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G1gat), .B(G8gat), .Z(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n479_), .B(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n473_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n471_), .A2(new_n482_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT78), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n471_), .A2(new_n482_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n485_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n484_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n471_), .A2(KEYINPUT78), .A3(new_n482_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n486_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G113gat), .B(G141gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT79), .ZN(new_n495_));
  INV_X1    g294(.A(G169gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(G197gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n493_), .A2(new_n498_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n463_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n384_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n473_), .A2(new_n448_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G232gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT34), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT35), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n471_), .A2(new_n448_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n506_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n509_), .A2(new_n510_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n514_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n506_), .A2(new_n516_), .A3(new_n511_), .A4(new_n512_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(KEYINPUT72), .A3(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G190gat), .B(G218gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT71), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(G134gat), .ZN(new_n521_));
  INV_X1    g320(.A(G162gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n523_), .A2(KEYINPUT36), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n518_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n515_), .A2(new_n517_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(KEYINPUT36), .A3(new_n523_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT37), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n526_), .A2(KEYINPUT37), .A3(new_n528_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n482_), .B(new_n393_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT74), .B(KEYINPUT75), .Z(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G127gat), .B(G155gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G183gat), .B(G211gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n539_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n544_), .A2(new_n545_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n539_), .A2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT77), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(KEYINPUT77), .A3(new_n549_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n505_), .A2(new_n534_), .A3(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n307_), .B(KEYINPUT100), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n476_), .A3(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT38), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n526_), .A2(KEYINPUT101), .A3(new_n528_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT101), .B1(new_n526_), .B2(new_n528_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT102), .ZN(new_n563_));
  INV_X1    g362(.A(new_n561_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n559_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT102), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n547_), .A2(new_n549_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n384_), .A2(new_n568_), .A3(new_n570_), .A4(new_n504_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT103), .Z(new_n572_));
  AND2_X1   g371(.A1(new_n572_), .A2(new_n307_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n558_), .B1(new_n573_), .B2(new_n476_), .ZN(G1324gat));
  AND3_X1   g373(.A1(new_n384_), .A2(new_n504_), .A3(new_n568_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT104), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n575_), .A2(new_n576_), .A3(new_n570_), .A4(new_n381_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT104), .B1(new_n571_), .B2(new_n382_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(G8gat), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT39), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT39), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n577_), .A2(new_n581_), .A3(new_n578_), .A4(G8gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n554_), .A2(new_n477_), .A3(new_n381_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT40), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(KEYINPUT40), .A3(new_n584_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(G1325gat));
  INV_X1    g388(.A(G15gat), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n554_), .A2(new_n590_), .A3(new_n372_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n572_), .A2(new_n372_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n592_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT41), .B1(new_n592_), .B2(G15gat), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n591_), .B1(new_n593_), .B2(new_n594_), .ZN(G1326gat));
  XNOR2_X1  g394(.A(new_n351_), .B(KEYINPUT105), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n554_), .A2(new_n319_), .A3(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n572_), .A2(new_n596_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n599_), .B1(new_n600_), .B2(G22gat), .ZN(new_n601_));
  AOI211_X1 g400(.A(new_n319_), .B(new_n598_), .C1(new_n572_), .C2(new_n596_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n597_), .B1(new_n601_), .B2(new_n602_), .ZN(G1327gat));
  INV_X1    g402(.A(new_n552_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(new_n550_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n565_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT107), .B1(new_n505_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT107), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n384_), .A2(new_n609_), .A3(new_n504_), .A4(new_n606_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(G29gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n307_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT43), .B1(new_n384_), .B2(new_n534_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT43), .ZN(new_n615_));
  AOI211_X1 g414(.A(new_n615_), .B(new_n533_), .C1(new_n371_), .C2(new_n383_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n617_), .A2(KEYINPUT44), .A3(new_n504_), .A4(new_n553_), .ZN(new_n618_));
  AOI211_X1 g417(.A(new_n307_), .B(new_n381_), .C1(new_n373_), .C2(new_n374_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n316_), .A2(new_n369_), .A3(new_n351_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n369_), .B1(new_n316_), .B2(new_n351_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n619_), .B1(new_n622_), .B2(new_n368_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n615_), .B1(new_n623_), .B2(new_n533_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n384_), .A2(KEYINPUT43), .A3(new_n534_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n624_), .A2(new_n504_), .A3(new_n553_), .A4(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT44), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n618_), .A2(new_n628_), .A3(new_n556_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n613_), .B1(new_n629_), .B2(new_n612_), .ZN(G1328gat));
  NAND3_X1  g429(.A1(new_n618_), .A2(new_n628_), .A3(new_n381_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(G36gat), .ZN(new_n632_));
  INV_X1    g431(.A(G36gat), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n608_), .A2(new_n633_), .A3(new_n381_), .A4(new_n610_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT45), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT46), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n632_), .A2(new_n635_), .A3(KEYINPUT46), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1329gat));
  NAND3_X1  g439(.A1(new_n618_), .A2(new_n628_), .A3(new_n372_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G43gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n611_), .A2(new_n468_), .A3(new_n372_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT47), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n642_), .A2(KEYINPUT47), .A3(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1330gat));
  NAND3_X1  g447(.A1(new_n611_), .A2(new_n317_), .A3(new_n596_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n351_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n618_), .A2(new_n628_), .A3(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n651_), .B2(new_n317_), .ZN(G1331gat));
  INV_X1    g451(.A(G57gat), .ZN(new_n653_));
  INV_X1    g452(.A(new_n463_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n623_), .A2(new_n502_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT108), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT108), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n657_), .B1(new_n623_), .B2(new_n502_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n654_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n553_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n653_), .B1(new_n661_), .B2(new_n555_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n568_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(new_n654_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n655_), .A2(new_n664_), .A3(new_n605_), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT109), .B(G57gat), .Z(new_n666_));
  OR3_X1    g465(.A1(new_n665_), .A2(new_n376_), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n662_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT110), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT110), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n662_), .A2(new_n670_), .A3(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1332gat));
  OAI21_X1  g471(.A(G64gat), .B1(new_n665_), .B2(new_n382_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT48), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n382_), .A2(G64gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n661_), .B2(new_n675_), .ZN(G1333gat));
  OAI21_X1  g475(.A(G71gat), .B1(new_n665_), .B2(new_n368_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT49), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n368_), .A2(G71gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n661_), .B2(new_n679_), .ZN(G1334gat));
  INV_X1    g479(.A(new_n596_), .ZN(new_n681_));
  OR3_X1    g480(.A1(new_n661_), .A2(G78gat), .A3(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G78gat), .B1(new_n665_), .B2(new_n681_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(KEYINPUT111), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(KEYINPUT111), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n684_), .A2(KEYINPUT50), .A3(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT50), .B1(new_n684_), .B2(new_n685_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n682_), .B1(new_n686_), .B2(new_n687_), .ZN(G1335gat));
  NOR2_X1   g487(.A1(new_n654_), .A2(new_n502_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n624_), .A2(new_n553_), .A3(new_n625_), .A4(new_n689_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n690_), .A2(new_n405_), .A3(new_n376_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n659_), .A2(new_n606_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(new_n556_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n691_), .B1(new_n694_), .B2(new_n405_), .ZN(G1336gat));
  NOR3_X1   g494(.A1(new_n690_), .A2(new_n301_), .A3(new_n382_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n381_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(new_n301_), .ZN(G1337gat));
  OAI21_X1  g497(.A(G99gat), .B1(new_n690_), .B2(new_n368_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n372_), .A2(new_n398_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n692_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g501(.A(KEYINPUT52), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n690_), .A2(new_n351_), .ZN(new_n704_));
  OAI211_X1 g503(.A(KEYINPUT112), .B(new_n703_), .C1(new_n704_), .C2(new_n399_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n659_), .A2(new_n399_), .A3(new_n650_), .A4(new_n606_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n617_), .A2(new_n650_), .A3(new_n553_), .A4(new_n689_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n703_), .A2(KEYINPUT112), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n703_), .A2(KEYINPUT112), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n707_), .A2(G106gat), .A3(new_n708_), .A4(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n705_), .A2(new_n706_), .A3(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n705_), .A2(new_n712_), .A3(new_n706_), .A4(new_n710_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1339gat));
  INV_X1    g515(.A(KEYINPUT54), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n660_), .A2(new_n654_), .A3(new_n717_), .A4(new_n503_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n526_), .A2(KEYINPUT37), .A3(new_n528_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT37), .B1(new_n526_), .B2(new_n528_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n605_), .B(new_n503_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(KEYINPUT54), .B1(new_n721_), .B2(new_n463_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n718_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n489_), .A2(new_n484_), .A3(new_n491_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n498_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT117), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n483_), .A2(new_n490_), .A3(new_n485_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n499_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT56), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n451_), .A2(new_n385_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n451_), .A2(new_n385_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT55), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n451_), .A2(new_n733_), .A3(new_n385_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n730_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n729_), .B1(new_n735_), .B2(new_n457_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n733_), .B1(new_n451_), .B2(new_n385_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n385_), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT55), .B(new_n738_), .C1(new_n447_), .C2(new_n450_), .ZN(new_n739_));
  OAI22_X1  g538(.A1(new_n737_), .A2(new_n739_), .B1(new_n385_), .B2(new_n451_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(KEYINPUT56), .A3(new_n456_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n459_), .B1(new_n736_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n728_), .A2(new_n742_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT58), .Z(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(new_n533_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n735_), .B2(new_n457_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n740_), .A2(KEYINPUT114), .A3(new_n456_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n729_), .A3(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT115), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n747_), .A2(new_n751_), .A3(new_n729_), .A4(new_n748_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n750_), .A2(new_n741_), .A3(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n459_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(KEYINPUT116), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT116), .B1(new_n753_), .B2(new_n754_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n728_), .A2(new_n462_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n755_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT57), .B1(new_n759_), .B2(new_n562_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n753_), .A2(new_n754_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n753_), .A2(KEYINPUT116), .A3(new_n754_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n757_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n565_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n745_), .B1(new_n760_), .B2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n723_), .B1(new_n768_), .B2(new_n570_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n373_), .A2(new_n555_), .A3(new_n381_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(G113gat), .B1(new_n771_), .B2(new_n502_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n718_), .A2(new_n722_), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n744_), .A2(new_n533_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n765_), .A2(new_n766_), .A3(new_n565_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n766_), .B1(new_n765_), .B2(new_n565_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n774_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n773_), .B1(new_n777_), .B2(new_n553_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT59), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n770_), .A2(new_n779_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n771_), .B2(new_n779_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT118), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n781_), .B(new_n784_), .C1(new_n771_), .C2(new_n779_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n503_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n772_), .B1(new_n786_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g586(.A(G120gat), .B1(new_n782_), .B2(new_n654_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n225_), .B1(new_n654_), .B2(KEYINPUT60), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n771_), .B(new_n789_), .C1(KEYINPUT60), .C2(new_n225_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1341gat));
  AOI21_X1  g590(.A(G127gat), .B1(new_n771_), .B2(new_n605_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n569_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g593(.A(G134gat), .B1(new_n771_), .B2(new_n663_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n533_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(G134gat), .ZN(G1343gat));
  AOI21_X1  g596(.A(new_n773_), .B1(new_n777_), .B2(new_n569_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n555_), .A2(new_n381_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n374_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT119), .B1(new_n798_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803_));
  INV_X1    g602(.A(new_n801_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n769_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n802_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n502_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT120), .B(G141gat), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT121), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n807_), .B(new_n809_), .ZN(G1344gat));
  NAND2_X1  g609(.A1(new_n806_), .A2(new_n463_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g611(.A(KEYINPUT61), .B(G155gat), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n806_), .B2(new_n605_), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n553_), .B(new_n813_), .C1(new_n802_), .C2(new_n805_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n815_), .A2(new_n816_), .A3(new_n818_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n798_), .A2(KEYINPUT119), .A3(new_n801_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n803_), .B1(new_n769_), .B2(new_n804_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n605_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n813_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n806_), .A2(new_n605_), .A3(new_n814_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n817_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n819_), .A2(new_n825_), .ZN(G1346gat));
  AOI21_X1  g625(.A(G162gat), .B1(new_n806_), .B2(new_n663_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n533_), .B1(new_n802_), .B2(new_n805_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(G162gat), .B2(new_n828_), .ZN(G1347gat));
  NOR3_X1   g628(.A1(new_n556_), .A2(new_n382_), .A3(new_n368_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n778_), .A2(new_n596_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n502_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G169gat), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT124), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n496_), .A2(KEYINPUT22), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n496_), .A2(KEYINPUT22), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n832_), .A2(new_n502_), .A3(new_n838_), .A4(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n835_), .A2(new_n836_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n833_), .A2(G169gat), .A3(new_n841_), .A4(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n837_), .A2(new_n840_), .A3(new_n843_), .ZN(G1348gat));
  AOI21_X1  g643(.A(G176gat), .B1(new_n832_), .B2(new_n463_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n798_), .A2(new_n650_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n830_), .A2(G176gat), .A3(new_n463_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n845_), .B1(new_n846_), .B2(new_n847_), .ZN(G1349gat));
  INV_X1    g647(.A(new_n778_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(new_n681_), .A3(new_n830_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n850_), .A2(new_n569_), .A3(new_n250_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n851_), .A2(KEYINPUT125), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(KEYINPUT125), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n831_), .A2(new_n553_), .ZN(new_n854_));
  AOI21_X1  g653(.A(G183gat), .B1(new_n846_), .B2(new_n854_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n852_), .A2(new_n853_), .A3(new_n855_), .ZN(G1350gat));
  OAI21_X1  g655(.A(G190gat), .B1(new_n850_), .B2(new_n533_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n832_), .A2(new_n251_), .A3(new_n663_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1351gat));
  NOR2_X1   g658(.A1(new_n798_), .A2(new_n374_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n382_), .A2(new_n307_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n502_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g664(.A1(new_n862_), .A2(new_n654_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT126), .B(G204gat), .Z(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1353gat));
  NOR2_X1   g667(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n869_));
  AND2_X1   g668(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n862_), .A2(new_n569_), .A3(new_n869_), .A4(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n863_), .A2(new_n570_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n869_), .ZN(G1354gat));
  INV_X1    g672(.A(KEYINPUT127), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n863_), .A2(new_n874_), .A3(new_n663_), .ZN(new_n875_));
  INV_X1    g674(.A(G218gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT127), .B1(new_n862_), .B2(new_n568_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n863_), .A2(G218gat), .A3(new_n534_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1355gat));
endmodule


