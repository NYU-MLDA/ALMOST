//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_;
  XOR2_X1   g000(.A(G43gat), .B(G50gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G29gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT15), .Z(new_n205_));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT72), .B(G1gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(G8gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(G15gat), .B(G22gat), .Z(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n210_), .B(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n205_), .A2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n213_), .A2(new_n204_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G229gat), .A2(G233gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT73), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n213_), .B(new_n204_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G229gat), .A3(G233gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G113gat), .B(G141gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G169gat), .B(G197gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n222_), .B(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT74), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G85gat), .B(G92gat), .Z(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  OR4_X1    g032(.A1(KEYINPUT66), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n235_));
  OAI22_X1  g034(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n230_), .B1(new_n233_), .B2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT8), .ZN(new_n239_));
  INV_X1    g038(.A(G85gat), .ZN(new_n240_));
  INV_X1    g039(.A(G92gat), .ZN(new_n241_));
  NOR3_X1   g040(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT9), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n242_), .B1(new_n230_), .B2(KEYINPUT9), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT10), .B(G99gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(KEYINPUT64), .B(G106gat), .Z(new_n245_));
  OAI21_X1  g044(.A(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n246_), .A2(new_n233_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n239_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT68), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT12), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G57gat), .B(G64gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT11), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT67), .Z(new_n253_));
  XOR2_X1   g052(.A(G71gat), .B(G78gat), .Z(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(KEYINPUT11), .B2(new_n251_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n253_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n248_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n250_), .A2(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n249_), .A2(KEYINPUT12), .A3(new_n248_), .A4(new_n256_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G230gat), .A2(G233gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n248_), .A2(new_n256_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .A4(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n261_), .B1(new_n250_), .B2(new_n257_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n266_), .A2(KEYINPUT69), .A3(new_n260_), .A4(new_n259_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n257_), .ZN(new_n269_));
  OAI211_X1 g068(.A(G230gat), .B(G233gat), .C1(new_n269_), .C2(new_n261_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G120gat), .B(G148gat), .ZN(new_n271_));
  INV_X1    g070(.A(G204gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT5), .B(G176gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  NAND3_X1  g074(.A1(new_n268_), .A2(new_n270_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n275_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n279_), .A2(KEYINPUT13), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(KEYINPUT13), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT26), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G190gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT76), .ZN(new_n285_));
  NAND2_X1  g084(.A1(KEYINPUT75), .A2(G183gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT25), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(KEYINPUT75), .A2(KEYINPUT25), .A3(G183gat), .ZN(new_n289_));
  INV_X1    g088(.A(G190gat), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n288_), .A2(new_n289_), .B1(KEYINPUT26), .B2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT77), .B1(new_n285_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n296_), .B(new_n297_), .C1(new_n299_), .C2(KEYINPUT24), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT78), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n299_), .A2(KEYINPUT24), .A3(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n300_), .A2(new_n301_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n285_), .A2(KEYINPUT77), .A3(new_n291_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n293_), .A2(new_n305_), .A3(new_n306_), .A4(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  AND2_X1   g108(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n303_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n296_), .B(new_n297_), .C1(G183gat), .C2(G190gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n308_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G71gat), .B(G99gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT30), .B(KEYINPUT31), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(G43gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G127gat), .B(G134gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(G113gat), .A2(G120gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G113gat), .A2(G120gat), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n326_), .A2(new_n327_), .A3(KEYINPUT81), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT81), .ZN(new_n329_));
  INV_X1    g128(.A(G113gat), .ZN(new_n330_));
  INV_X1    g129(.A(G120gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G113gat), .A2(G120gat), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n329_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n325_), .B1(new_n328_), .B2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT81), .B1(new_n326_), .B2(new_n327_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n332_), .A2(new_n329_), .A3(new_n333_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(new_n324_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT80), .B(G15gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G227gat), .A2(G233gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n342_), .B(KEYINPUT79), .Z(new_n343_));
  XNOR2_X1  g142(.A(new_n341_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n323_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n323_), .A2(new_n345_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n336_), .A2(new_n337_), .A3(new_n324_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n324_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT100), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT100), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n335_), .A2(new_n352_), .A3(new_n338_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(G141gat), .ZN(new_n355_));
  INV_X1    g154(.A(G148gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G141gat), .A2(G148gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(KEYINPUT1), .B2(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n361_), .A2(KEYINPUT1), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n359_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365_));
  AND2_X1   g164(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n366_));
  NOR2_X1   g165(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT83), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n370_), .B(new_n365_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(KEYINPUT84), .A2(KEYINPUT2), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(G141gat), .A3(G148gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n358_), .A2(KEYINPUT84), .A3(KEYINPUT2), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(KEYINPUT84), .A2(KEYINPUT2), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n376_), .B1(new_n357_), .B2(KEYINPUT3), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n369_), .A2(new_n371_), .A3(new_n375_), .A4(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G155gat), .B(G162gat), .Z(new_n379_));
  AOI21_X1  g178(.A(new_n364_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT101), .B1(new_n354_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n354_), .A2(KEYINPUT101), .A3(new_n380_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT102), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT99), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n380_), .B2(new_n339_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n375_), .A2(new_n371_), .A3(new_n377_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n370_), .B1(new_n390_), .B2(new_n365_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n379_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n364_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n339_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(KEYINPUT99), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n388_), .A2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .A4(new_n397_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n354_), .A2(KEYINPUT101), .A3(new_n380_), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT99), .B1(new_n394_), .B2(new_n395_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n380_), .A2(new_n387_), .A3(new_n339_), .ZN(new_n401_));
  OAI22_X1  g200(.A1(new_n399_), .A2(new_n381_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n386_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT102), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT4), .B1(new_n394_), .B2(new_n395_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(new_n402_), .B2(KEYINPUT4), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n398_), .B(new_n404_), .C1(new_n406_), .C2(new_n386_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(G85gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT0), .B(G57gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n407_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n411_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G8gat), .B(G36gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(new_n241_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT18), .B(G64gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n417_), .B(new_n418_), .Z(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G226gat), .A2(G233gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT19), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT26), .B(G190gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT25), .B(G183gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n304_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(KEYINPUT95), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n300_), .B1(new_n427_), .B2(KEYINPUT95), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT96), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n313_), .B1(new_n430_), .B2(new_n315_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n315_), .A2(new_n430_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n428_), .A2(new_n429_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(G197gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n434_), .A2(G204gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT87), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n434_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n435_), .B1(new_n439_), .B2(G204gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(G211gat), .B(G218gat), .Z(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT21), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n440_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n437_), .A2(KEYINPUT88), .A3(new_n272_), .A4(new_n438_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(G197gat), .B2(new_n272_), .ZN(new_n447_));
  AND2_X1   g246(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n448_));
  NOR2_X1   g247(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT88), .B1(new_n450_), .B2(new_n272_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT21), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(KEYINPUT89), .B(KEYINPUT21), .Z(new_n453_));
  AOI21_X1  g252(.A(new_n441_), .B1(new_n440_), .B2(new_n453_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n452_), .A2(KEYINPUT90), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT90), .B1(new_n452_), .B2(new_n454_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n433_), .B(new_n445_), .C1(new_n455_), .C2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT20), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n458_), .A2(KEYINPUT105), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n445_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n458_), .A2(KEYINPUT105), .B1(new_n317_), .B2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n423_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n452_), .A2(new_n454_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT90), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n452_), .A2(KEYINPUT90), .A3(new_n454_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n444_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT20), .B1(new_n467_), .B2(new_n433_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n460_), .A2(new_n317_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n468_), .A2(new_n469_), .A3(new_n422_), .ZN(new_n470_));
  OAI211_X1 g269(.A(KEYINPUT32), .B(new_n420_), .C1(new_n462_), .C2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT20), .ZN(new_n472_));
  INV_X1    g271(.A(new_n433_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n472_), .B1(new_n460_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n307_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n475_), .A2(new_n292_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n306_), .A2(new_n304_), .A3(new_n302_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n476_), .A2(new_n477_), .B1(new_n315_), .B2(new_n314_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n467_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n423_), .B1(new_n474_), .B2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n423_), .B1(new_n467_), .B2(new_n478_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(new_n458_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT32), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n483_), .B1(new_n484_), .B2(new_n419_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n415_), .A2(new_n471_), .A3(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n397_), .B(new_n403_), .C1(new_n381_), .C2(new_n399_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT104), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n411_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n489_), .B1(new_n406_), .B2(new_n403_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n488_), .B1(new_n487_), .B2(new_n411_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n492_), .B1(new_n412_), .B2(KEYINPUT33), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(new_n407_), .B2(new_n411_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT103), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n419_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n422_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n422_), .B1(new_n460_), .B2(new_n317_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(KEYINPUT20), .A3(new_n457_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n420_), .A3(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n502_), .A3(KEYINPUT97), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT98), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT97), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n483_), .A2(new_n505_), .A3(new_n420_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  OAI211_X1 g306(.A(KEYINPUT103), .B(new_n494_), .C1(new_n407_), .C2(new_n411_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n493_), .A2(new_n497_), .A3(new_n507_), .A4(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n504_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n486_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT106), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n394_), .A2(KEYINPUT29), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n460_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G228gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT86), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n516_), .A2(KEYINPUT91), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n460_), .A2(new_n513_), .B1(KEYINPUT91), .B2(new_n516_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(new_n517_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G78gat), .B(G106gat), .Z(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT92), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n524_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n394_), .A2(KEYINPUT29), .ZN(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G22gat), .B(G50gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n526_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n523_), .A2(new_n525_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n520_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT93), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n521_), .B1(new_n520_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT94), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n536_), .A2(KEYINPUT94), .A3(new_n538_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n531_), .B1(new_n535_), .B2(new_n521_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n534_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n511_), .A2(new_n512_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n541_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n547_), .B1(new_n533_), .B2(new_n532_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n419_), .B1(new_n462_), .B2(new_n470_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(KEYINPUT27), .A3(new_n502_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT27), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n503_), .A2(new_n551_), .A3(new_n506_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n415_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n548_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n546_), .A2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n512_), .B1(new_n511_), .B2(new_n545_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n348_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  OR3_X1    g358(.A1(new_n548_), .A2(KEYINPUT107), .A3(new_n553_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n348_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT107), .B1(new_n548_), .B2(new_n553_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n555_), .A4(new_n562_), .ZN(new_n563_));
  AOI211_X1 g362(.A(new_n229_), .B(new_n282_), .C1(new_n559_), .C2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n248_), .A2(new_n205_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT34), .ZN(new_n567_));
  OAI221_X1 g366(.A(new_n565_), .B1(KEYINPUT35), .B2(new_n567_), .C1(new_n204_), .C2(new_n248_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(KEYINPUT35), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT36), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n572_), .B(new_n573_), .Z(new_n574_));
  AND3_X1   g373(.A1(new_n570_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n571_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n570_), .A2(new_n576_), .ZN(new_n577_));
  OAI22_X1  g376(.A1(new_n575_), .A2(new_n577_), .B1(KEYINPUT70), .B2(KEYINPUT37), .ZN(new_n578_));
  NAND2_X1  g377(.A1(KEYINPUT70), .A2(KEYINPUT37), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT71), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n578_), .B(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n213_), .B(new_n583_), .Z(new_n584_));
  INV_X1    g383(.A(new_n256_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(G211gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT16), .B(G183gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT68), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n592_), .A3(KEYINPUT17), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(KEYINPUT17), .B2(new_n591_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n587_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n586_), .A2(new_n593_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n582_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n564_), .A2(new_n599_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n600_), .A2(new_n207_), .A3(new_n555_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n601_), .A2(KEYINPUT38), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(KEYINPUT38), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n575_), .A2(new_n577_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT108), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(new_n598_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n564_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G1gat), .B1(new_n607_), .B2(new_n555_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n602_), .A2(new_n603_), .A3(new_n608_), .ZN(G1324gat));
  OR3_X1    g408(.A1(new_n600_), .A2(G8gat), .A3(new_n554_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G8gat), .B1(new_n607_), .B2(new_n554_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n611_), .A2(KEYINPUT39), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(KEYINPUT39), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n610_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g414(.A(G15gat), .B1(new_n607_), .B2(new_n348_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n616_), .A2(KEYINPUT41), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(KEYINPUT41), .ZN(new_n618_));
  OR3_X1    g417(.A1(new_n600_), .A2(G15gat), .A3(new_n348_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .ZN(G1326gat));
  OAI21_X1  g419(.A(G22gat), .B1(new_n607_), .B2(new_n545_), .ZN(new_n621_));
  XOR2_X1   g420(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n545_), .A2(G22gat), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n623_), .B1(new_n600_), .B2(new_n624_), .ZN(G1327gat));
  INV_X1    g424(.A(new_n604_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n597_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n564_), .A2(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n628_), .A2(G29gat), .A3(new_n555_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n282_), .A2(new_n229_), .A3(new_n597_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n559_), .A2(new_n563_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n632_), .B2(new_n582_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n582_), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT43), .B(new_n634_), .C1(new_n559_), .C2(new_n563_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n630_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT44), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(KEYINPUT44), .B(new_n630_), .C1(new_n633_), .C2(new_n635_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n415_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n629_), .B1(new_n640_), .B2(G29gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT110), .ZN(G1328gat));
  NAND3_X1  g441(.A1(new_n638_), .A2(new_n553_), .A3(new_n639_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT111), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n638_), .A2(KEYINPUT111), .A3(new_n553_), .A4(new_n639_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(G36gat), .A3(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n628_), .A2(G36gat), .A3(new_n554_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT45), .Z(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT46), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n647_), .A2(new_n649_), .A3(KEYINPUT46), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1329gat));
  NAND2_X1  g453(.A1(new_n638_), .A2(new_n639_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G43gat), .B1(new_n655_), .B2(new_n348_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n561_), .A2(new_n322_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n628_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n658_), .B(new_n660_), .ZN(G1330gat));
  OAI21_X1  g460(.A(G50gat), .B1(new_n655_), .B2(new_n545_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n545_), .A2(G50gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n662_), .B1(new_n628_), .B2(new_n663_), .ZN(G1331gat));
  INV_X1    g463(.A(new_n282_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(new_n228_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n666_), .A2(new_n632_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(new_n599_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G57gat), .B1(new_n668_), .B2(new_n415_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n667_), .A2(new_n606_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n555_), .A2(KEYINPUT113), .ZN(new_n671_));
  MUX2_X1   g470(.A(KEYINPUT113), .B(new_n671_), .S(G57gat), .Z(new_n672_));
  AOI21_X1  g471(.A(new_n669_), .B1(new_n670_), .B2(new_n672_), .ZN(G1332gat));
  INV_X1    g472(.A(G64gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n670_), .B2(new_n553_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT48), .Z(new_n676_));
  NAND2_X1  g475(.A1(new_n553_), .A2(new_n674_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT114), .Z(new_n678_));
  NAND2_X1  g477(.A1(new_n668_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(G1333gat));
  INV_X1    g479(.A(G71gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n670_), .B2(new_n561_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT49), .Z(new_n683_));
  NAND3_X1  g482(.A1(new_n668_), .A2(new_n681_), .A3(new_n561_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1334gat));
  INV_X1    g484(.A(G78gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n670_), .B2(new_n548_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT50), .Z(new_n688_));
  NAND3_X1  g487(.A1(new_n668_), .A2(new_n686_), .A3(new_n548_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1335gat));
  AND2_X1   g489(.A1(new_n667_), .A2(new_n627_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G85gat), .B1(new_n691_), .B2(new_n415_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n632_), .A2(new_n582_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT43), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n632_), .A2(new_n631_), .A3(new_n582_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n696_), .A2(new_n598_), .A3(new_n666_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n555_), .A2(new_n240_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n692_), .B1(new_n697_), .B2(new_n698_), .ZN(G1336gat));
  AOI21_X1  g498(.A(G92gat), .B1(new_n691_), .B2(new_n553_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n554_), .A2(new_n241_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n697_), .B2(new_n701_), .ZN(G1337gat));
  INV_X1    g501(.A(G99gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n697_), .B2(new_n561_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n667_), .A2(new_n627_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n705_), .A2(new_n244_), .A3(new_n348_), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n704_), .A2(new_n706_), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n707_));
  NAND2_X1  g506(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(G1338gat));
  OR3_X1    g508(.A1(new_n705_), .A2(new_n245_), .A3(new_n545_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n696_), .A2(new_n548_), .A3(new_n598_), .A4(new_n666_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT52), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n711_), .A2(new_n712_), .A3(G106gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n711_), .B2(G106gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g515(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n717_), .A2(new_n555_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n718_), .A2(KEYINPUT59), .ZN(new_n719_));
  INV_X1    g518(.A(new_n275_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT55), .B1(new_n265_), .B2(new_n267_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n266_), .A2(KEYINPUT55), .A3(new_n260_), .A4(new_n259_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n266_), .A2(new_n259_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n260_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n721_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT56), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT56), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n727_), .B(new_n720_), .C1(new_n721_), .C2(new_n724_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n726_), .A2(new_n228_), .A3(new_n276_), .A4(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n222_), .A2(new_n225_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n216_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(new_n218_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n226_), .B1(new_n220_), .B2(new_n218_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n730_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n604_), .B1(new_n729_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT57), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n726_), .A2(new_n276_), .A3(new_n734_), .A4(new_n728_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT58), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n728_), .A2(new_n276_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n742_), .A2(KEYINPUT58), .A3(new_n734_), .A4(new_n726_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n741_), .A2(new_n582_), .A3(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(KEYINPUT57), .B2(new_n736_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT117), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n738_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n736_), .A2(KEYINPUT57), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(KEYINPUT117), .A3(new_n744_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n597_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n665_), .A2(new_n599_), .A3(new_n229_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT54), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n719_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n745_), .B2(new_n738_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n748_), .A2(KEYINPUT116), .A3(new_n737_), .A4(new_n744_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n598_), .A3(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n751_), .B(KEYINPUT54), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n718_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT59), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n754_), .B(new_n228_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G113gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(new_n330_), .A3(new_n228_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT118), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n763_), .A2(new_n764_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1340gat));
  OAI21_X1  g568(.A(new_n331_), .B1(new_n665_), .B2(KEYINPUT60), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n760_), .B(new_n770_), .C1(KEYINPUT60), .C2(new_n331_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n760_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n747_), .A2(new_n749_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n598_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n759_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n772_), .A2(KEYINPUT59), .B1(new_n775_), .B2(new_n719_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n282_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n771_), .B1(new_n778_), .B2(new_n331_), .ZN(G1341gat));
  NOR2_X1   g578(.A1(new_n759_), .A2(new_n598_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n718_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G127gat), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT119), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n597_), .A2(G127gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n776_), .B2(new_n784_), .ZN(G1342gat));
  AOI21_X1  g584(.A(G134gat), .B1(new_n760_), .B2(new_n605_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n582_), .A2(G134gat), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT120), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n786_), .B1(new_n776_), .B2(new_n788_), .ZN(G1343gat));
  NAND2_X1  g588(.A1(new_n758_), .A2(new_n759_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n548_), .A2(new_n348_), .A3(new_n415_), .A4(new_n554_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT121), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n228_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n282_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g596(.A1(new_n780_), .A2(new_n792_), .ZN(new_n798_));
  XOR2_X1   g597(.A(KEYINPUT61), .B(G155gat), .Z(new_n799_));
  XNOR2_X1  g598(.A(new_n798_), .B(new_n799_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(G1346gat));
  AOI21_X1  g601(.A(G162gat), .B1(new_n793_), .B2(new_n605_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n582_), .A2(G162gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n793_), .B2(new_n804_), .ZN(G1347gat));
  NOR3_X1   g604(.A1(new_n548_), .A2(new_n348_), .A3(new_n415_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n553_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n775_), .A2(new_n228_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT62), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(KEYINPUT124), .A3(new_n810_), .A4(G169gat), .ZN(new_n811_));
  INV_X1    g610(.A(G169gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n807_), .B1(new_n774_), .B2(new_n759_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n228_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n811_), .B1(new_n814_), .B2(new_n810_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT124), .B1(new_n814_), .B2(new_n810_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n310_), .A2(new_n311_), .ZN(new_n817_));
  OAI22_X1  g616(.A1(new_n815_), .A2(new_n816_), .B1(new_n817_), .B2(new_n809_), .ZN(G1348gat));
  AOI21_X1  g617(.A(G176gat), .B1(new_n813_), .B2(new_n282_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n665_), .A2(new_n309_), .A3(new_n807_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n790_), .B2(new_n820_), .ZN(G1349gat));
  AOI21_X1  g620(.A(G183gat), .B1(new_n780_), .B2(new_n808_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n598_), .A2(new_n425_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n813_), .B2(new_n823_), .ZN(G1350gat));
  NAND3_X1  g623(.A1(new_n813_), .A2(new_n424_), .A3(new_n605_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n813_), .A2(new_n582_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n290_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT125), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT125), .B(new_n825_), .C1(new_n826_), .C2(new_n290_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1351gat));
  NOR4_X1   g630(.A1(new_n561_), .A2(new_n545_), .A3(new_n554_), .A4(new_n415_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n790_), .A2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(new_n229_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(new_n434_), .ZN(G1352gat));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n665_), .ZN(new_n836_));
  XOR2_X1   g635(.A(KEYINPUT126), .B(G204gat), .Z(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1353gat));
  AND2_X1   g637(.A1(new_n790_), .A2(new_n832_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT127), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n598_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n841_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT127), .B1(new_n833_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1354gat));
  AND3_X1   g646(.A1(new_n839_), .A2(G218gat), .A3(new_n582_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G218gat), .B1(new_n839_), .B2(new_n605_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1355gat));
endmodule


