//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n205_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n204_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(new_n212_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G229gat), .A2(G233gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT69), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n214_), .B(new_n212_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n218_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n213_), .A2(new_n222_), .A3(new_n217_), .A4(new_n215_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n219_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G141gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G169gat), .B(G197gat), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n225_), .B(new_n226_), .Z(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n219_), .A2(new_n221_), .A3(new_n223_), .A4(new_n227_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G169gat), .ZN(new_n233_));
  INV_X1    g032(.A(G176gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT87), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT23), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n241_));
  INV_X1    g040(.A(G183gat), .ZN(new_n242_));
  INV_X1    g041(.A(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n235_), .A2(new_n237_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n238_), .B(KEYINPUT23), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT24), .ZN(new_n249_));
  INV_X1    g048(.A(G169gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(new_n234_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n242_), .A2(KEYINPUT25), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G183gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT84), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT85), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n243_), .A2(KEYINPUT26), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT26), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(G190gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n258_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT84), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n253_), .A2(new_n255_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(G190gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n243_), .A2(KEYINPUT26), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(KEYINPUT85), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n257_), .A2(new_n262_), .A3(new_n264_), .A4(new_n267_), .ZN(new_n268_));
  OR3_X1    g067(.A1(KEYINPUT71), .A2(G169gat), .A3(G176gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT71), .B1(G169gat), .B2(G176gat), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n269_), .A2(KEYINPUT24), .A3(new_n236_), .A4(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n252_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n271_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n264_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n263_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n265_), .A2(new_n266_), .A3(KEYINPUT85), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT85), .B1(new_n265_), .B2(new_n266_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n275_), .B1(new_n278_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT86), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n247_), .B1(new_n274_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G211gat), .B(G218gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G204gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G197gat), .ZN(new_n288_));
  INV_X1    g087(.A(G197gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G204gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n286_), .A2(KEYINPUT21), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT81), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(new_n287_), .A3(G197gat), .ZN(new_n294_));
  OAI211_X1 g093(.A(KEYINPUT21), .B(new_n294_), .C1(new_n291_), .C2(new_n293_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n285_), .B1(new_n291_), .B2(KEYINPUT21), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n292_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT88), .B1(new_n284_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT88), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n286_), .A2(KEYINPUT21), .A3(new_n291_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n294_), .A2(KEYINPUT21), .ZN(new_n302_));
  INV_X1    g101(.A(new_n291_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(KEYINPUT81), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n301_), .B1(new_n304_), .B2(new_n296_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n268_), .A2(KEYINPUT86), .A3(new_n271_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT86), .B1(new_n268_), .B2(new_n271_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n306_), .A2(new_n307_), .A3(new_n252_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n300_), .B(new_n305_), .C1(new_n308_), .C2(new_n247_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT19), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n245_), .A2(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n240_), .A2(new_n244_), .A3(KEYINPUT72), .A4(new_n241_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(G169gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n270_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(KEYINPUT71), .A2(G169gat), .A3(G176gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n249_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n253_), .B(new_n255_), .C1(new_n259_), .C2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT70), .B1(new_n265_), .B2(new_n266_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n321_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n271_), .A2(new_n248_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n318_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT20), .B1(new_n327_), .B2(new_n305_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT83), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI211_X1 g129(.A(KEYINPUT83), .B(KEYINPUT20), .C1(new_n327_), .C2(new_n305_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n299_), .A2(new_n309_), .A3(new_n312_), .A4(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n252_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(new_n282_), .B2(KEYINPUT86), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n298_), .B(new_n246_), .C1(new_n335_), .C2(new_n306_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT20), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n337_), .B1(new_n327_), .B2(new_n305_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(new_n311_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n333_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n341_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT92), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n341_), .A2(KEYINPUT92), .A3(new_n346_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT27), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n336_), .A2(new_n312_), .A3(new_n338_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n299_), .A2(new_n309_), .A3(new_n332_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n352_), .B1(new_n353_), .B2(new_n311_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n346_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n351_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n349_), .A2(new_n350_), .A3(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n354_), .A2(new_n355_), .ZN(new_n358_));
  AOI211_X1 g157(.A(new_n346_), .B(new_n352_), .C1(new_n353_), .C2(new_n311_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n351_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT93), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n364_));
  INV_X1    g163(.A(G155gat), .ZN(new_n365_));
  INV_X1    g164(.A(G162gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n367_), .A2(KEYINPUT79), .A3(new_n368_), .A4(new_n369_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n374_));
  INV_X1    g173(.A(G141gat), .ZN(new_n375_));
  INV_X1    g174(.A(G148gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT3), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n374_), .A2(new_n379_), .A3(new_n375_), .A4(new_n376_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n378_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT78), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n372_), .B(new_n373_), .C1(new_n382_), .C2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G141gat), .A2(G148gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n375_), .A2(new_n376_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n368_), .A2(KEYINPUT76), .A3(KEYINPUT1), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT76), .B1(new_n368_), .B2(KEYINPUT1), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n367_), .B(new_n369_), .C1(KEYINPUT1), .C2(new_n368_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n386_), .B(new_n387_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n385_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n298_), .B1(new_n393_), .B2(KEYINPUT29), .ZN(new_n394_));
  AND2_X1   g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n394_), .A2(new_n396_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n363_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n394_), .A2(new_n396_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n394_), .A2(new_n396_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n363_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT82), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n399_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(KEYINPUT82), .B(new_n363_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G22gat), .B(G50gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT28), .B1(new_n393_), .B2(KEYINPUT29), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT28), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n385_), .A2(new_n409_), .A3(new_n410_), .A4(new_n392_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n407_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n408_), .A2(new_n411_), .A3(new_n407_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n413_), .A2(KEYINPUT80), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT80), .B1(new_n413_), .B2(new_n414_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n405_), .B(new_n406_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n399_), .A2(new_n403_), .A3(new_n414_), .A4(new_n413_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G113gat), .B(G120gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G134gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(G127gat), .ZN(new_n423_));
  INV_X1    g222(.A(G127gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G134gat), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n423_), .A2(new_n425_), .A3(KEYINPUT73), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT73), .B1(new_n423_), .B2(new_n425_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n421_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n423_), .A2(new_n425_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT73), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n423_), .A2(new_n425_), .A3(KEYINPUT73), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n420_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G71gat), .B(G99gat), .ZN(new_n435_));
  INV_X1    g234(.A(G43gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n327_), .B(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G227gat), .A2(G233gat), .ZN(new_n440_));
  INV_X1    g239(.A(G15gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT30), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT31), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT74), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT31), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n443_), .B(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n327_), .A2(new_n437_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n327_), .A2(new_n437_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n445_), .A2(new_n446_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n446_), .B1(new_n445_), .B2(new_n451_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n434_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n445_), .A2(new_n451_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT74), .ZN(new_n457_));
  INV_X1    g256(.A(new_n434_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(new_n452_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G1gat), .B(G29gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(G85gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT0), .B(G57gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n462_), .B(new_n463_), .Z(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G225gat), .A2(G233gat), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n385_), .A2(new_n434_), .A3(new_n392_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n434_), .B1(new_n385_), .B2(new_n392_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT4), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n393_), .A2(new_n470_), .A3(new_n458_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n467_), .A2(new_n468_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n471_), .B1(new_n472_), .B2(KEYINPUT4), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n465_), .B(new_n469_), .C1(new_n473_), .C2(new_n466_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n393_), .A2(new_n458_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n385_), .A2(new_n434_), .A3(new_n392_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(KEYINPUT4), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n468_), .A2(new_n470_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n466_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n469_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n464_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n474_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n460_), .A2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n361_), .A2(new_n362_), .A3(new_n419_), .A4(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n357_), .A2(new_n419_), .A3(new_n360_), .A4(new_n483_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT93), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n482_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n357_), .A2(new_n488_), .A3(new_n360_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n417_), .A2(new_n418_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n355_), .A2(KEYINPUT32), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n341_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT91), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n354_), .A2(new_n491_), .B1(new_n481_), .B2(new_n474_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n341_), .A2(KEYINPUT91), .A3(new_n492_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT33), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT90), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n469_), .B1(new_n473_), .B2(new_n466_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n501_), .B2(new_n464_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n464_), .B(new_n500_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n477_), .A2(new_n466_), .A3(new_n478_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n475_), .A2(new_n476_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n504_), .B(new_n465_), .C1(new_n466_), .C2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n502_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n353_), .A2(new_n311_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n352_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n346_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n354_), .A2(new_n355_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n508_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n490_), .B1(new_n498_), .B2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n460_), .B1(new_n489_), .B2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n232_), .B1(new_n487_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G230gat), .A2(G233gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G85gat), .B(G92gat), .Z(new_n520_));
  NOR2_X1   g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT7), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT6), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n520_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT8), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT10), .B(G99gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT64), .ZN(new_n530_));
  INV_X1    g329(.A(G106gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n526_), .ZN(new_n533_));
  XOR2_X1   g332(.A(KEYINPUT65), .B(G85gat), .Z(new_n534_));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT66), .B(G92gat), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G85gat), .A2(G92gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT9), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n532_), .B(new_n533_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n528_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G57gat), .B(G64gat), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n544_), .A2(KEYINPUT11), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(KEYINPUT11), .ZN(new_n546_));
  XOR2_X1   g345(.A(G71gat), .B(G78gat), .Z(new_n547_));
  NAND3_X1  g346(.A1(new_n545_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n546_), .A2(new_n547_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n543_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n528_), .A2(new_n542_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(new_n549_), .A3(new_n548_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(KEYINPUT12), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT12), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n552_), .A2(new_n555_), .A3(new_n549_), .A4(new_n548_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n519_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n518_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n559_), .A2(new_n563_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT13), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n564_), .A2(KEYINPUT13), .A3(new_n565_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G134gat), .B(G162gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n573_), .A2(new_n574_), .ZN(new_n576_));
  XOR2_X1   g375(.A(KEYINPUT67), .B(KEYINPUT34), .Z(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT35), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n543_), .A2(new_n214_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n205_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n552_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n581_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT68), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n552_), .A2(new_n204_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n583_), .B2(new_n552_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n579_), .A2(new_n580_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n585_), .A2(new_n586_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n575_), .B(new_n576_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n586_), .A2(new_n585_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT68), .B1(new_n589_), .B2(new_n581_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n595_), .A2(new_n574_), .A3(new_n573_), .A4(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n594_), .A2(new_n597_), .A3(KEYINPUT37), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n550_), .B(new_n212_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n603_), .B(new_n604_), .Z(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT17), .ZN(new_n607_));
  XOR2_X1   g406(.A(G127gat), .B(G155gat), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT16), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  OR3_X1    g410(.A1(new_n606_), .A2(new_n607_), .A3(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(KEYINPUT17), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n606_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n570_), .A2(new_n602_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n517_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT94), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n517_), .A2(KEYINPUT94), .A3(new_n616_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n619_), .A2(new_n207_), .A3(new_n482_), .A4(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT95), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n623_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n598_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n487_), .B2(new_n516_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n570_), .A2(new_n232_), .A3(new_n615_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n482_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n624_), .A2(new_n625_), .A3(new_n631_), .ZN(G1324gat));
  INV_X1    g431(.A(new_n361_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n627_), .A2(new_n633_), .A3(new_n628_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(G8gat), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT96), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(new_n637_), .A3(G8gat), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n636_), .A2(KEYINPUT39), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n635_), .A2(KEYINPUT96), .A3(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n619_), .A2(new_n208_), .A3(new_n633_), .A4(new_n620_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT98), .B1(new_n639_), .B2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n636_), .A2(KEYINPUT39), .A3(new_n638_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n641_), .A4(new_n642_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n644_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1325gat));
  OAI21_X1  g452(.A(G15gat), .B1(new_n629_), .B2(new_n460_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT99), .Z(new_n655_));
  OR2_X1    g454(.A1(new_n655_), .A2(KEYINPUT41), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(KEYINPUT41), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n619_), .A2(new_n620_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n460_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n441_), .A3(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n656_), .A2(new_n657_), .A3(new_n660_), .ZN(G1326gat));
  XNOR2_X1  g460(.A(new_n490_), .B(KEYINPUT100), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n627_), .A2(new_n628_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G22gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT42), .ZN(new_n665_));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n662_), .A2(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT101), .Z(new_n668_));
  NAND2_X1  g467(.A1(new_n658_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n665_), .A2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT102), .Z(G1327gat));
  NAND2_X1  g470(.A1(new_n626_), .A2(new_n615_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n570_), .A2(new_n672_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n517_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n675_), .A2(G29gat), .A3(new_n630_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n568_), .A2(new_n231_), .A3(new_n569_), .A4(new_n615_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT103), .ZN(new_n678_));
  INV_X1    g477(.A(new_n602_), .ZN(new_n679_));
  AOI211_X1 g478(.A(KEYINPUT43), .B(new_n679_), .C1(new_n487_), .C2(new_n516_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n485_), .A2(KEYINPUT93), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n485_), .A2(KEYINPUT93), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n516_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n681_), .B1(new_n684_), .B2(new_n602_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n678_), .B1(new_n680_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n678_), .B(KEYINPUT44), .C1(new_n680_), .C2(new_n685_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n482_), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n676_), .B1(new_n690_), .B2(G29gat), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT104), .ZN(G1328gat));
  INV_X1    g491(.A(G36gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n674_), .A2(new_n693_), .A3(new_n633_), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n688_), .A2(new_n633_), .A3(new_n689_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(KEYINPUT105), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n688_), .A2(new_n699_), .A3(new_n633_), .A4(new_n689_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G36gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n696_), .B1(new_n698_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(KEYINPUT46), .B(new_n696_), .C1(new_n698_), .C2(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  AND2_X1   g505(.A1(new_n688_), .A2(new_n689_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(G43gat), .A3(new_n659_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n436_), .B1(new_n675_), .B2(new_n460_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(KEYINPUT47), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT47), .B1(new_n708_), .B2(new_n709_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1330gat));
  AOI21_X1  g511(.A(G50gat), .B1(new_n674_), .B2(new_n662_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n490_), .A2(G50gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n707_), .B2(new_n714_), .ZN(G1331gat));
  INV_X1    g514(.A(new_n615_), .ZN(new_n716_));
  AND4_X1   g515(.A1(new_n232_), .A2(new_n627_), .A3(new_n570_), .A4(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(G57gat), .A3(new_n482_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n718_), .A2(new_n719_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n231_), .B1(new_n487_), .B2(new_n516_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n722_), .A2(new_n570_), .A3(new_n716_), .A4(new_n679_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n482_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n720_), .A2(new_n721_), .A3(new_n725_), .ZN(G1332gat));
  NOR2_X1   g525(.A1(new_n361_), .A2(G64gat), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT109), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n724_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n717_), .A2(new_n633_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G64gat), .ZN(new_n731_));
  XOR2_X1   g530(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n731_), .A2(new_n732_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT110), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n737_), .B(new_n729_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1333gat));
  INV_X1    g538(.A(G71gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n717_), .B2(new_n659_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT49), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n724_), .A2(new_n740_), .A3(new_n659_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1334gat));
  INV_X1    g543(.A(G78gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n717_), .B2(new_n662_), .ZN(new_n746_));
  XOR2_X1   g545(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n724_), .A2(new_n745_), .A3(new_n662_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1335gat));
  INV_X1    g549(.A(new_n722_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n570_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n672_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G85gat), .B1(new_n753_), .B2(new_n482_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n680_), .A2(new_n685_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n570_), .A2(new_n232_), .A3(new_n615_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT112), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n482_), .A2(new_n534_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n754_), .B1(new_n759_), .B2(new_n760_), .ZN(G1336gat));
  AOI21_X1  g560(.A(G92gat), .B1(new_n753_), .B2(new_n633_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n633_), .A2(new_n536_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT113), .Z(new_n764_));
  AOI21_X1  g563(.A(new_n762_), .B1(new_n759_), .B2(new_n764_), .ZN(G1337gat));
  NAND3_X1  g564(.A1(new_n755_), .A2(new_n659_), .A3(new_n757_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n659_), .A2(new_n530_), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n766_), .A2(G99gat), .B1(new_n753_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n768_), .A2(KEYINPUT114), .A3(new_n769_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n768_), .A2(KEYINPUT115), .A3(new_n769_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT115), .B1(new_n768_), .B2(new_n769_), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n772_), .A2(new_n773_), .B1(new_n774_), .B2(new_n775_), .ZN(G1338gat));
  NAND3_X1  g575(.A1(new_n753_), .A2(new_n531_), .A3(new_n490_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n755_), .A2(new_n490_), .A3(new_n757_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(new_n779_), .A3(G106gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G106gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n784_), .B(new_n777_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1339gat));
  NOR2_X1   g585(.A1(new_n633_), .A2(new_n490_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n460_), .A2(new_n630_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n565_), .A2(new_n231_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n554_), .A2(new_n556_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n518_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n554_), .A2(new_n556_), .A3(new_n519_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(KEYINPUT55), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n563_), .B1(new_n557_), .B2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n796_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n790_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n227_), .B1(new_n220_), .B2(new_n217_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n230_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n626_), .B1(new_n800_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT116), .B1(new_n806_), .B2(KEYINPUT57), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  INV_X1    g608(.A(new_n799_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n797_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n804_), .B1(new_n811_), .B2(new_n790_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n808_), .B(new_n809_), .C1(new_n812_), .C2(new_n626_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n803_), .B1(new_n559_), .B2(new_n563_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n815_), .B(KEYINPUT58), .C1(new_n798_), .C2(new_n799_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n602_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT58), .B1(new_n811_), .B2(new_n815_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n814_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n807_), .A2(new_n813_), .A3(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n602_), .A2(new_n816_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n811_), .A2(new_n815_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(new_n824_), .A3(KEYINPUT117), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n806_), .A2(KEYINPUT57), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n615_), .B1(new_n820_), .B2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n752_), .A2(new_n232_), .A3(new_n716_), .A4(new_n679_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT54), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n789_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(G113gat), .B1(new_n831_), .B2(new_n231_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n831_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT59), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT59), .ZN(new_n835_));
  INV_X1    g634(.A(new_n789_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(KEYINPUT118), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(KEYINPUT118), .B2(new_n836_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n830_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n806_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n840_), .A2(new_n809_), .B1(new_n821_), .B2(new_n824_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n716_), .B1(new_n841_), .B2(new_n826_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n838_), .B1(new_n839_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n834_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n231_), .A2(G113gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT119), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n832_), .B1(new_n845_), .B2(new_n847_), .ZN(G1340gat));
  INV_X1    g647(.A(KEYINPUT60), .ZN(new_n849_));
  AOI21_X1  g648(.A(G120gat), .B1(new_n570_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT120), .B1(new_n849_), .B2(G120gat), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n831_), .B(new_n852_), .C1(new_n850_), .C2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n843_), .B(new_n570_), .C1(new_n831_), .C2(new_n835_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G120gat), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n855_), .A2(new_n856_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n854_), .B1(new_n858_), .B2(new_n859_), .ZN(G1341gat));
  OAI21_X1  g659(.A(new_n424_), .B1(new_n833_), .B2(new_n615_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n615_), .A2(KEYINPUT122), .ZN(new_n862_));
  MUX2_X1   g661(.A(KEYINPUT122), .B(new_n862_), .S(G127gat), .Z(new_n863_));
  OAI211_X1 g662(.A(new_n843_), .B(new_n863_), .C1(new_n831_), .C2(new_n835_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n861_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT123), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n861_), .A2(new_n864_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1342gat));
  OAI21_X1  g668(.A(G134gat), .B1(new_n844_), .B2(new_n679_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n831_), .A2(new_n422_), .A3(new_n626_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1343gat));
  NAND2_X1  g671(.A1(new_n828_), .A2(new_n830_), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n633_), .A2(new_n419_), .A3(new_n630_), .A4(new_n659_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n232_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n375_), .ZN(G1344gat));
  NOR2_X1   g676(.A1(new_n875_), .A2(new_n752_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n376_), .ZN(G1345gat));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n875_), .B2(new_n615_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n873_), .A2(KEYINPUT124), .A3(new_n716_), .A4(new_n874_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1346gat));
  OAI21_X1  g684(.A(G162gat), .B1(new_n875_), .B2(new_n679_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n626_), .A2(new_n366_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n875_), .B2(new_n887_), .ZN(G1347gat));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  INV_X1    g688(.A(new_n842_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n830_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n633_), .A2(new_n483_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n662_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n232_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n889_), .B1(new_n895_), .B2(new_n250_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n233_), .ZN(new_n897_));
  OAI211_X1 g696(.A(KEYINPUT62), .B(G169gat), .C1(new_n894_), .C2(new_n232_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(G1348gat));
  INV_X1    g698(.A(new_n894_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G176gat), .B1(new_n900_), .B2(new_n570_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n490_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n752_), .A2(new_n892_), .A3(new_n234_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1349gat));
  NOR2_X1   g703(.A1(new_n615_), .A2(new_n278_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n891_), .A2(new_n893_), .A3(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n892_), .A2(new_n615_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n873_), .A2(KEYINPUT125), .A3(new_n419_), .A4(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n242_), .ZN(new_n909_));
  AOI21_X1  g708(.A(KEYINPUT125), .B1(new_n902_), .B2(new_n907_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n906_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(KEYINPUT126), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n913_), .B(new_n906_), .C1(new_n909_), .C2(new_n910_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n894_), .B2(new_n679_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n626_), .A2(new_n281_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n894_), .B2(new_n917_), .ZN(G1351gat));
  NOR4_X1   g717(.A1(new_n361_), .A2(new_n419_), .A3(new_n482_), .A4(new_n659_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n873_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n232_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(new_n289_), .ZN(G1352gat));
  NOR2_X1   g721(.A1(new_n920_), .A2(new_n752_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(new_n287_), .ZN(G1353gat));
  AOI21_X1  g723(.A(new_n615_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  OAI21_X1  g725(.A(KEYINPUT127), .B1(new_n920_), .B2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n873_), .A2(new_n928_), .A3(new_n919_), .A4(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n930_), .B(new_n931_), .ZN(G1354gat));
  OAI21_X1  g731(.A(G218gat), .B1(new_n920_), .B2(new_n679_), .ZN(new_n933_));
  OR2_X1    g732(.A1(new_n598_), .A2(G218gat), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n920_), .B2(new_n934_), .ZN(G1355gat));
endmodule


