//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n968_, new_n969_, new_n971_, new_n972_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n980_,
    new_n981_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n991_, new_n992_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G85gat), .B(G92gat), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT6), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n208_), .B(new_n210_), .C1(KEYINPUT9), .C2(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n206_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(KEYINPUT69), .A2(KEYINPUT8), .ZN(new_n214_));
  INV_X1    g013(.A(G99gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT7), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n215_), .B(new_n203_), .C1(new_n216_), .C2(KEYINPUT66), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT7), .ZN(new_n220_));
  OR3_X1    g019(.A1(new_n217_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n218_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n210_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n207_), .B(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n214_), .B1(new_n225_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n210_), .A2(new_n224_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n230_), .B1(new_n222_), .B2(new_n221_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n214_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n227_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n213_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G57gat), .B(G64gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT11), .ZN(new_n238_));
  XOR2_X1   g037(.A(G71gat), .B(G78gat), .Z(new_n239_));
  OR2_X1    g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n235_), .B(KEYINPUT70), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT11), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n238_), .A2(new_n243_), .A3(new_n239_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n234_), .A2(KEYINPUT12), .A3(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n206_), .A2(new_n212_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n225_), .A2(new_n214_), .A3(new_n228_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n232_), .B1(new_n231_), .B2(new_n227_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n240_), .A2(new_n244_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n246_), .A2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n250_), .A2(new_n251_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT72), .B1(new_n254_), .B2(KEYINPUT12), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G230gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT64), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n234_), .A2(new_n245_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT72), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT12), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n253_), .A2(new_n255_), .A3(new_n257_), .A4(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT73), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n259_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n246_), .A2(new_n252_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n267_), .A2(KEYINPUT73), .A3(new_n257_), .A4(new_n261_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n258_), .A2(new_n252_), .A3(KEYINPUT71), .ZN(new_n269_));
  OR3_X1    g068(.A1(new_n234_), .A2(new_n245_), .A3(KEYINPUT71), .ZN(new_n270_));
  INV_X1    g069(.A(new_n257_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n264_), .A2(new_n268_), .A3(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G120gat), .B(G148gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT5), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G176gat), .B(G204gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n275_), .B(new_n276_), .Z(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n277_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n264_), .A2(new_n268_), .A3(new_n272_), .A4(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(KEYINPUT13), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT13), .B1(new_n278_), .B2(new_n280_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G231gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n245_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G1gat), .ZN(new_n288_));
  INV_X1    g087(.A(G8gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT14), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT75), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n292_), .B(KEYINPUT14), .C1(new_n288_), .C2(new_n289_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n291_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n295_), .A2(KEYINPUT76), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(KEYINPUT76), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(G1gat), .B(G8gat), .Z(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n296_), .A2(new_n299_), .A3(new_n297_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n287_), .B(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G127gat), .B(G155gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT16), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G183gat), .B(G211gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT17), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n304_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n309_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n304_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G232gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT34), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT35), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(new_n316_), .B2(KEYINPUT35), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G29gat), .B(G36gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G43gat), .B(G50gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n319_), .B1(new_n250_), .B2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(KEYINPUT15), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n234_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n317_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G190gat), .B(G218gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G134gat), .B(G162gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(KEYINPUT36), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n323_), .A2(new_n317_), .A3(new_n325_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n327_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n330_), .B(KEYINPUT36), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(new_n327_), .B2(new_n332_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT37), .B1(new_n334_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n337_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT37), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(new_n333_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n285_), .A2(new_n314_), .A3(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G127gat), .B(G134gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G113gat), .B(G120gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT31), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n347_), .B(KEYINPUT82), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT31), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT83), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n350_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n354_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G169gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT23), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(G183gat), .A3(G190gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n360_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT78), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT25), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(KEYINPUT79), .A3(G183gat), .ZN(new_n380_));
  INV_X1    g179(.A(G190gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT26), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT26), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G190gat), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(G183gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT25), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n379_), .A2(G183gat), .B1(KEYINPUT79), .B2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n370_), .B(new_n374_), .C1(new_n386_), .C2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n362_), .A2(KEYINPUT81), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n392_), .B1(new_n361_), .B2(KEYINPUT23), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n364_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  OR3_X1    g193(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n390_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n374_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n382_), .A2(new_n384_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n387_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n401_), .B2(KEYINPUT79), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n377_), .A2(KEYINPUT25), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n375_), .A2(KEYINPUT78), .ZN(new_n404_));
  OAI21_X1  g203(.A(G183gat), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n388_), .A2(KEYINPUT79), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n399_), .B1(new_n402_), .B2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n408_), .A2(new_n370_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n369_), .B1(new_n398_), .B2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G71gat), .B(G99gat), .ZN(new_n411_));
  INV_X1    g210(.A(G43gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n396_), .B1(new_n408_), .B2(new_n370_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n374_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT80), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n368_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n413_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421_));
  INV_X1    g220(.A(G15gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT30), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n414_), .A2(new_n420_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n414_), .B2(new_n420_), .ZN(new_n427_));
  OAI211_X1 g226(.A(KEYINPUT84), .B(new_n357_), .C1(new_n426_), .C2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n424_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n410_), .A2(new_n413_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n418_), .A2(new_n419_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n432_), .A2(new_n425_), .A3(new_n350_), .A4(new_n353_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n425_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT84), .B1(new_n435_), .B2(new_n357_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G22gat), .B(G50gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(G155gat), .A2(G162gat), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT85), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G155gat), .A2(G162gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n446_));
  NOR4_X1   g245(.A1(new_n446_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G141gat), .A2(G148gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT3), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT86), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G141gat), .A2(G148gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT2), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT2), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(G141gat), .A3(G148gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G141gat), .ZN(new_n457_));
  INV_X1    g256(.A(G148gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT3), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n456_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n445_), .B1(new_n451_), .B2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n449_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n446_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n448_), .A2(KEYINPUT86), .A3(new_n449_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n453_), .A2(new_n455_), .B1(new_n459_), .B2(KEYINPUT3), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(KEYINPUT87), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n444_), .B1(new_n462_), .B2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n443_), .B(KEYINPUT1), .Z(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n442_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n471_), .A2(new_n459_), .A3(new_n452_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT88), .B1(new_n469_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n444_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n466_), .A2(KEYINPUT87), .A3(new_n467_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT87), .B1(new_n466_), .B2(new_n467_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n471_), .A2(new_n459_), .A3(new_n452_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n473_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT29), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT28), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT28), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n481_), .A2(new_n485_), .A3(new_n482_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n439_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n485_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n488_));
  AOI211_X1 g287(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n473_), .C2(new_n480_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n438_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT21), .ZN(new_n491_));
  INV_X1    g290(.A(G204gat), .ZN(new_n492_));
  INV_X1    g291(.A(G197gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT89), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(G197gat), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n492_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(G197gat), .A2(G204gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n491_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(G218gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G211gat), .ZN(new_n501_));
  INV_X1    g300(.A(G211gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(G218gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n494_), .A2(new_n496_), .A3(new_n492_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n491_), .B1(G197gat), .B2(G204gat), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n499_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n497_), .A2(new_n498_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(KEYINPUT21), .A3(new_n504_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(G228gat), .B2(G233gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n513_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G78gat), .B(G106gat), .Z(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT90), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n508_), .A2(new_n510_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n482_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n521_));
  OAI211_X1 g320(.A(G228gat), .B(G233gat), .C1(new_n520_), .C2(new_n521_), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n514_), .A2(new_n516_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n516_), .B1(new_n514_), .B2(new_n522_), .ZN(new_n524_));
  OAI22_X1  g323(.A1(new_n487_), .A2(new_n490_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n514_), .A2(new_n522_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n515_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n484_), .A2(new_n486_), .A3(new_n439_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n438_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n514_), .A2(new_n516_), .A3(new_n522_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .A4(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n525_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G1gat), .B(G29gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(G85gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT0), .B(G57gat), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n534_), .B(new_n535_), .Z(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n473_), .A2(new_n480_), .A3(new_n351_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n477_), .A2(new_n479_), .A3(new_n347_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G225gat), .A2(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n538_), .A2(KEYINPUT4), .A3(new_n539_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT4), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n473_), .A2(new_n480_), .A3(new_n544_), .A4(new_n351_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n540_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n537_), .B(new_n542_), .C1(new_n543_), .C2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G8gat), .B(G36gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT18), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G64gat), .B(G92gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G226gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT20), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n360_), .B1(new_n394_), .B2(new_n367_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n365_), .A2(new_n395_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT92), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n365_), .A2(new_n561_), .A3(new_n395_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT25), .B(G183gat), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n385_), .A2(new_n564_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT93), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n365_), .A2(new_n561_), .A3(new_n395_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n561_), .B1(new_n365_), .B2(new_n395_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n565_), .B(KEYINPUT93), .C1(new_n567_), .C2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n558_), .B1(new_n566_), .B2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n556_), .B1(new_n571_), .B2(new_n511_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n512_), .B(new_n369_), .C1(new_n398_), .C2(new_n409_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n555_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n554_), .A2(new_n556_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n571_), .B2(new_n511_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n415_), .A2(new_n417_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n512_), .B1(new_n577_), .B2(new_n369_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n551_), .B1(new_n574_), .B2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n565_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n557_), .B1(new_n583_), .B2(new_n569_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT20), .B1(new_n584_), .B2(new_n512_), .ZN(new_n585_));
  AOI211_X1 g384(.A(new_n511_), .B(new_n368_), .C1(new_n415_), .C2(new_n417_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n554_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n551_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n575_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(new_n584_), .B2(new_n512_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n410_), .A2(new_n511_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n587_), .A2(new_n588_), .A3(new_n592_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n547_), .A2(new_n580_), .A3(new_n593_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n545_), .A2(new_n541_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n538_), .A2(KEYINPUT4), .A3(new_n539_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n595_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n599_), .A2(KEYINPUT94), .A3(KEYINPUT33), .A4(new_n536_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT94), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n602_), .B(new_n536_), .C1(new_n543_), .C2(new_n596_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n601_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n604_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n594_), .A2(new_n600_), .A3(new_n605_), .A4(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n602_), .B1(new_n543_), .B2(new_n596_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n537_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n603_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n588_), .A2(KEYINPUT32), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n585_), .A2(new_n586_), .A3(new_n554_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n557_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n556_), .B1(new_n520_), .B2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n555_), .B1(new_n614_), .B2(new_n591_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n611_), .B1(new_n612_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT95), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n574_), .A2(new_n579_), .A3(new_n611_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n616_), .B1(new_n619_), .B2(new_n617_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n610_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n532_), .B1(new_n607_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n580_), .A2(new_n593_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT27), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n573_), .B(KEYINPUT20), .C1(new_n512_), .C2(new_n584_), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n625_), .A2(new_n554_), .B1(new_n591_), .B2(new_n590_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n624_), .B1(new_n626_), .B2(new_n588_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n551_), .B1(new_n612_), .B2(new_n615_), .ZN(new_n628_));
  AOI22_X1  g427(.A1(new_n623_), .A2(new_n624_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n610_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n629_), .A2(new_n532_), .A3(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n437_), .B1(new_n622_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n628_), .A2(KEYINPUT27), .A3(new_n593_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT27), .B1(new_n580_), .B2(new_n593_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n633_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n587_), .A2(new_n588_), .A3(new_n592_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n588_), .B1(new_n587_), .B2(new_n592_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n624_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n628_), .A2(KEYINPUT27), .A3(new_n593_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(KEYINPUT96), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n636_), .A2(new_n641_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n525_), .A2(new_n531_), .A3(new_n603_), .A4(new_n609_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(new_n437_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n642_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n632_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n303_), .A2(new_n322_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n322_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n301_), .A2(new_n302_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n649_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n301_), .A2(new_n302_), .A3(new_n324_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n650_), .A2(new_n649_), .A3(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(G113gat), .B(G141gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT77), .ZN(new_n659_));
  XNOR2_X1  g458(.A(G169gat), .B(G197gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n657_), .B(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n344_), .A2(new_n648_), .A3(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT98), .Z(new_n664_));
  OR2_X1    g463(.A1(new_n610_), .A2(KEYINPUT99), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n610_), .A2(KEYINPUT99), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(new_n288_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT38), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n662_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n285_), .A2(new_n672_), .A3(new_n314_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n607_), .A2(new_n621_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n525_), .A2(new_n531_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n631_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n639_), .A2(KEYINPUT96), .A3(new_n640_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT96), .B1(new_n639_), .B2(new_n640_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n435_), .A2(new_n357_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT84), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n433_), .A3(new_n428_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n675_), .A2(new_n630_), .A3(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT97), .B1(new_n681_), .B2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n642_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n688_));
  AOI22_X1  g487(.A1(new_n678_), .A2(new_n437_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n339_), .A2(new_n333_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT100), .Z(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n689_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n673_), .A2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G1gat), .B1(new_n694_), .B2(new_n630_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n669_), .A2(new_n670_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n671_), .A2(new_n695_), .A3(new_n696_), .ZN(G1324gat));
  NAND3_X1  g496(.A1(new_n664_), .A2(new_n289_), .A3(new_n681_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G8gat), .B1(new_n694_), .B2(new_n642_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT39), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT40), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(G1325gat));
  OAI21_X1  g502(.A(G15gat), .B1(new_n694_), .B2(new_n437_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT101), .Z(new_n705_));
  OR2_X1    g504(.A1(new_n705_), .A2(KEYINPUT41), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(KEYINPUT41), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n664_), .A2(new_n422_), .A3(new_n685_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(G1326gat));
  XNOR2_X1  g508(.A(new_n532_), .B(KEYINPUT102), .ZN(new_n710_));
  INV_X1    g509(.A(G22gat), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT103), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n664_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n673_), .A2(new_n693_), .A3(new_n710_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G22gat), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT42), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n717_), .ZN(G1327gat));
  INV_X1    g517(.A(new_n690_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n314_), .ZN(new_n720_));
  NOR4_X1   g519(.A1(new_n689_), .A2(new_n285_), .A3(new_n672_), .A4(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G29gat), .B1(new_n721_), .B2(new_n610_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n314_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n285_), .A2(new_n672_), .A3(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n338_), .A2(new_n341_), .A3(KEYINPUT104), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(KEYINPUT43), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n687_), .A2(new_n688_), .ZN(new_n727_));
  AOI211_X1 g526(.A(new_n342_), .B(new_n726_), .C1(new_n727_), .C2(new_n632_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n726_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n648_), .B2(new_n343_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n724_), .B(KEYINPUT44), .C1(new_n728_), .C2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n726_), .B1(new_n689_), .B2(new_n342_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n648_), .A2(new_n343_), .A3(new_n729_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n736_), .A2(KEYINPUT105), .A3(KEYINPUT44), .A4(new_n724_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n724_), .B1(new_n728_), .B2(new_n730_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n733_), .A2(new_n737_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n668_), .A2(G29gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n722_), .B1(new_n740_), .B2(new_n741_), .ZN(G1328gat));
  INV_X1    g541(.A(G36gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n721_), .A2(new_n743_), .A3(new_n681_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT45), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n733_), .A2(new_n737_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n642_), .B1(new_n739_), .B2(new_n738_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n746_), .B1(new_n749_), .B2(G36gat), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT106), .B(new_n743_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n745_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  OAI211_X1 g553(.A(KEYINPUT46), .B(new_n745_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1329gat));
  NAND3_X1  g555(.A1(new_n740_), .A2(G43gat), .A3(new_n685_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n721_), .A2(new_n685_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n412_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g560(.A(G50gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n721_), .A2(new_n762_), .A3(new_n710_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n675_), .B1(new_n739_), .B2(new_n738_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n747_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G50gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n764_), .B1(new_n747_), .B2(new_n765_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n763_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT108), .B(new_n763_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1331gat));
  INV_X1    g572(.A(G57gat), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n693_), .A2(new_n672_), .A3(new_n285_), .A4(new_n723_), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n775_), .A2(KEYINPUT109), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(KEYINPUT109), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n774_), .B1(new_n778_), .B2(new_n610_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n689_), .A2(new_n662_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n284_), .A2(new_n314_), .A3(new_n343_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n782_), .A2(G57gat), .A3(new_n667_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n779_), .A2(new_n783_), .ZN(G1332gat));
  OR3_X1    g583(.A1(new_n782_), .A2(G64gat), .A3(new_n642_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n776_), .A2(new_n681_), .A3(new_n777_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT48), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(G64gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(G64gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT110), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(new_n785_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1333gat));
  OR3_X1    g593(.A1(new_n782_), .A2(G71gat), .A3(new_n437_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n778_), .A2(new_n685_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(G71gat), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(KEYINPUT49), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(KEYINPUT49), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(G1334gat));
  INV_X1    g599(.A(G78gat), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n780_), .A2(new_n801_), .A3(new_n781_), .A4(new_n710_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n778_), .A2(new_n710_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(G78gat), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n804_), .A2(KEYINPUT50), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(KEYINPUT50), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n802_), .B1(new_n805_), .B2(new_n806_), .ZN(G1335gat));
  NOR2_X1   g606(.A1(new_n284_), .A2(new_n720_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n780_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(G85gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n811_), .A3(new_n668_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n285_), .A2(new_n672_), .A3(new_n314_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n610_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n812_), .B1(new_n816_), .B2(new_n811_), .ZN(G1336gat));
  NOR3_X1   g616(.A1(new_n809_), .A2(G92gat), .A3(new_n642_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n814_), .A2(new_n681_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(G92gat), .B2(new_n819_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT111), .Z(G1337gat));
  AOI21_X1  g620(.A(new_n215_), .B1(new_n814_), .B2(new_n685_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n685_), .A2(new_n202_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n810_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n824_), .B(new_n825_), .ZN(G1338gat));
  NAND3_X1  g625(.A1(new_n810_), .A2(new_n203_), .A3(new_n532_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n814_), .A2(new_n532_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n828_), .A2(G106gat), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n828_), .B2(G106gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n827_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g632(.A(G113gat), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n681_), .A2(new_n667_), .A3(new_n437_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837_));
  INV_X1    g636(.A(new_n655_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n651_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n650_), .A2(KEYINPUT117), .A3(new_n655_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n649_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n840_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n650_), .A2(new_n652_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n661_), .B1(new_n844_), .B2(new_n649_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n654_), .A2(new_n656_), .A3(new_n661_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n846_), .A2(KEYINPUT118), .A3(new_n847_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n852_), .A2(new_n280_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n264_), .A2(new_n268_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n253_), .A2(new_n255_), .A3(new_n261_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n271_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n854_), .B2(new_n262_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n277_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n853_), .B1(new_n859_), .B2(KEYINPUT56), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n262_), .A2(new_n854_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n257_), .B1(new_n267_), .B2(new_n261_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n264_), .A2(new_n268_), .A3(new_n854_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n279_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT56), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n836_), .B1(new_n860_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n859_), .A2(KEYINPUT56), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n865_), .A2(new_n866_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n869_), .A2(KEYINPUT58), .A3(new_n870_), .A4(new_n853_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n868_), .A2(new_n343_), .A3(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n278_), .A2(new_n280_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n852_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n874_), .B2(new_n852_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n873_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n662_), .A2(new_n280_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n662_), .A2(new_n280_), .A3(KEYINPUT115), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n859_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT116), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n866_), .B1(new_n865_), .B2(new_n886_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n884_), .A2(new_n885_), .A3(new_n887_), .ZN(new_n888_));
  OAI22_X1  g687(.A1(new_n879_), .A2(new_n888_), .B1(KEYINPUT120), .B2(new_n690_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n872_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  OAI221_X1 g690(.A(KEYINPUT57), .B1(KEYINPUT120), .B2(new_n690_), .C1(new_n879_), .C2(new_n888_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n723_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n723_), .A2(new_n672_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT114), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n284_), .A3(new_n342_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT54), .Z(new_n897_));
  OAI211_X1 g696(.A(new_n675_), .B(new_n835_), .C1(new_n893_), .C2(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n834_), .B1(new_n898_), .B2(new_n672_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  OAI211_X1 g700(.A(KEYINPUT121), .B(new_n834_), .C1(new_n898_), .C2(new_n672_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n897_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n891_), .A2(new_n892_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n723_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n905_), .A2(KEYINPUT59), .A3(new_n675_), .A4(new_n835_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n898_), .A2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n672_), .A2(new_n834_), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n901_), .A2(new_n902_), .B1(new_n909_), .B2(new_n910_), .ZN(G1340gat));
  INV_X1    g710(.A(G120gat), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(KEYINPUT60), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n914_));
  AOI21_X1  g713(.A(G120gat), .B1(new_n285_), .B2(new_n914_), .ZN(new_n915_));
  OR3_X1    g714(.A1(new_n898_), .A2(new_n913_), .A3(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n284_), .B1(new_n906_), .B2(new_n908_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n912_), .ZN(G1341gat));
  AOI21_X1  g717(.A(new_n314_), .B1(new_n906_), .B2(new_n908_), .ZN(new_n919_));
  INV_X1    g718(.A(G127gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n723_), .A2(new_n920_), .ZN(new_n921_));
  OAI22_X1  g720(.A1(new_n919_), .A2(new_n920_), .B1(new_n898_), .B2(new_n921_), .ZN(G1342gat));
  XNOR2_X1  g721(.A(KEYINPUT122), .B(G134gat), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n342_), .A2(new_n923_), .ZN(new_n924_));
  OR2_X1    g723(.A1(new_n898_), .A2(new_n691_), .ZN(new_n925_));
  INV_X1    g724(.A(G134gat), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n909_), .A2(new_n924_), .B1(new_n925_), .B2(new_n926_), .ZN(G1343gat));
  NOR3_X1   g726(.A1(new_n681_), .A2(new_n667_), .A3(new_n675_), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n437_), .B(new_n928_), .C1(new_n893_), .C2(new_n897_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(new_n672_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(new_n457_), .ZN(G1344gat));
  NOR2_X1   g730(.A1(new_n929_), .A2(new_n284_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(new_n458_), .ZN(G1345gat));
  NOR2_X1   g732(.A1(new_n929_), .A2(new_n314_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(KEYINPUT61), .B(G155gat), .ZN(new_n935_));
  XOR2_X1   g734(.A(new_n934_), .B(new_n935_), .Z(G1346gat));
  INV_X1    g735(.A(G162gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n937_), .B1(new_n929_), .B2(new_n691_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n343_), .A2(G162gat), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(KEYINPUT123), .ZN(new_n940_));
  NAND4_X1  g739(.A1(new_n905_), .A2(new_n437_), .A3(new_n928_), .A4(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n938_), .A2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(KEYINPUT124), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n938_), .A2(new_n941_), .A3(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n945_), .ZN(G1347gat));
  INV_X1    g745(.A(G169gat), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n668_), .A2(new_n437_), .A3(new_n642_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(new_n710_), .ZN(new_n950_));
  OAI211_X1 g749(.A(new_n662_), .B(new_n950_), .C1(new_n893_), .C2(new_n897_), .ZN(new_n951_));
  OAI211_X1 g750(.A(KEYINPUT62), .B(new_n947_), .C1(new_n951_), .C2(KEYINPUT22), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  OAI21_X1  g752(.A(KEYINPUT62), .B1(new_n951_), .B2(KEYINPUT22), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n951_), .A2(KEYINPUT62), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n955_), .A2(new_n947_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n953_), .B1(new_n954_), .B2(new_n956_), .ZN(G1348gat));
  NAND3_X1  g756(.A1(new_n905_), .A2(KEYINPUT125), .A3(new_n675_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n893_), .A2(new_n897_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n960_), .B2(new_n532_), .ZN(new_n961_));
  INV_X1    g760(.A(G176gat), .ZN(new_n962_));
  NOR3_X1   g761(.A1(new_n949_), .A2(new_n284_), .A3(new_n962_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n958_), .A2(new_n961_), .A3(new_n963_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n905_), .A2(new_n950_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n962_), .B1(new_n965_), .B2(new_n284_), .ZN(new_n966_));
  AND2_X1   g765(.A1(new_n964_), .A2(new_n966_), .ZN(G1349gat));
  NOR3_X1   g766(.A1(new_n965_), .A2(new_n564_), .A3(new_n314_), .ZN(new_n968_));
  NAND4_X1  g767(.A1(new_n958_), .A2(new_n961_), .A3(new_n723_), .A4(new_n948_), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n968_), .B1(new_n969_), .B2(new_n387_), .ZN(G1350gat));
  OAI21_X1  g769(.A(G190gat), .B1(new_n965_), .B2(new_n342_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n692_), .A2(new_n385_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n965_), .B2(new_n972_), .ZN(G1351gat));
  NOR3_X1   g772(.A1(new_n642_), .A2(new_n675_), .A3(new_n610_), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n905_), .A2(new_n437_), .A3(new_n974_), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n493_), .B1(new_n975_), .B2(new_n672_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n960_), .A2(new_n685_), .ZN(new_n977_));
  NAND4_X1  g776(.A1(new_n977_), .A2(G197gat), .A3(new_n662_), .A4(new_n974_), .ZN(new_n978_));
  AND2_X1   g777(.A1(new_n976_), .A2(new_n978_), .ZN(G1352gat));
  OAI21_X1  g778(.A(G204gat), .B1(new_n975_), .B2(new_n284_), .ZN(new_n980_));
  NAND4_X1  g779(.A1(new_n977_), .A2(new_n492_), .A3(new_n285_), .A4(new_n974_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n980_), .A2(new_n981_), .ZN(G1353gat));
  INV_X1    g781(.A(KEYINPUT63), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n983_), .A2(new_n502_), .ZN(new_n984_));
  XNOR2_X1  g783(.A(new_n984_), .B(KEYINPUT127), .ZN(new_n985_));
  OAI21_X1  g784(.A(new_n723_), .B1(new_n983_), .B2(new_n502_), .ZN(new_n986_));
  XNOR2_X1  g785(.A(new_n986_), .B(KEYINPUT126), .ZN(new_n987_));
  OR3_X1    g786(.A1(new_n975_), .A2(new_n985_), .A3(new_n987_), .ZN(new_n988_));
  OAI21_X1  g787(.A(new_n985_), .B1(new_n975_), .B2(new_n987_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n988_), .A2(new_n989_), .ZN(G1354gat));
  OAI21_X1  g789(.A(G218gat), .B1(new_n975_), .B2(new_n342_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n692_), .A2(new_n500_), .ZN(new_n992_));
  OAI21_X1  g791(.A(new_n991_), .B1(new_n975_), .B2(new_n992_), .ZN(G1355gat));
endmodule


