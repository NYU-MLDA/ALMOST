//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n949_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G29gat), .B(G36gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G43gat), .B(G50gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n203_), .A2(new_n205_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT75), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G1gat), .B(G8gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT74), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(KEYINPUT74), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216_));
  INV_X1    g015(.A(G8gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n215_), .A2(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n213_), .A2(new_n218_), .A3(new_n216_), .A4(new_n214_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n211_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT76), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n211_), .A2(new_n222_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT77), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n223_), .A2(KEYINPUT76), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n223_), .A2(KEYINPUT76), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n225_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT77), .B1(new_n234_), .B2(new_n229_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n209_), .B(KEYINPUT15), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n238_), .A2(new_n222_), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n239_), .B(KEYINPUT78), .Z(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(new_n224_), .A3(new_n229_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G113gat), .B(G141gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G169gat), .B(G197gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT79), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n236_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n242_), .A2(KEYINPUT79), .A3(new_n246_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT10), .B(G99gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G106gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G85gat), .B(G92gat), .Z(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT9), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G99gat), .A2(G106gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT6), .ZN(new_n262_));
  INV_X1    g061(.A(G85gat), .ZN(new_n263_));
  INV_X1    g062(.A(G92gat), .ZN(new_n264_));
  OR3_X1    g063(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT9), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n260_), .A2(new_n262_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n258_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n270_));
  OR3_X1    g069(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n262_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n259_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n259_), .A2(KEYINPUT66), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT8), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n273_), .B(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n269_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n237_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G232gat), .A2(G233gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n280_), .B(KEYINPUT34), .Z(new_n281_));
  XOR2_X1   g080(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(new_n267_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n209_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n281_), .A2(new_n282_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n279_), .A2(new_n287_), .A3(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n238_), .B1(new_n269_), .B2(new_n277_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n288_), .B1(new_n291_), .B2(new_n286_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G190gat), .B(G218gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(G134gat), .B(G162gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT36), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT72), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n290_), .A2(new_n292_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT73), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n290_), .A2(new_n292_), .A3(new_n301_), .A4(new_n298_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n290_), .A2(new_n292_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n295_), .A2(new_n296_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n297_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G71gat), .B(G99gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(G43gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT30), .ZN(new_n311_));
  NOR2_X1   g110(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n312_));
  INV_X1    g111(.A(G169gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT23), .ZN(new_n318_));
  INV_X1    g117(.A(G183gat), .ZN(new_n319_));
  INV_X1    g118(.A(G190gat), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT81), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n316_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n324_), .B(new_n325_), .C1(G183gat), .C2(G190gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT81), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n322_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n319_), .A2(KEYINPUT25), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(G183gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n320_), .A2(KEYINPUT26), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT26), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(G190gat), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n329_), .A2(new_n331_), .A3(new_n332_), .A4(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NOR3_X1   g136(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n339_), .A2(KEYINPUT24), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n338_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT25), .B(G183gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT26), .B(G190gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(KEYINPUT80), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n337_), .A2(new_n318_), .A3(new_n343_), .A4(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n328_), .A2(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n311_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n311_), .A2(new_n348_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G227gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(G15gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n349_), .A2(new_n354_), .A3(new_n350_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n359_), .A2(KEYINPUT31), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(KEYINPUT31), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G113gat), .B(G120gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n365_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n360_), .A2(new_n367_), .A3(new_n361_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370_));
  INV_X1    g169(.A(G228gat), .ZN(new_n371_));
  INV_X1    g170(.A(G233gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT87), .ZN(new_n374_));
  INV_X1    g173(.A(G197gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n376_));
  INV_X1    g175(.A(G204gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(KEYINPUT86), .A2(G204gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n375_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(G197gat), .A2(G204gat), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n374_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(KEYINPUT86), .A2(G204gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(KEYINPUT86), .A2(G204gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(G197gat), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n381_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(KEYINPUT87), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G211gat), .B(G218gat), .Z(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT21), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT21), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n378_), .A2(new_n375_), .A3(new_n379_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT21), .B1(new_n375_), .B2(new_n377_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n389_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n388_), .A2(new_n391_), .B1(new_n393_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT83), .ZN(new_n400_));
  AND2_X1   g199(.A1(G155gat), .A2(G162gat), .ZN(new_n401_));
  NOR2_X1   g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n401_), .A2(new_n402_), .A3(KEYINPUT1), .ZN(new_n403_));
  INV_X1    g202(.A(G141gat), .ZN(new_n404_));
  INV_X1    g203(.A(G148gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G141gat), .A2(G148gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n400_), .B1(new_n403_), .B2(new_n409_), .ZN(new_n410_));
  OR2_X1    g209(.A1(G155gat), .A2(G162gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT1), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n408_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(G141gat), .A2(G148gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n414_), .A2(new_n417_), .A3(KEYINPUT83), .A4(new_n407_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n410_), .A2(new_n418_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n401_), .A2(new_n402_), .A3(KEYINPUT84), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n415_), .A2(KEYINPUT2), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT3), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n416_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT2), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n408_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n424_), .A2(new_n426_), .A3(new_n428_), .A4(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n423_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n399_), .B1(new_n419_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n373_), .B1(new_n398_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n419_), .A2(new_n431_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT29), .ZN(new_n435_));
  INV_X1    g234(.A(new_n373_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n380_), .A2(new_n374_), .A3(new_n381_), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT87), .B1(new_n385_), .B2(new_n386_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n391_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n397_), .A2(new_n393_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n435_), .A2(new_n436_), .A3(new_n441_), .ZN(new_n442_));
  AOI211_X1 g241(.A(KEYINPUT88), .B(new_n370_), .C1(new_n433_), .C2(new_n442_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n398_), .A2(new_n432_), .A3(new_n373_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n436_), .B1(new_n435_), .B2(new_n441_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n370_), .B(KEYINPUT88), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G22gat), .B(G50gat), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n410_), .A2(new_n418_), .B1(new_n423_), .B2(new_n430_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(new_n399_), .ZN(new_n452_));
  AND4_X1   g251(.A1(new_n399_), .A2(new_n419_), .A3(new_n431_), .A4(new_n450_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n449_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n450_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n455_), .B1(new_n434_), .B2(KEYINPUT29), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n451_), .A2(new_n399_), .A3(new_n450_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n448_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  OR3_X1    g258(.A1(new_n443_), .A2(new_n447_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n370_), .A2(KEYINPUT89), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n433_), .A2(new_n442_), .A3(new_n461_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n459_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT90), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n463_), .A2(new_n459_), .A3(KEYINPUT90), .A4(new_n464_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G57gat), .B(G85gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT97), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(G1gat), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n470_), .A2(KEYINPUT97), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(KEYINPUT97), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n202_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n477_));
  INV_X1    g276(.A(G29gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n476_), .B(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n434_), .A2(new_n367_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n451_), .A2(new_n365_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(KEYINPUT4), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G225gat), .A2(G233gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n365_), .B1(new_n419_), .B2(new_n431_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT4), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n484_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(KEYINPUT95), .A3(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n481_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT95), .B1(new_n483_), .B2(new_n487_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n480_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n483_), .A2(new_n487_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT95), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n479_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n476_), .B(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n495_), .A2(new_n497_), .A3(new_n489_), .A4(new_n488_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n492_), .A2(KEYINPUT99), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT99), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n500_), .B(new_n480_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n460_), .A2(new_n469_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT27), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n439_), .A2(new_n440_), .A3(new_n328_), .A4(new_n347_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n316_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n326_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n325_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n338_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n335_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT92), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n339_), .A2(new_n512_), .A3(KEYINPUT24), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n512_), .B1(new_n339_), .B2(KEYINPUT24), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n341_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n506_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n390_), .B1(new_n382_), .B2(new_n387_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G211gat), .B(G218gat), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n383_), .A2(new_n384_), .A3(G197gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(new_n395_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT21), .B1(new_n385_), .B2(new_n386_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n516_), .B1(new_n517_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n504_), .A2(new_n523_), .A3(KEYINPUT20), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G226gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT19), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT91), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT93), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n335_), .A2(new_n336_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT80), .B1(new_n344_), .B2(new_n345_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n343_), .A2(new_n318_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n532_), .A2(new_n533_), .B1(new_n327_), .B2(new_n322_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT94), .B1(new_n534_), .B2(new_n398_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT20), .ZN(new_n536_));
  INV_X1    g335(.A(new_n516_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n398_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n526_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT94), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n441_), .A2(new_n540_), .A3(new_n348_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n535_), .A2(new_n538_), .A3(new_n539_), .A4(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n524_), .A2(new_n543_), .A3(new_n527_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G8gat), .B(G36gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT18), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G64gat), .B(G92gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  NAND4_X1  g347(.A1(new_n529_), .A2(new_n542_), .A3(new_n544_), .A4(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT101), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n524_), .A2(new_n527_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n535_), .A2(new_n541_), .A3(new_n538_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(new_n539_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n548_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n549_), .A2(new_n550_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n542_), .A2(new_n544_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n543_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(KEYINPUT101), .A3(new_n548_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n503_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n554_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(new_n503_), .A3(new_n549_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n502_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n469_), .A2(new_n460_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n484_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n481_), .A2(new_n482_), .A3(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT98), .B1(new_n497_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT98), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n481_), .A2(new_n482_), .A3(new_n566_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n480_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n483_), .B(new_n484_), .C1(KEYINPUT4), .C2(new_n481_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n568_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n561_), .A2(new_n549_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n498_), .A2(KEYINPUT33), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n488_), .A2(new_n489_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT33), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n497_), .A4(new_n495_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n548_), .A2(KEYINPUT32), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n558_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n553_), .A2(KEYINPUT32), .A3(new_n548_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n499_), .A2(new_n501_), .A3(new_n582_), .A4(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n565_), .B1(new_n580_), .B2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n564_), .B1(new_n585_), .B2(KEYINPUT100), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT100), .ZN(new_n587_));
  AOI211_X1 g386(.A(new_n587_), .B(new_n565_), .C1(new_n580_), .C2(new_n584_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n369_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n499_), .A2(new_n501_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n369_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n560_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n562_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n565_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n591_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n308_), .B1(new_n589_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n222_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT67), .B(G71gat), .ZN(new_n599_));
  INV_X1    g398(.A(G78gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G57gat), .B(G64gat), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n602_), .A2(KEYINPUT11), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n602_), .A2(KEYINPUT11), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n601_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n598_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT17), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT16), .ZN(new_n611_));
  XOR2_X1   g410(.A(G183gat), .B(G211gat), .Z(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n608_), .A2(new_n609_), .A3(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(KEYINPUT17), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n608_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT70), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n284_), .A2(new_n607_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n607_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT12), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n618_), .B1(new_n278_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT64), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n284_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n620_), .B1(new_n626_), .B2(new_n619_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n622_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n619_), .B1(new_n277_), .B2(new_n267_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n624_), .B1(new_n629_), .B2(new_n618_), .ZN(new_n630_));
  XOR2_X1   g429(.A(G120gat), .B(G148gat), .Z(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n628_), .A2(new_n630_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n636_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n617_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n639_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(KEYINPUT70), .A3(new_n637_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT13), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(new_n642_), .A3(KEYINPUT13), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AND4_X1   g447(.A1(new_n253_), .A2(new_n596_), .A3(new_n616_), .A4(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n202_), .B1(new_n649_), .B2(new_n590_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n589_), .A2(new_n595_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n253_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT37), .B1(new_n303_), .B2(new_n306_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n303_), .A2(KEYINPUT37), .A3(new_n306_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n616_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n654_), .A2(new_n660_), .A3(new_n648_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n590_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(G1gat), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n650_), .B1(new_n665_), .B2(KEYINPUT38), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n665_), .A2(KEYINPUT103), .A3(KEYINPUT38), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT38), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n664_), .B2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n667_), .B2(new_n670_), .ZN(G1324gat));
  INV_X1    g470(.A(new_n593_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n661_), .A2(new_n217_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n649_), .A2(new_n672_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(G8gat), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(KEYINPUT39), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(KEYINPUT39), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(G1325gat));
  INV_X1    g479(.A(new_n369_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n353_), .B1(new_n649_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT41), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n661_), .A2(new_n353_), .A3(new_n681_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1326gat));
  INV_X1    g484(.A(G22gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n649_), .B2(new_n565_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT42), .Z(new_n688_));
  NAND3_X1  g487(.A1(new_n661_), .A2(new_n686_), .A3(new_n565_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1327gat));
  NOR3_X1   g489(.A1(new_n647_), .A2(new_n307_), .A3(new_n616_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n654_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n478_), .B1(new_n692_), .B2(new_n662_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n647_), .A2(new_n252_), .A3(new_n616_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n651_), .B2(new_n658_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n303_), .A2(KEYINPUT37), .A3(new_n306_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n655_), .ZN(new_n698_));
  AOI211_X1 g497(.A(KEYINPUT43), .B(new_n698_), .C1(new_n589_), .C2(new_n595_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n696_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT44), .B(new_n694_), .C1(new_n696_), .C2(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n590_), .A2(G29gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n693_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT104), .Z(G1328gat));
  NOR2_X1   g506(.A1(new_n593_), .A2(G36gat), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n652_), .A2(new_n653_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT102), .B1(new_n651_), .B2(new_n253_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n691_), .B(new_n708_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n702_), .A2(new_n672_), .A3(new_n703_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(new_n715_), .A3(G36gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n714_), .B2(G36gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT46), .B(new_n713_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1329gat));
  NOR2_X1   g521(.A1(new_n692_), .A2(new_n369_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n681_), .A2(G43gat), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n723_), .A2(G43gat), .B1(new_n704_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g525(.A1(new_n692_), .A2(new_n594_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(G50gat), .ZN(new_n728_));
  INV_X1    g527(.A(new_n704_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n565_), .A2(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n729_), .B2(new_n730_), .ZN(G1331gat));
  NOR2_X1   g530(.A1(new_n648_), .A2(new_n253_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n732_), .A2(new_n651_), .A3(new_n660_), .ZN(new_n733_));
  INV_X1    g532(.A(G57gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n590_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(new_n616_), .A3(new_n596_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT107), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n737_), .A2(new_n590_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n738_), .B2(new_n734_), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n733_), .A2(new_n740_), .A3(new_n672_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n672_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(G64gat), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n742_), .B2(G64gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n733_), .A2(new_n747_), .A3(new_n681_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n737_), .A2(new_n681_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G71gat), .ZN(new_n751_));
  AOI211_X1 g550(.A(KEYINPUT49), .B(new_n747_), .C1(new_n737_), .C2(new_n681_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1334gat));
  NAND3_X1  g552(.A1(new_n733_), .A2(new_n600_), .A3(new_n565_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n737_), .A2(new_n565_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G78gat), .ZN(new_n757_));
  AOI211_X1 g556(.A(KEYINPUT50), .B(new_n600_), .C1(new_n737_), .C2(new_n565_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1335gat));
  OR2_X1    g558(.A1(new_n696_), .A2(new_n699_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n732_), .A2(new_n659_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n763_), .A2(new_n263_), .A3(new_n662_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n732_), .A2(new_n651_), .A3(new_n308_), .A4(new_n659_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT109), .ZN(new_n766_));
  AOI21_X1  g565(.A(G85gat), .B1(new_n766_), .B2(new_n590_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n768_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n764_), .B1(new_n769_), .B2(new_n770_), .ZN(G1336gat));
  NAND3_X1  g570(.A1(new_n766_), .A2(new_n264_), .A3(new_n672_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G92gat), .B1(new_n763_), .B2(new_n593_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1337gat));
  NAND3_X1  g573(.A1(new_n766_), .A2(new_n681_), .A3(new_n256_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n760_), .A2(new_n681_), .A3(new_n762_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(G99gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G99gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n781_), .A2(KEYINPUT112), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n780_), .B(new_n782_), .ZN(G1338gat));
  NAND3_X1  g582(.A1(new_n766_), .A2(new_n257_), .A3(new_n565_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n760_), .A2(new_n565_), .A3(new_n762_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n785_), .A2(new_n786_), .A3(G106gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n785_), .B2(G106gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g589(.A(G113gat), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n672_), .A2(new_n662_), .A3(new_n369_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n246_), .B1(new_n234_), .B2(new_n230_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(KEYINPUT117), .B(new_n246_), .C1(new_n234_), .C2(new_n230_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n240_), .A2(new_n224_), .A3(new_n230_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n249_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT118), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n249_), .A2(new_n798_), .A3(new_n801_), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n800_), .A2(new_n802_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n622_), .A2(KEYINPUT55), .A3(new_n625_), .A4(new_n627_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT116), .ZN(new_n806_));
  XNOR2_X1  g605(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n628_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n622_), .A2(new_n627_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n624_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n806_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n804_), .B1(new_n812_), .B2(new_n636_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n805_), .B(new_n814_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n808_), .A2(new_n810_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n636_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT56), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n813_), .A2(new_n818_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n250_), .A2(new_n251_), .A3(new_n637_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n803_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n308_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n800_), .A2(new_n802_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n643_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n815_), .A2(new_n816_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT56), .B1(new_n826_), .B2(new_n635_), .ZN(new_n827_));
  AOI211_X1 g626(.A(new_n804_), .B(new_n636_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n250_), .A2(new_n251_), .A3(new_n637_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n825_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT57), .B1(new_n831_), .B2(new_n307_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n823_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n817_), .B2(KEYINPUT56), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT119), .B(new_n804_), .C1(new_n812_), .C2(new_n636_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n818_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n638_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT58), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n837_), .A2(KEYINPUT58), .A3(new_n838_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n658_), .A3(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n616_), .B1(new_n833_), .B2(new_n842_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n844_));
  NAND4_X1  g643(.A1(new_n648_), .A2(new_n660_), .A3(KEYINPUT114), .A4(new_n252_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n698_), .A2(new_n645_), .A3(new_n616_), .A4(new_n646_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n253_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n844_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n845_), .A2(new_n848_), .A3(new_n844_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n594_), .B(new_n792_), .C1(new_n843_), .C2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n791_), .B1(new_n853_), .B2(new_n252_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(KEYINPUT120), .B(new_n791_), .C1(new_n853_), .C2(new_n252_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n853_), .A2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n822_), .B1(new_n821_), .B2(new_n308_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n831_), .A2(KEYINPUT57), .A3(new_n307_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n841_), .A2(new_n658_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n860_), .B(new_n861_), .C1(new_n862_), .C2(new_n839_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n659_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n845_), .A2(new_n848_), .A3(new_n844_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n849_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n565_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(KEYINPUT59), .A3(new_n792_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n859_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n253_), .A2(G113gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT121), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n856_), .A2(new_n857_), .B1(new_n869_), .B2(new_n871_), .ZN(G1340gat));
  NOR2_X1   g671(.A1(new_n648_), .A2(KEYINPUT60), .ZN(new_n873_));
  INV_X1    g672(.A(G120gat), .ZN(new_n874_));
  MUX2_X1   g673(.A(KEYINPUT60), .B(new_n873_), .S(new_n874_), .Z(new_n875_));
  NAND3_X1  g674(.A1(new_n867_), .A2(new_n792_), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n867_), .A2(KEYINPUT122), .A3(new_n792_), .A4(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n648_), .B1(new_n859_), .B2(new_n868_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n874_), .ZN(G1341gat));
  AOI21_X1  g681(.A(new_n659_), .B1(new_n859_), .B2(new_n868_), .ZN(new_n883_));
  INV_X1    g682(.A(G127gat), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n616_), .A2(new_n884_), .ZN(new_n885_));
  OAI22_X1  g684(.A1(new_n883_), .A2(new_n884_), .B1(new_n853_), .B2(new_n885_), .ZN(G1342gat));
  AOI21_X1  g685(.A(new_n698_), .B1(new_n859_), .B2(new_n868_), .ZN(new_n887_));
  INV_X1    g686(.A(G134gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n308_), .A2(new_n888_), .ZN(new_n889_));
  OAI22_X1  g688(.A1(new_n887_), .A2(new_n888_), .B1(new_n853_), .B2(new_n889_), .ZN(G1343gat));
  NAND2_X1  g689(.A1(new_n864_), .A2(new_n866_), .ZN(new_n891_));
  NOR4_X1   g690(.A1(new_n672_), .A2(new_n681_), .A3(new_n594_), .A4(new_n662_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n252_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(new_n404_), .ZN(G1344gat));
  NOR2_X1   g694(.A1(new_n893_), .A2(new_n648_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(new_n405_), .ZN(G1345gat));
  OAI211_X1 g696(.A(new_n616_), .B(new_n892_), .C1(new_n843_), .C2(new_n852_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT123), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n891_), .A2(new_n900_), .A3(new_n616_), .A4(new_n892_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT61), .B(G155gat), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n899_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n899_), .B2(new_n901_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1346gat));
  OAI21_X1  g704(.A(G162gat), .B1(new_n893_), .B2(new_n698_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n307_), .A2(G162gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n893_), .B2(new_n907_), .ZN(G1347gat));
  NAND2_X1  g707(.A1(new_n591_), .A2(new_n672_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n867_), .A2(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT22), .B(G169gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(new_n253_), .A3(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n909_), .A2(new_n252_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT124), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n867_), .A2(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n914_), .B1(new_n917_), .B2(G169gat), .ZN(new_n918_));
  AOI211_X1 g717(.A(KEYINPUT62), .B(new_n313_), .C1(new_n867_), .C2(new_n916_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n913_), .B1(new_n918_), .B2(new_n919_), .ZN(G1348gat));
  NAND3_X1  g719(.A1(new_n867_), .A2(new_n647_), .A3(new_n910_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT125), .B(G176gat), .Z(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1349gat));
  NAND3_X1  g722(.A1(new_n867_), .A2(new_n616_), .A3(new_n910_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n344_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(new_n319_), .B2(new_n924_), .ZN(G1350gat));
  NAND3_X1  g725(.A1(new_n911_), .A2(new_n345_), .A3(new_n308_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n867_), .A2(new_n658_), .A3(new_n910_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929_));
  AND3_X1   g728(.A1(new_n928_), .A2(new_n929_), .A3(G190gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n928_), .B2(G190gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n927_), .B1(new_n930_), .B2(new_n931_), .ZN(G1351gat));
  AND3_X1   g731(.A1(new_n672_), .A2(new_n502_), .A3(new_n369_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n891_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n252_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n375_), .ZN(G1352gat));
  AOI211_X1 g735(.A(new_n648_), .B(new_n934_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n891_), .A2(new_n933_), .ZN(new_n938_));
  AOI21_X1  g737(.A(G204gat), .B1(new_n938_), .B2(new_n647_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n937_), .A2(new_n939_), .ZN(G1353gat));
  OR2_X1    g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  NAND2_X1  g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  AND4_X1   g741(.A1(new_n616_), .A2(new_n938_), .A3(new_n941_), .A4(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n941_), .B1(new_n938_), .B2(new_n616_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1354gat));
  AND3_X1   g744(.A1(new_n938_), .A2(G218gat), .A3(new_n658_), .ZN(new_n946_));
  AND3_X1   g745(.A1(new_n891_), .A2(new_n308_), .A3(new_n933_), .ZN(new_n947_));
  OR2_X1    g746(.A1(new_n947_), .A2(KEYINPUT127), .ZN(new_n948_));
  AOI21_X1  g747(.A(G218gat), .B1(new_n947_), .B2(KEYINPUT127), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n946_), .B1(new_n948_), .B2(new_n949_), .ZN(G1355gat));
endmodule


