//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_;
  OR2_X1    g000(.A1(G197gat), .A2(G204gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G197gat), .A2(G204gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(KEYINPUT21), .A3(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT21), .ZN(new_n205_));
  AND2_X1   g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n204_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NOR3_X1   g009(.A1(new_n206_), .A2(new_n207_), .A3(new_n205_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G211gat), .B(G218gat), .Z(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n215_), .B1(KEYINPUT1), .B2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(KEYINPUT1), .B2(new_n216_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G141gat), .B(G148gat), .Z(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  INV_X1    g020(.A(G141gat), .ZN(new_n222_));
  INV_X1    g021(.A(G148gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n224_), .A2(new_n226_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n215_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n230_), .A2(new_n216_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n220_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT29), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n214_), .B1(new_n234_), .B2(KEYINPUT88), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G228gat), .A2(G233gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT87), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n214_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT86), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n210_), .A2(new_n213_), .A3(KEYINPUT87), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT88), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n242_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT87), .B1(new_n210_), .B2(new_n213_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n237_), .A2(new_n241_), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n245_), .A2(new_n237_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n234_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n238_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G78gat), .B(G106gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(KEYINPUT89), .A3(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G22gat), .B(G50gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT28), .B1(new_n233_), .B2(KEYINPUT29), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NOR3_X1   g058(.A1(new_n233_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n257_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n260_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(new_n258_), .A3(new_n256_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n253_), .B(KEYINPUT89), .Z(new_n265_));
  OAI211_X1 g064(.A(new_n255_), .B(new_n264_), .C1(new_n252_), .C2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n254_), .A2(KEYINPUT90), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n264_), .B1(new_n252_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT91), .ZN(new_n269_));
  OAI221_X1 g068(.A(new_n238_), .B1(KEYINPUT90), .B2(new_n254_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n266_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G8gat), .B(G36gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT18), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G64gat), .B(G92gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  NAND2_X1  g078(.A1(G226gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT93), .ZN(new_n281_));
  XOR2_X1   g080(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  AND3_X1   g083(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G183gat), .ZN(new_n288_));
  INV_X1    g087(.A(G190gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G169gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT22), .ZN(new_n293_));
  INV_X1    g092(.A(G176gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(G169gat), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n287_), .A2(new_n290_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n294_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(KEYINPUT24), .A3(new_n298_), .ZN(new_n299_));
  OR3_X1    g098(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n287_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n289_), .A2(KEYINPUT26), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT26), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G190gat), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT25), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G183gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n288_), .A2(KEYINPUT25), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT82), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n288_), .A2(KEYINPUT82), .A3(KEYINPUT25), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n305_), .A2(new_n307_), .A3(new_n310_), .A4(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n296_), .B1(new_n301_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n313_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n214_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n302_), .A2(new_n304_), .A3(new_n308_), .A4(new_n307_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n316_), .A2(new_n299_), .A3(new_n287_), .A4(new_n300_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT94), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n296_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n301_), .A2(KEYINPUT94), .A3(new_n316_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n315_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n314_), .B(KEYINPUT20), .C1(new_n321_), .C2(KEYINPUT95), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n320_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n214_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT95), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n284_), .B1(new_n322_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT96), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT96), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n329_), .B(new_n284_), .C1(new_n322_), .C2(new_n326_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n246_), .A2(new_n313_), .A3(new_n247_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n319_), .A2(new_n315_), .A3(new_n320_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n333_), .A2(KEYINPUT20), .A3(new_n283_), .A4(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n279_), .B1(new_n331_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n279_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n335_), .ZN(new_n338_));
  AOI211_X1 g137(.A(new_n337_), .B(new_n338_), .C1(new_n328_), .C2(new_n330_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n275_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n331_), .A2(new_n279_), .A3(new_n335_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n296_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n315_), .A2(new_n317_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT20), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n284_), .B1(new_n332_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT99), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  OAI211_X1 g146(.A(KEYINPUT99), .B(new_n284_), .C1(new_n332_), .C2(new_n344_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n324_), .A2(new_n325_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n321_), .A2(KEYINPUT95), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n349_), .A2(KEYINPUT20), .A3(new_n350_), .A4(new_n314_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n347_), .B(new_n348_), .C1(new_n351_), .C2(new_n284_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n337_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n341_), .A2(KEYINPUT27), .A3(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G85gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT0), .B(G57gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362_));
  XOR2_X1   g161(.A(G127gat), .B(G134gat), .Z(new_n363_));
  XOR2_X1   g162(.A(G113gat), .B(G120gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(new_n233_), .B2(KEYINPUT97), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n363_), .B(new_n364_), .Z(new_n367_));
  INV_X1    g166(.A(KEYINPUT97), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n218_), .A2(new_n219_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n362_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT98), .B(KEYINPUT4), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n367_), .A2(new_n233_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n361_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n366_), .A2(new_n370_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n377_), .A2(new_n361_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n359_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n378_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n375_), .A2(new_n380_), .A3(new_n358_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n273_), .A2(new_n340_), .A3(new_n354_), .A4(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT101), .ZN(new_n384_));
  INV_X1    g183(.A(new_n273_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT33), .ZN(new_n386_));
  AOI211_X1 g185(.A(new_n386_), .B(new_n358_), .C1(new_n375_), .C2(new_n380_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n377_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n358_), .B1(new_n388_), .B2(new_n360_), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n371_), .A2(new_n361_), .A3(new_n374_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT33), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n387_), .B1(new_n379_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n330_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n329_), .B1(new_n351_), .B2(new_n284_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n335_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n337_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n392_), .A2(new_n396_), .A3(new_n341_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n279_), .A2(KEYINPUT32), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n379_), .A2(new_n381_), .B1(new_n352_), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n383_), .A2(new_n384_), .B1(new_n385_), .B2(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n340_), .A2(new_n354_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n403_), .A2(KEYINPUT101), .A3(new_n273_), .A4(new_n382_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(KEYINPUT84), .B(G43gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(new_n313_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G227gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(G15gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(G71gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n409_), .B(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT31), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n415_), .B1(new_n365_), .B2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n416_), .B2(new_n365_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(G99gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n414_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n414_), .A2(new_n420_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n403_), .A2(new_n385_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n382_), .ZN(new_n425_));
  OAI22_X1  g224(.A1(new_n405_), .A2(new_n423_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G15gat), .B(G22gat), .ZN(new_n428_));
  INV_X1    g227(.A(G1gat), .ZN(new_n429_));
  INV_X1    g228(.A(G8gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT14), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G1gat), .B(G8gat), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n432_), .B(new_n433_), .Z(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G29gat), .B(G36gat), .Z(new_n436_));
  XOR2_X1   g235(.A(G43gat), .B(G50gat), .Z(new_n437_));
  XOR2_X1   g236(.A(new_n436_), .B(new_n437_), .Z(new_n438_));
  OR2_X1    g237(.A1(new_n435_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G229gat), .A2(G233gat), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n438_), .B(KEYINPUT15), .Z(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n435_), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n434_), .B(new_n438_), .Z(new_n444_));
  INV_X1    g243(.A(new_n440_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n441_), .A2(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G113gat), .B(G141gat), .Z(new_n447_));
  XNOR2_X1  g246(.A(G169gat), .B(G197gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n446_), .A2(new_n449_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n427_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G106gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(KEYINPUT10), .B(G99gat), .Z(new_n458_));
  AOI21_X1  g257(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT9), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT65), .B(G85gat), .ZN(new_n461_));
  INV_X1    g260(.A(G92gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n460_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n463_), .B(KEYINPUT66), .Z(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT67), .B1(G85gat), .B2(G92gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n466_));
  MUX2_X1   g265(.A(KEYINPUT67), .B(new_n465_), .S(new_n466_), .Z(new_n467_));
  OAI21_X1  g266(.A(new_n459_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT8), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G85gat), .B(G92gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT69), .ZN(new_n472_));
  NOR2_X1   g271(.A1(G99gat), .A2(G106gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n472_), .B1(new_n473_), .B2(KEYINPUT68), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT7), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT68), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n476_), .B1(new_n475_), .B2(KEYINPUT69), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n474_), .A2(new_n475_), .B1(new_n473_), .B2(new_n477_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n469_), .B(new_n471_), .C1(new_n478_), .C2(new_n456_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n454_), .ZN(new_n480_));
  AND2_X1   g279(.A1(KEYINPUT70), .A2(KEYINPUT6), .ZN(new_n481_));
  NOR2_X1   g280(.A1(KEYINPUT70), .A2(KEYINPUT6), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT70), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n455_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(KEYINPUT70), .A2(KEYINPUT6), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n454_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT71), .B1(new_n483_), .B2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n485_), .A2(new_n454_), .A3(new_n486_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT71), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n474_), .A2(new_n475_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n477_), .A2(new_n473_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n488_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n469_), .B1(new_n496_), .B2(new_n471_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n479_), .B1(new_n497_), .B2(KEYINPUT72), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT72), .ZN(new_n499_));
  AOI211_X1 g298(.A(new_n499_), .B(new_n469_), .C1(new_n496_), .C2(new_n471_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n468_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n442_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n468_), .B(new_n438_), .C1(new_n498_), .C2(new_n500_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G232gat), .A2(G233gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT34), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT35), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G190gat), .B(G218gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT74), .ZN(new_n511_));
  XOR2_X1   g310(.A(G134gat), .B(G162gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n514_), .A2(KEYINPUT36), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n503_), .A2(new_n504_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n506_), .A2(KEYINPUT35), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n508_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT75), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT75), .ZN(new_n520_));
  INV_X1    g319(.A(new_n518_), .ZN(new_n521_));
  AOI211_X1 g320(.A(new_n520_), .B(new_n521_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n509_), .B(new_n515_), .C1(new_n519_), .C2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT37), .ZN(new_n524_));
  INV_X1    g323(.A(new_n509_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n504_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n491_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n527_), .A2(new_n478_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n470_), .B1(new_n528_), .B2(new_n492_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n499_), .B1(new_n529_), .B2(new_n469_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n496_), .A2(new_n471_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(KEYINPUT72), .A3(KEYINPUT8), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n532_), .A3(new_n479_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n442_), .B1(new_n533_), .B2(new_n468_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n518_), .B1(new_n526_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n520_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n516_), .A2(KEYINPUT75), .A3(new_n518_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n525_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n513_), .B(KEYINPUT36), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n523_), .B(new_n524_), .C1(new_n538_), .C2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT77), .B1(new_n538_), .B2(new_n540_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT76), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n523_), .A2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n509_), .B1(new_n519_), .B2(new_n522_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT77), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n539_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n536_), .A2(new_n537_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n549_), .A2(KEYINPUT76), .A3(new_n509_), .A4(new_n515_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n543_), .A2(new_n545_), .A3(new_n548_), .A4(new_n550_), .ZN(new_n551_));
  AOI211_X1 g350(.A(KEYINPUT78), .B(new_n542_), .C1(KEYINPUT37), .C2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT78), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n543_), .A2(new_n548_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n545_), .A2(new_n550_), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT37), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n553_), .B1(new_n556_), .B2(new_n541_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G231gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n434_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G57gat), .B(G64gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT11), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G71gat), .B(G78gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n561_), .A2(KEYINPUT11), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n567_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n560_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G127gat), .B(G155gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT16), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G183gat), .B(G211gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(KEYINPUT79), .A2(KEYINPUT17), .ZN(new_n575_));
  OR3_X1    g374(.A1(new_n570_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  MUX2_X1   g375(.A(new_n575_), .B(KEYINPUT17), .S(new_n574_), .Z(new_n577_));
  NAND2_X1  g376(.A1(new_n570_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT80), .Z(new_n580_));
  NOR2_X1   g379(.A1(new_n558_), .A2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n568_), .B1(new_n533_), .B2(new_n468_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(KEYINPUT12), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT73), .Z(new_n584_));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT64), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n533_), .A2(new_n568_), .A3(new_n468_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(KEYINPUT12), .B2(new_n582_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n584_), .A2(new_n587_), .A3(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n586_), .B1(new_n589_), .B2(new_n582_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G120gat), .B(G148gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT5), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n597_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n591_), .A2(new_n592_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n598_), .A2(KEYINPUT13), .A3(new_n600_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n581_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n453_), .B1(new_n607_), .B2(KEYINPUT81), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(KEYINPUT81), .B2(new_n607_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n382_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n429_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT38), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT102), .B1(new_n605_), .B2(new_n452_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n523_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n427_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n579_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT102), .ZN(new_n619_));
  INV_X1    g418(.A(new_n452_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n603_), .A2(new_n619_), .A3(new_n604_), .A4(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n614_), .A2(new_n617_), .A3(new_n618_), .A4(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G1gat), .B1(new_n622_), .B2(new_n382_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n611_), .A2(new_n612_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n613_), .A2(new_n623_), .A3(new_n624_), .ZN(G1324gat));
  OAI21_X1  g424(.A(G8gat), .B1(new_n622_), .B2(new_n403_), .ZN(new_n626_));
  XOR2_X1   g425(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n403_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n609_), .A2(new_n430_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n626_), .A2(new_n628_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n629_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g433(.A(new_n423_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G15gat), .B1(new_n622_), .B2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT41), .Z(new_n637_));
  NAND3_X1  g436(.A1(new_n609_), .A2(new_n411_), .A3(new_n423_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1326gat));
  OAI21_X1  g438(.A(G22gat), .B1(new_n622_), .B2(new_n385_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT42), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n385_), .A2(G22gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT104), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n609_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(G1327gat));
  NAND2_X1  g444(.A1(new_n580_), .A2(new_n616_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n605_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n453_), .A2(new_n647_), .ZN(new_n648_));
  OR3_X1    g447(.A1(new_n648_), .A2(G29gat), .A3(new_n382_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n556_), .A2(new_n541_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT78), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n556_), .A2(new_n553_), .A3(new_n541_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n423_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n424_), .A2(new_n425_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n655_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n654_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n652_), .A2(KEYINPUT105), .A3(new_n653_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n661_), .B1(new_n552_), .B2(new_n557_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(new_n662_), .A3(new_n426_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n659_), .B1(new_n663_), .B2(KEYINPUT43), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n614_), .A2(new_n580_), .A3(new_n621_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n650_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(KEYINPUT43), .ZN(new_n668_));
  INV_X1    g467(.A(new_n659_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n665_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(KEYINPUT44), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT106), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(KEYINPUT44), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n667_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(new_n610_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n678_), .A2(KEYINPUT107), .ZN(new_n679_));
  OAI21_X1  g478(.A(G29gat), .B1(new_n678_), .B2(KEYINPUT107), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n649_), .B1(new_n679_), .B2(new_n680_), .ZN(G1328gat));
  NOR3_X1   g480(.A1(new_n648_), .A2(G36gat), .A3(new_n403_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT45), .Z(new_n683_));
  NAND2_X1  g482(.A1(new_n666_), .A2(new_n630_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686_));
  INV_X1    g485(.A(G36gat), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n685_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n675_), .B1(new_n674_), .B2(KEYINPUT44), .ZN(new_n689_));
  NOR4_X1   g488(.A1(new_n664_), .A2(KEYINPUT106), .A3(new_n665_), .A4(new_n650_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n630_), .B(new_n666_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT108), .B1(new_n691_), .B2(G36gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n683_), .B1(new_n688_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT109), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n694_), .A2(KEYINPUT109), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n693_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n686_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n691_), .A2(KEYINPUT108), .A3(G36gat), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n700_), .A2(KEYINPUT109), .A3(new_n694_), .A4(new_n683_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n697_), .A2(new_n701_), .ZN(G1329gat));
  NAND3_X1  g501(.A1(new_n677_), .A2(G43gat), .A3(new_n423_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n648_), .A2(new_n635_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(G43gat), .B2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(G1330gat));
  INV_X1    g506(.A(G50gat), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n385_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n453_), .A2(new_n273_), .A3(new_n647_), .ZN(new_n710_));
  AOI22_X1  g509(.A1(new_n677_), .A2(new_n709_), .B1(new_n708_), .B2(new_n710_), .ZN(G1331gat));
  INV_X1    g510(.A(new_n580_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n606_), .A2(new_n620_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n617_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G57gat), .B1(new_n714_), .B2(new_n382_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n426_), .A2(new_n452_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT111), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(new_n605_), .A3(new_n581_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n382_), .A2(G57gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n715_), .B1(new_n718_), .B2(new_n719_), .ZN(G1332gat));
  OAI21_X1  g519(.A(G64gat), .B1(new_n714_), .B2(new_n403_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT48), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n403_), .A2(G64gat), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT112), .Z(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(new_n718_), .B2(new_n724_), .ZN(G1333gat));
  OAI21_X1  g524(.A(G71gat), .B1(new_n714_), .B2(new_n635_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT49), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n635_), .A2(G71gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n718_), .B2(new_n728_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT113), .Z(G1334gat));
  OAI21_X1  g529(.A(G78gat), .B1(new_n714_), .B2(new_n385_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT50), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n385_), .A2(G78gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n718_), .B2(new_n733_), .ZN(G1335gat));
  NAND4_X1  g533(.A1(new_n717_), .A2(new_n605_), .A3(new_n616_), .A4(new_n580_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G85gat), .B1(new_n736_), .B2(new_n610_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n713_), .A2(new_n580_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n664_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n740_), .A2(new_n461_), .A3(new_n382_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n737_), .A2(new_n741_), .ZN(G1336gat));
  OAI21_X1  g541(.A(G92gat), .B1(new_n740_), .B2(new_n403_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n630_), .A2(new_n462_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n735_), .B2(new_n744_), .ZN(G1337gat));
  OAI21_X1  g544(.A(G99gat), .B1(new_n740_), .B2(new_n635_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n423_), .A2(new_n458_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n735_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g548(.A1(new_n736_), .A2(new_n457_), .A3(new_n273_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n739_), .B2(new_n273_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n754_));
  INV_X1    g553(.A(new_n738_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n670_), .A2(new_n751_), .A3(new_n273_), .A4(new_n755_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n753_), .A2(new_n754_), .A3(G106gat), .A4(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(G106gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT115), .B1(new_n759_), .B2(new_n752_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n757_), .A2(new_n758_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n758_), .B1(new_n757_), .B2(new_n760_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n750_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT53), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n750_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  NOR3_X1   g566(.A1(new_n424_), .A2(new_n382_), .A3(new_n635_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n607_), .A2(new_n620_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n443_), .A2(new_n439_), .A3(new_n445_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n449_), .B1(new_n444_), .B2(new_n440_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n450_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n600_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n584_), .A2(KEYINPUT55), .A3(new_n590_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n777_), .A2(KEYINPUT118), .A3(new_n587_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n778_), .A2(new_n599_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n591_), .A2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(new_n777_), .C1(KEYINPUT118), .C2(new_n587_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT56), .B1(new_n779_), .B2(new_n782_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n776_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT58), .B(new_n776_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n601_), .A2(new_n790_), .A3(new_n775_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n790_), .B1(new_n601_), .B2(new_n775_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n600_), .A2(new_n620_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n616_), .B1(new_n794_), .B2(new_n798_), .ZN(new_n799_));
  OAI22_X1  g598(.A1(new_n789_), .A2(new_n654_), .B1(new_n799_), .B2(KEYINPUT57), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n799_), .A2(KEYINPUT57), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n579_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n769_), .B1(new_n772_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(G113gat), .B1(new_n803_), .B2(new_n620_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n772_), .A2(new_n802_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n768_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT120), .B1(new_n806_), .B2(KEYINPUT59), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n803_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n801_), .B1(new_n800_), .B2(KEYINPUT121), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n813_));
  OAI221_X1 g612(.A(new_n813_), .B1(new_n799_), .B2(KEYINPUT57), .C1(new_n789_), .C2(new_n654_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n712_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n772_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n809_), .B(new_n768_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n811_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n620_), .A2(G113gat), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT122), .Z(new_n821_));
  AOI21_X1  g620(.A(new_n804_), .B1(new_n819_), .B2(new_n821_), .ZN(G1340gat));
  OAI211_X1 g621(.A(new_n605_), .B(new_n817_), .C1(new_n807_), .C2(new_n810_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(G120gat), .ZN(new_n824_));
  INV_X1    g623(.A(G120gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n606_), .B2(KEYINPUT60), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n803_), .B(new_n826_), .C1(KEYINPUT60), .C2(new_n825_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n824_), .A2(new_n827_), .ZN(G1341gat));
  OAI211_X1 g627(.A(new_n618_), .B(new_n817_), .C1(new_n807_), .C2(new_n810_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G127gat), .ZN(new_n830_));
  OR3_X1    g629(.A1(new_n806_), .A2(G127gat), .A3(new_n580_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1342gat));
  AOI21_X1  g631(.A(G134gat), .B1(new_n803_), .B2(new_n616_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT123), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n558_), .A2(G134gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n819_), .B2(new_n835_), .ZN(G1343gat));
  NOR4_X1   g635(.A1(new_n630_), .A2(new_n385_), .A3(new_n382_), .A4(new_n423_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n805_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n620_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n605_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT124), .B(G148gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1345gat));
  NAND3_X1  g642(.A1(new_n805_), .A2(new_n712_), .A3(new_n837_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n844_), .A2(KEYINPUT125), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(KEYINPUT125), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1346gat));
  AOI21_X1  g649(.A(G162gat), .B1(new_n838_), .B2(new_n616_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n660_), .A2(new_n662_), .A3(G162gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n838_), .B2(new_n852_), .ZN(G1347gat));
  NOR2_X1   g652(.A1(new_n403_), .A2(new_n425_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT126), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n385_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n620_), .B(new_n857_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT62), .B(new_n291_), .C1(new_n858_), .C2(KEYINPUT22), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(KEYINPUT62), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n291_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT62), .B1(new_n858_), .B2(KEYINPUT22), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n862_), .B2(new_n863_), .ZN(G1348gat));
  NOR2_X1   g663(.A1(new_n815_), .A2(new_n816_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n856_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G176gat), .B1(new_n866_), .B2(new_n605_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n856_), .B1(new_n772_), .B2(new_n802_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n606_), .A2(new_n294_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n868_), .B2(new_n869_), .ZN(G1349gat));
  AOI21_X1  g669(.A(G183gat), .B1(new_n868_), .B2(new_n712_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n579_), .B1(new_n308_), .B2(new_n307_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n866_), .B2(new_n872_), .ZN(G1350gat));
  NAND3_X1  g672(.A1(new_n866_), .A2(new_n616_), .A3(new_n305_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n865_), .A2(new_n654_), .A3(new_n856_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n289_), .B2(new_n875_), .ZN(G1351gat));
  NAND4_X1  g675(.A1(new_n630_), .A2(new_n273_), .A3(new_n382_), .A4(new_n635_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n772_), .B2(new_n802_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n620_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n605_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g681(.A(KEYINPUT63), .B(G211gat), .Z(new_n883_));
  NAND3_X1  g682(.A1(new_n878_), .A2(new_n618_), .A3(new_n883_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n884_), .A2(KEYINPUT127), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n884_), .A2(KEYINPUT127), .ZN(new_n886_));
  AOI211_X1 g685(.A(KEYINPUT63), .B(G211gat), .C1(new_n878_), .C2(new_n618_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n885_), .A2(new_n886_), .A3(new_n887_), .ZN(G1354gat));
  INV_X1    g687(.A(G218gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n878_), .A2(new_n889_), .A3(new_n616_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n878_), .A2(new_n558_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n889_), .ZN(G1355gat));
endmodule


