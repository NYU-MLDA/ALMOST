//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n959_, new_n960_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_;
  XNOR2_X1  g000(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT35), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT8), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT66), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n209_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(KEYINPUT66), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n215_));
  AOI22_X1  g014(.A1(new_n214_), .A2(new_n215_), .B1(G99gat), .B2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  INV_X1    g016(.A(G99gat), .ZN(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NOR3_X1   g021(.A1(new_n213_), .A2(new_n216_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G85gat), .ZN(new_n224_));
  INV_X1    g023(.A(G92gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n207_), .B1(new_n223_), .B2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G29gat), .B(G36gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G43gat), .B(G50gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n213_), .A2(new_n216_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT9), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n226_), .A2(new_n227_), .B1(new_n234_), .B2(G92gat), .ZN(new_n235_));
  AND2_X1   g034(.A1(G85gat), .A2(G92gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G85gat), .A2(G92gat), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n236_), .A2(new_n237_), .A3(KEYINPUT9), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT65), .B1(new_n235_), .B2(new_n238_), .ZN(new_n239_));
  OAI22_X1  g038(.A1(new_n236_), .A2(new_n237_), .B1(KEYINPUT9), .B2(new_n225_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n240_), .B(new_n241_), .C1(KEYINPUT9), .C2(new_n228_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT10), .B(G99gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT64), .B(G106gat), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n233_), .A2(new_n239_), .A3(new_n242_), .A4(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n222_), .A2(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n214_), .A2(new_n215_), .A3(G99gat), .A4(G106gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n220_), .A2(KEYINPUT67), .A3(new_n221_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n212_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .A4(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n228_), .A2(new_n207_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n229_), .A2(new_n232_), .A3(new_n246_), .A4(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n204_), .A2(new_n205_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(KEYINPUT73), .A3(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n229_), .A2(new_n254_), .A3(new_n246_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n232_), .B(KEYINPUT15), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT73), .B1(new_n255_), .B2(new_n256_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n206_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT74), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n265_), .B(new_n206_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n255_), .A2(new_n256_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n206_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n260_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n264_), .A2(new_n266_), .A3(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G190gat), .B(G218gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT75), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G134gat), .B(G162gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT36), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n274_), .A2(new_n275_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n270_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n269_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n263_), .B2(KEYINPUT74), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n280_), .A2(new_n275_), .A3(new_n274_), .A4(new_n266_), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n278_), .A2(KEYINPUT37), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT37), .B1(new_n278_), .B2(new_n281_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G127gat), .B(G155gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(G183gat), .B(G211gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT17), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT77), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G15gat), .B(G22gat), .ZN(new_n293_));
  INV_X1    g092(.A(G1gat), .ZN(new_n294_));
  INV_X1    g093(.A(G8gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT14), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n298_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G231gat), .A2(G233gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  XNOR2_X1  g102(.A(G57gat), .B(G64gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT11), .ZN(new_n305_));
  XOR2_X1   g104(.A(G71gat), .B(G78gat), .Z(new_n306_));
  OR2_X1    g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n304_), .A2(KEYINPUT11), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n306_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n307_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n303_), .B(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n292_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n310_), .B(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n303_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n303_), .A2(new_n314_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n289_), .A2(new_n290_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n291_), .A4(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n312_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n284_), .A2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n321_), .B(KEYINPUT78), .Z(new_n322_));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G197gat), .B(G204gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT21), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G211gat), .B(G218gat), .Z(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(G197gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT21), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT91), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n331_), .B1(new_n332_), .B2(new_n324_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G211gat), .B(G218gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(G204gat), .ZN(new_n335_));
  INV_X1    g134(.A(G204gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G197gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n334_), .B1(new_n338_), .B2(KEYINPUT21), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n328_), .B1(new_n333_), .B2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT22), .B(G169gat), .ZN(new_n341_));
  INV_X1    g140(.A(G176gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n346_), .B(new_n347_), .C1(G183gat), .C2(G190gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n343_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n340_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT97), .ZN(new_n353_));
  INV_X1    g152(.A(G183gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT25), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G183gat), .ZN(new_n357_));
  INV_X1    g156(.A(G190gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT26), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT26), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(G190gat), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n355_), .A2(new_n357_), .A3(new_n359_), .A4(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G169gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n342_), .ZN(new_n364_));
  AND2_X1   g163(.A1(KEYINPUT95), .A2(KEYINPUT24), .ZN(new_n365_));
  NOR2_X1   g164(.A1(KEYINPUT95), .A2(KEYINPUT24), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n364_), .B(new_n349_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT96), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT96), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n362_), .A2(new_n367_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n344_), .B(new_n345_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n353_), .B1(new_n372_), .B2(new_n375_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n362_), .A2(new_n367_), .A3(new_n370_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n370_), .B1(new_n362_), .B2(new_n367_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n353_), .B(new_n375_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n352_), .B1(new_n376_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT98), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n327_), .B1(new_n325_), .B2(new_n324_), .ZN(new_n383_));
  OAI211_X1 g182(.A(KEYINPUT21), .B(new_n330_), .C1(new_n338_), .C2(KEYINPUT91), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n383_), .A2(new_n384_), .B1(new_n327_), .B2(new_n326_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n350_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n375_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT97), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n386_), .B1(new_n388_), .B2(new_n379_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT98), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT20), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT94), .ZN(new_n394_));
  XOR2_X1   g193(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT26), .B(G190gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n355_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT25), .B(G183gat), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n397_), .B(new_n399_), .C1(new_n400_), .C2(new_n398_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n344_), .B(KEYINPUT23), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n364_), .A2(KEYINPUT24), .A3(new_n349_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n364_), .A2(KEYINPUT24), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .A4(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n363_), .A2(KEYINPUT84), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT22), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT22), .B1(new_n407_), .B2(G169gat), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n409_), .B(new_n342_), .C1(new_n410_), .C2(new_n406_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(new_n349_), .A3(new_n348_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n405_), .A2(new_n412_), .ZN(new_n413_));
  AOI211_X1 g212(.A(new_n392_), .B(new_n396_), .C1(new_n413_), .C2(new_n340_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n382_), .A2(new_n391_), .A3(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT20), .B1(new_n413_), .B2(new_n340_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n351_), .B1(new_n388_), .B2(new_n379_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(new_n385_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n396_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT18), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G64gat), .B(G92gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n415_), .A2(new_n420_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n425_), .B1(new_n415_), .B2(new_n420_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n323_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n415_), .A2(new_n420_), .A3(new_n425_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n396_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n417_), .B(new_n430_), .C1(new_n418_), .C2(new_n385_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n352_), .A2(new_n387_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n405_), .A2(new_n412_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT20), .B1(new_n433_), .B2(new_n385_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n396_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n424_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n429_), .A2(new_n437_), .A3(KEYINPUT27), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n428_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT85), .B(G43gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT31), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n433_), .A2(KEYINPUT30), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT30), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n413_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(G15gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(G71gat), .ZN(new_n449_));
  INV_X1    g248(.A(G15gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n447_), .B(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(G71gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n449_), .A2(new_n453_), .A3(G99gat), .ZN(new_n454_));
  AOI21_X1  g253(.A(G99gat), .B1(new_n449_), .B2(new_n453_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n446_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G127gat), .B(G134gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G113gat), .B(G120gat), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n459_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n443_), .B(new_n445_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n457_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n462_), .B1(new_n457_), .B2(new_n463_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n442_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(new_n441_), .A3(new_n464_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G141gat), .ZN(new_n472_));
  INV_X1    g271(.A(G148gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G141gat), .A2(G148gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n477_));
  INV_X1    g276(.A(G155gat), .ZN(new_n478_));
  INV_X1    g277(.A(G162gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G155gat), .A2(G162gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT1), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n476_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n472_), .A2(new_n473_), .A3(KEYINPUT3), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT3), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(G141gat), .B2(G148gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT88), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT2), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n491_), .A2(new_n492_), .B1(new_n475_), .B2(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(KEYINPUT88), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n490_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n480_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n496_), .A2(KEYINPUT89), .A3(new_n497_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n486_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT29), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n486_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n496_), .A2(KEYINPUT89), .A3(new_n497_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT89), .B1(new_n496_), .B2(new_n497_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n503_), .B(new_n506_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n504_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n505_), .A2(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G22gat), .B(G50gat), .Z(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n505_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G78gat), .B(G106gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n340_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n520_));
  INV_X1    g319(.A(G228gat), .ZN(new_n521_));
  INV_X1    g320(.A(G233gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  OAI221_X1 g323(.A(new_n340_), .B1(new_n521_), .B2(new_n522_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n519_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT92), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n517_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n525_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n518_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n525_), .A3(new_n519_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n530_), .A2(new_n517_), .A3(new_n527_), .A4(new_n531_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G225gat), .A2(G233gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n462_), .A2(KEYINPUT99), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT99), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n460_), .A2(new_n538_), .A3(new_n461_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n502_), .B2(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n506_), .B(new_n539_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n537_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n536_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G1gat), .B(G29gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(G85gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT0), .B(G57gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT4), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n541_), .A2(new_n542_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n500_), .A2(new_n501_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n552_), .A2(new_n506_), .A3(new_n537_), .A4(new_n539_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n550_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n506_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n462_), .A2(KEYINPUT4), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n536_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n544_), .B(new_n549_), .C1(new_n554_), .C2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n558_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT4), .B1(new_n540_), .B2(new_n543_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n536_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n560_), .B1(new_n564_), .B2(new_n549_), .ZN(new_n565_));
  NOR4_X1   g364(.A1(new_n439_), .A2(new_n471_), .A3(new_n535_), .A4(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n425_), .A2(KEYINPUT32), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n415_), .A2(new_n420_), .A3(KEYINPUT103), .A4(new_n567_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n415_), .A2(new_n420_), .A3(new_n567_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT103), .ZN(new_n570_));
  INV_X1    g369(.A(new_n567_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n570_), .B1(new_n436_), .B2(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n565_), .B(new_n568_), .C1(new_n569_), .C2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n350_), .B1(new_n376_), .B2(new_n380_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n416_), .B1(new_n574_), .B2(new_n340_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n414_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n576_));
  AOI211_X1 g375(.A(KEYINPUT98), .B(new_n386_), .C1(new_n388_), .C2(new_n379_), .ZN(new_n577_));
  OAI22_X1  g376(.A1(new_n575_), .A2(new_n430_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n424_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT101), .B(KEYINPUT33), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n560_), .A2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n558_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n549_), .B1(new_n562_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT102), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n584_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n551_), .A2(new_n553_), .A3(KEYINPUT102), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n558_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n579_), .A2(new_n581_), .A3(new_n429_), .A4(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT100), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n590_), .B1(new_n560_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n562_), .A2(new_n563_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n561_), .A2(new_n548_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n593_), .A2(new_n594_), .A3(KEYINPUT100), .A4(KEYINPUT33), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n573_), .B1(new_n589_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n535_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n579_), .A2(new_n429_), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT20), .B(new_n430_), .C1(new_n433_), .C2(new_n385_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n381_), .B2(KEYINPUT98), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n602_), .A2(new_n391_), .B1(new_n419_), .B2(new_n396_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n323_), .B1(new_n603_), .B2(new_n425_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n600_), .A2(new_n323_), .B1(new_n604_), .B2(new_n437_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n565_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n599_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n470_), .B(KEYINPUT86), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n566_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611_));
  INV_X1    g410(.A(new_n258_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n611_), .B1(new_n314_), .B2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n310_), .B(KEYINPUT68), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n258_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(KEYINPUT12), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT12), .ZN(new_n617_));
  INV_X1    g416(.A(new_n310_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n258_), .B2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n613_), .B1(new_n616_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT69), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n614_), .B2(new_n258_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n314_), .A2(KEYINPUT69), .A3(new_n612_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n615_), .A3(new_n623_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n624_), .A2(KEYINPUT70), .A3(new_n611_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT70), .B1(new_n624_), .B2(new_n611_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n620_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT5), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n629_), .B(new_n630_), .Z(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n631_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n620_), .B(new_n633_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT13), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n632_), .B(new_n634_), .C1(KEYINPUT71), .C2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n259_), .A2(new_n301_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT80), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n259_), .A2(KEYINPUT80), .A3(new_n301_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G229gat), .A2(G233gat), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT79), .ZN(new_n647_));
  INV_X1    g446(.A(new_n301_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n648_), .B2(new_n232_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n647_), .A3(new_n232_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n645_), .B(new_n646_), .C1(new_n649_), .C2(new_n651_), .ZN(new_n652_));
  OAI22_X1  g451(.A1(new_n651_), .A2(new_n649_), .B1(new_n648_), .B2(new_n232_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n646_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(G113gat), .B(G141gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT81), .ZN(new_n658_));
  XNOR2_X1  g457(.A(G169gat), .B(G197gat), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n658_), .B(new_n659_), .Z(new_n660_));
  NAND2_X1  g459(.A1(new_n656_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n660_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n652_), .A2(new_n655_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n640_), .A2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n610_), .A2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n322_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n294_), .A3(new_n565_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT38), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n278_), .A2(new_n281_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n610_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n665_), .A2(new_n319_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n565_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G1gat), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n668_), .A2(new_n669_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n670_), .A2(new_n677_), .A3(new_n678_), .ZN(G1324gat));
  NAND3_X1  g478(.A1(new_n673_), .A2(new_n674_), .A3(new_n439_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n680_), .A2(new_n681_), .A3(G8gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n680_), .B2(G8gat), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n686_), .A3(KEYINPUT39), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n686_), .A2(KEYINPUT39), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n667_), .A2(new_n295_), .A3(new_n439_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n687_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n687_), .A2(new_n688_), .A3(KEYINPUT40), .A4(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1325gat));
  OAI21_X1  g493(.A(G15gat), .B1(new_n675_), .B2(new_n609_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT41), .Z(new_n696_));
  XOR2_X1   g495(.A(new_n470_), .B(KEYINPUT86), .Z(new_n697_));
  NAND3_X1  g496(.A1(new_n667_), .A2(new_n450_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1326gat));
  OAI21_X1  g498(.A(G22gat), .B1(new_n675_), .B2(new_n598_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT42), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n598_), .A2(G22gat), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT106), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n667_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(G1327gat));
  NOR2_X1   g504(.A1(new_n671_), .A2(new_n320_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n666_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G29gat), .B1(new_n708_), .B2(new_n565_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n640_), .A2(new_n664_), .A3(new_n319_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n610_), .B2(new_n284_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n439_), .A2(new_n535_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(new_n676_), .A3(new_n470_), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n597_), .A2(new_n598_), .B1(new_n606_), .B2(new_n605_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(new_n697_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n716_));
  INV_X1    g515(.A(new_n284_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n710_), .B1(new_n711_), .B2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n720_));
  INV_X1    g519(.A(new_n710_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n426_), .A2(new_n427_), .ZN(new_n722_));
  AOI22_X1  g521(.A1(new_n560_), .A2(new_n580_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n722_), .A2(new_n723_), .A3(new_n592_), .A4(new_n595_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n535_), .B1(new_n724_), .B2(new_n573_), .ZN(new_n725_));
  AND4_X1   g524(.A1(new_n535_), .A2(new_n676_), .A3(new_n428_), .A4(new_n438_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n609_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  AOI211_X1 g526(.A(KEYINPUT43), .B(new_n284_), .C1(new_n727_), .C2(new_n713_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n716_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT44), .B(new_n721_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n721_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n734_));
  AOI22_X1  g533(.A1(new_n720_), .A2(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n565_), .A2(G29gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n709_), .B1(new_n735_), .B2(new_n736_), .ZN(G1328gat));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739_));
  INV_X1    g538(.A(G36gat), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n666_), .A2(new_n740_), .A3(new_n439_), .A4(new_n706_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n605_), .B1(new_n734_), .B2(new_n733_), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT107), .B1(new_n719_), .B2(KEYINPUT44), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n730_), .A2(new_n731_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n744_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n743_), .B1(new_n747_), .B2(G36gat), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n738_), .B(new_n739_), .C1(new_n748_), .C2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n743_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n439_), .B1(new_n719_), .B2(KEYINPUT44), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n732_), .B2(new_n720_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n751_), .B1(new_n753_), .B2(new_n740_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT109), .B1(new_n754_), .B2(KEYINPUT108), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT46), .B1(new_n748_), .B2(new_n738_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n750_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(G1329gat));
  AOI21_X1  g557(.A(G43gat), .B1(new_n708_), .B2(new_n697_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n470_), .A2(G43gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n735_), .B2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(G1330gat));
  OR3_X1    g562(.A1(new_n707_), .A2(G50gat), .A3(new_n598_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n735_), .A2(new_n535_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n765_), .A2(KEYINPUT111), .ZN(new_n766_));
  OAI21_X1  g565(.A(G50gat), .B1(new_n765_), .B2(KEYINPUT111), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n764_), .B1(new_n766_), .B2(new_n767_), .ZN(G1331gat));
  INV_X1    g567(.A(new_n640_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n664_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n610_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n322_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(G57gat), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n565_), .ZN(new_n776_));
  NOR4_X1   g575(.A1(new_n771_), .A2(new_n610_), .A3(new_n319_), .A4(new_n672_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(new_n565_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n776_), .B1(new_n775_), .B2(new_n778_), .ZN(G1332gat));
  INV_X1    g578(.A(G64gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n777_), .B2(new_n439_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT48), .Z(new_n782_));
  NAND3_X1  g581(.A1(new_n774_), .A2(new_n780_), .A3(new_n439_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1333gat));
  AOI21_X1  g583(.A(new_n452_), .B1(new_n777_), .B2(new_n697_), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT49), .Z(new_n786_));
  NAND3_X1  g585(.A1(new_n774_), .A2(new_n452_), .A3(new_n697_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(G1334gat));
  INV_X1    g587(.A(G78gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n777_), .B2(new_n535_), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT50), .Z(new_n791_));
  NAND3_X1  g590(.A1(new_n774_), .A2(new_n789_), .A3(new_n535_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT112), .ZN(G1335gat));
  NAND2_X1  g593(.A1(new_n711_), .A2(new_n718_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n771_), .A2(new_n320_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n795_), .A2(KEYINPUT113), .A3(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(G85gat), .B1(new_n802_), .B2(new_n676_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n772_), .A2(new_n706_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n224_), .A3(new_n565_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(G1336gat));
  OAI21_X1  g606(.A(G92gat), .B1(new_n802_), .B2(new_n605_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(new_n225_), .A3(new_n439_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1337gat));
  OR2_X1    g609(.A1(new_n471_), .A2(new_n243_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n812_));
  OAI22_X1  g611(.A1(new_n804_), .A2(new_n811_), .B1(KEYINPUT115), .B2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n218_), .B1(new_n801_), .B2(new_n697_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(KEYINPUT114), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(KEYINPUT115), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n609_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n218_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n815_), .A2(new_n816_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n816_), .B1(new_n815_), .B2(new_n819_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1338gat));
  OR3_X1    g621(.A1(new_n804_), .A2(new_n598_), .A3(new_n244_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n795_), .A2(new_n535_), .A3(new_n796_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(G106gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n824_), .B2(G106gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n823_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n616_), .A2(new_n619_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n622_), .A2(new_n623_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n611_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n620_), .A2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n613_), .B(KEYINPUT55), .C1(new_n616_), .C2(new_n619_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(KEYINPUT56), .A3(new_n631_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT56), .B1(new_n837_), .B2(new_n631_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n662_), .B1(new_n653_), .B2(new_n646_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n643_), .A2(new_n644_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n654_), .B1(new_n651_), .B2(new_n649_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n663_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n663_), .A2(new_n845_), .A3(KEYINPUT116), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n634_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n830_), .B1(new_n841_), .B2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n837_), .A2(new_n631_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n838_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n856_), .A2(KEYINPUT58), .A3(new_n634_), .A4(new_n850_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n852_), .A2(new_n857_), .A3(new_n717_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n664_), .A2(new_n634_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n855_), .B2(new_n838_), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT117), .B1(new_n635_), .B2(new_n850_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n635_), .A2(KEYINPUT117), .A3(new_n850_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n671_), .A2(KEYINPUT57), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n858_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n863_), .ZN(new_n867_));
  OAI22_X1  g666(.A1(new_n867_), .A2(new_n861_), .B1(new_n841_), .B2(new_n859_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n868_), .B2(new_n671_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n319_), .B1(new_n866_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n321_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n871_), .A2(new_n872_), .A3(new_n770_), .A4(new_n640_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n640_), .A2(new_n770_), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT54), .B1(new_n874_), .B2(new_n321_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n870_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n471_), .A2(new_n676_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n712_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n877_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(G113gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n882_), .A2(new_n883_), .A3(new_n664_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n879_), .A2(KEYINPUT59), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n876_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n870_), .B2(KEYINPUT118), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n889_), .B(new_n319_), .C1(new_n866_), .C2(new_n869_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n886_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n877_), .B2(new_n880_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n891_), .A2(new_n893_), .A3(new_n770_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n884_), .B1(new_n894_), .B2(new_n883_), .ZN(G1340gat));
  INV_X1    g694(.A(G120gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n640_), .B2(KEYINPUT60), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n882_), .B(new_n897_), .C1(KEYINPUT60), .C2(new_n896_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n891_), .A2(new_n893_), .A3(new_n640_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900_));
  OAI21_X1  g699(.A(G120gat), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  NOR4_X1   g700(.A1(new_n891_), .A2(new_n893_), .A3(KEYINPUT119), .A4(new_n640_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n898_), .B1(new_n901_), .B2(new_n902_), .ZN(G1341gat));
  NAND2_X1  g702(.A1(new_n888_), .A2(new_n890_), .ZN(new_n904_));
  AOI22_X1  g703(.A1(new_n904_), .A2(new_n885_), .B1(new_n881_), .B2(KEYINPUT59), .ZN(new_n905_));
  INV_X1    g704(.A(G127gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n319_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909_));
  OAI211_X1 g708(.A(KEYINPUT120), .B(new_n906_), .C1(new_n881_), .C2(new_n319_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n319_), .B(new_n879_), .C1(new_n870_), .C2(new_n876_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(G127gat), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n908_), .A2(new_n909_), .A3(new_n910_), .A4(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n910_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n907_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n891_), .A2(new_n893_), .A3(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(KEYINPUT121), .B1(new_n915_), .B2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n914_), .A2(new_n918_), .ZN(G1342gat));
  AOI21_X1  g718(.A(G134gat), .B1(new_n882_), .B2(new_n672_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n717_), .A2(G134gat), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(KEYINPUT122), .Z(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n905_), .B2(new_n922_), .ZN(G1343gat));
  NOR3_X1   g722(.A1(new_n697_), .A2(new_n598_), .A3(new_n676_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n877_), .A2(new_n605_), .A3(new_n924_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n770_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(new_n472_), .ZN(G1344gat));
  NOR2_X1   g726(.A1(new_n925_), .A2(new_n640_), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT123), .B(G148gat), .Z(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1345gat));
  NOR2_X1   g729(.A1(new_n925_), .A2(new_n319_), .ZN(new_n931_));
  XOR2_X1   g730(.A(KEYINPUT61), .B(G155gat), .Z(new_n932_));
  XNOR2_X1  g731(.A(new_n931_), .B(new_n932_), .ZN(G1346gat));
  OAI21_X1  g732(.A(G162gat), .B1(new_n925_), .B2(new_n284_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n672_), .A2(new_n479_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n925_), .B2(new_n935_), .ZN(G1347gat));
  NOR4_X1   g735(.A1(new_n609_), .A2(new_n535_), .A3(new_n565_), .A4(new_n605_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n904_), .A2(new_n937_), .ZN(new_n938_));
  OAI21_X1  g737(.A(G169gat), .B1(new_n938_), .B2(new_n770_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n938_), .A2(new_n942_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n904_), .A2(KEYINPUT125), .A3(new_n937_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n943_), .A2(new_n341_), .A3(new_n664_), .A4(new_n944_), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(KEYINPUT62), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n941_), .B(new_n945_), .C1(new_n939_), .C2(new_n947_), .ZN(G1348gat));
  NAND3_X1  g747(.A1(new_n943_), .A2(new_n769_), .A3(new_n944_), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n877_), .A2(new_n937_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n640_), .A2(new_n342_), .ZN(new_n951_));
  AOI22_X1  g750(.A1(new_n949_), .A2(new_n342_), .B1(new_n950_), .B2(new_n951_), .ZN(G1349gat));
  AOI21_X1  g751(.A(G183gat), .B1(new_n950_), .B2(new_n320_), .ZN(new_n953_));
  AND3_X1   g752(.A1(new_n904_), .A2(KEYINPUT125), .A3(new_n937_), .ZN(new_n954_));
  AOI21_X1  g753(.A(KEYINPUT125), .B1(new_n904_), .B2(new_n937_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n319_), .A2(new_n400_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n953_), .B1(new_n956_), .B2(new_n957_), .ZN(G1350gat));
  NAND4_X1  g757(.A1(new_n943_), .A2(new_n397_), .A3(new_n672_), .A4(new_n944_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n954_), .A2(new_n955_), .A3(new_n284_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n960_), .B2(new_n358_), .ZN(G1351gat));
  AND3_X1   g760(.A1(new_n609_), .A2(new_n606_), .A3(new_n439_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n877_), .A2(new_n962_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n963_), .A2(new_n770_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n964_), .B(new_n329_), .ZN(G1352gat));
  NOR2_X1   g764(.A1(new_n963_), .A2(new_n640_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(new_n336_), .ZN(G1353gat));
  INV_X1    g766(.A(new_n963_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n319_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n969_));
  XOR2_X1   g768(.A(new_n969_), .B(KEYINPUT126), .Z(new_n970_));
  NAND2_X1  g769(.A1(new_n968_), .A2(new_n970_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n971_), .B1(KEYINPUT127), .B2(new_n972_), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n972_), .B(KEYINPUT127), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n973_), .B1(new_n971_), .B2(new_n974_), .ZN(G1354gat));
  OR3_X1    g774(.A1(new_n963_), .A2(G218gat), .A3(new_n671_), .ZN(new_n976_));
  OAI21_X1  g775(.A(G218gat), .B1(new_n963_), .B2(new_n284_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n976_), .A2(new_n977_), .ZN(G1355gat));
endmodule


