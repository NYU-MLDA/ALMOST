//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n844_, new_n845_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G134gat), .ZN(new_n203_));
  INV_X1    g002(.A(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT36), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT35), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT15), .ZN(new_n208_));
  INV_X1    g007(.A(G50gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G29gat), .A2(G36gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n211_), .A2(new_n212_), .A3(G43gat), .ZN(new_n213_));
  INV_X1    g012(.A(G43gat), .ZN(new_n214_));
  INV_X1    g013(.A(G29gat), .ZN(new_n215_));
  INV_X1    g014(.A(G36gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n214_), .B1(new_n217_), .B2(new_n210_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n209_), .B1(new_n213_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n220_));
  OAI21_X1  g019(.A(G43gat), .B1(new_n211_), .B2(new_n212_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n217_), .A2(new_n214_), .A3(new_n210_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(G50gat), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n219_), .A2(new_n220_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n220_), .B1(new_n219_), .B2(new_n223_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n208_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n223_), .ZN(new_n227_));
  AOI21_X1  g026(.A(G50gat), .B1(new_n221_), .B2(new_n222_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT68), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n219_), .A2(new_n220_), .A3(new_n223_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(KEYINPUT15), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G85gat), .B(G92gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT9), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(KEYINPUT10), .B(G99gat), .Z(new_n235_));
  INV_X1    g034(.A(G106gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G99gat), .A2(G106gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT6), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT6), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(G99gat), .A3(G106gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n233_), .A2(G85gat), .A3(G92gat), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n234_), .A2(new_n237_), .A3(new_n242_), .A4(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(G99gat), .A2(G106gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT7), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n245_), .B1(KEYINPUT64), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT64), .B(KEYINPUT7), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n242_), .B(new_n247_), .C1(new_n245_), .C2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT8), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n232_), .A2(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n249_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n250_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n244_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n226_), .A2(new_n231_), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n207_), .B1(new_n256_), .B2(KEYINPUT69), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n253_), .A2(new_n254_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n227_), .A2(new_n228_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n244_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G232gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT34), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n257_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n263_), .A2(KEYINPUT35), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n256_), .A2(new_n260_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n266_), .B1(new_n257_), .B2(new_n263_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n206_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n256_), .A2(KEYINPUT69), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(KEYINPUT35), .A3(new_n263_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n266_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n273_));
  NAND3_X1  g072(.A1(new_n257_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .A4(new_n205_), .ZN(new_n275_));
  XOR2_X1   g074(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n276_));
  NAND3_X1  g075(.A1(new_n268_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT74), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n268_), .A2(KEYINPUT71), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n280_), .B(new_n206_), .C1(new_n264_), .C2(new_n267_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n275_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT37), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(KEYINPUT72), .A3(KEYINPUT37), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n278_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G57gat), .B(G64gat), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n288_), .A2(KEYINPUT11), .ZN(new_n289_));
  XOR2_X1   g088(.A(G71gat), .B(G78gat), .Z(new_n290_));
  OR2_X1    g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n288_), .A2(KEYINPUT11), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n290_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n255_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT66), .B(KEYINPUT12), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT66), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n255_), .B(new_n294_), .C1(new_n298_), .C2(KEYINPUT12), .ZN(new_n299_));
  INV_X1    g098(.A(new_n294_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n258_), .A2(new_n244_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G230gat), .A2(G233gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  OR3_X1    g103(.A1(new_n297_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n301_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n304_), .B1(new_n306_), .B2(new_n295_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G120gat), .B(G148gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G176gat), .B(G204gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n305_), .A2(new_n307_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n313_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n317_), .A2(KEYINPUT13), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(KEYINPUT13), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G231gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n294_), .B(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(KEYINPUT75), .B(KEYINPUT76), .Z(new_n323_));
  XNOR2_X1  g122(.A(G1gat), .B(G8gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G15gat), .ZN(new_n326_));
  INV_X1    g125(.A(G22gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G15gat), .A2(G22gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G1gat), .A2(G8gat), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n328_), .A2(new_n329_), .B1(KEYINPUT14), .B2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n325_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n322_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G127gat), .B(G155gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G183gat), .B(G211gat), .Z(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n338_), .A2(KEYINPUT17), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n340_), .A3(KEYINPUT17), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n333_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n333_), .A2(new_n341_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n287_), .A2(new_n320_), .A3(new_n346_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n347_), .A2(KEYINPUT79), .ZN(new_n348_));
  INV_X1    g147(.A(G204gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G197gat), .ZN(new_n350_));
  INV_X1    g149(.A(G197gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G204gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT21), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT21), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(new_n352_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G211gat), .ZN(new_n357_));
  INV_X1    g156(.A(G218gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G211gat), .A2(G218gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n354_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n360_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G211gat), .A2(G218gat), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT87), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT87), .B1(new_n359_), .B2(new_n360_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT21), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n353_), .A2(KEYINPUT88), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT88), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n350_), .A2(new_n352_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n362_), .B1(new_n368_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT2), .ZN(new_n374_));
  INV_X1    g173(.A(G141gat), .ZN(new_n375_));
  INV_X1    g174(.A(G148gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n374_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n377_), .A2(new_n379_), .A3(new_n380_), .A4(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT85), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(G155gat), .A3(G162gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n382_), .A2(new_n383_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT1), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n385_), .A2(new_n387_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT86), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(KEYINPUT1), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT86), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n385_), .A2(new_n387_), .A3(new_n394_), .A4(new_n390_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n392_), .A2(new_n393_), .A3(new_n383_), .A4(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G141gat), .B(G148gat), .Z(new_n397_));
  AOI21_X1  g196(.A(new_n389_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n373_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G78gat), .B(G106gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G228gat), .A2(G233gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n401_), .B(new_n402_), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n373_), .B(new_n403_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT89), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT89), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(new_n409_), .A3(new_n406_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n396_), .A2(new_n397_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n389_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(G50gat), .B1(new_n413_), .B2(KEYINPUT29), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n398_), .A2(new_n399_), .A3(new_n209_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT28), .B(G22gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n417_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n414_), .A2(new_n419_), .A3(new_n415_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n408_), .A2(new_n410_), .A3(new_n418_), .A4(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n420_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n410_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G183gat), .A2(G190gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT23), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n431_));
  INV_X1    g230(.A(G169gat), .ZN(new_n432_));
  INV_X1    g231(.A(G176gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n430_), .B(new_n431_), .C1(new_n434_), .C2(KEYINPUT24), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G169gat), .A2(G176gat), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n436_), .A2(KEYINPUT92), .A3(KEYINPUT24), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT92), .B1(new_n436_), .B2(KEYINPUT24), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n435_), .B1(new_n439_), .B2(new_n434_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT25), .B(G183gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT91), .ZN(new_n442_));
  NOR2_X1   g241(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n442_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n445_), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n447_), .A2(new_n443_), .A3(KEYINPUT91), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n441_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G183gat), .ZN(new_n453_));
  INV_X1    g252(.A(G190gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n433_), .A2(KEYINPUT82), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT82), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(G176gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT22), .B(G169gat), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n452_), .A2(new_n455_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n436_), .B(KEYINPUT93), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n440_), .A2(new_n449_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n361_), .A2(new_n365_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n359_), .A2(KEYINPUT87), .A3(new_n360_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n355_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n371_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n370_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n350_), .A2(new_n352_), .A3(new_n355_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n355_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n466_), .A2(new_n469_), .B1(new_n472_), .B2(new_n361_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n427_), .B1(new_n463_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G226gat), .A2(G233gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n475_), .B(KEYINPUT90), .Z(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT19), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT25), .B1(new_n453_), .B2(KEYINPUT81), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT81), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT25), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(G183gat), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n478_), .B(new_n481_), .C1(new_n443_), .C2(new_n447_), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n434_), .A2(KEYINPUT24), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n434_), .A2(KEYINPUT24), .A3(new_n436_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n482_), .A2(new_n452_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n459_), .A2(new_n460_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n430_), .A2(new_n455_), .A3(new_n431_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n436_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT94), .B1(new_n373_), .B2(new_n489_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n373_), .A2(KEYINPUT94), .A3(new_n489_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n474_), .B(new_n477_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT95), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n473_), .A2(new_n488_), .A3(new_n485_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n494_), .B(KEYINPUT20), .C1(new_n473_), .C2(new_n463_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n477_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n373_), .A2(new_n489_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT94), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n373_), .A2(new_n489_), .A3(KEYINPUT94), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT95), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n477_), .A4(new_n474_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n493_), .A2(new_n497_), .A3(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G8gat), .B(G36gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT18), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(G64gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(G92gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n493_), .A2(new_n511_), .A3(new_n504_), .A4(new_n497_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n495_), .A2(new_n496_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n477_), .B1(new_n502_), .B2(new_n474_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n509_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n512_), .A2(new_n518_), .A3(KEYINPUT27), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(G127gat), .ZN(new_n522_));
  INV_X1    g321(.A(G134gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G127gat), .A2(G134gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(G113gat), .ZN(new_n527_));
  INV_X1    g326(.A(G113gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n524_), .A2(new_n528_), .A3(new_n525_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(G120gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n413_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n530_), .B(G120gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n398_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(KEYINPUT4), .A3(new_n535_), .ZN(new_n536_));
  OR3_X1    g335(.A1(new_n398_), .A2(new_n534_), .A3(KEYINPUT4), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G225gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT96), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n536_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n533_), .A2(new_n541_), .A3(new_n535_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G1gat), .B(G29gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(G85gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT0), .ZN(new_n546_));
  INV_X1    g345(.A(G57gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n543_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT97), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n540_), .A2(new_n548_), .A3(new_n542_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n543_), .A2(KEYINPUT97), .A3(new_n549_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n426_), .B1(new_n521_), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G71gat), .B(G99gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT30), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G227gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(G15gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n558_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n489_), .A2(G43gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n485_), .A2(new_n488_), .A3(new_n214_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n561_), .B1(new_n563_), .B2(new_n562_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT84), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n561_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n562_), .A2(new_n563_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT84), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n564_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n534_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n567_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n574_), .A2(new_n571_), .A3(new_n570_), .A4(new_n564_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n516_), .A2(new_n517_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n511_), .A2(KEYINPUT32), .ZN(new_n580_));
  MUX2_X1   g379(.A(new_n579_), .B(new_n505_), .S(new_n580_), .Z(new_n581_));
  NAND2_X1  g380(.A1(new_n555_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n536_), .A2(new_n537_), .A3(new_n541_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n533_), .A2(new_n539_), .A3(new_n535_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n549_), .A3(new_n584_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n510_), .A2(new_n512_), .A3(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n553_), .B(KEYINPUT33), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n582_), .A2(new_n588_), .A3(new_n425_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n556_), .A2(new_n578_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT97), .B1(new_n543_), .B2(new_n549_), .ZN(new_n591_));
  AOI211_X1 g390(.A(new_n551_), .B(new_n548_), .C1(new_n540_), .C2(new_n542_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n553_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n578_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n594_), .A2(new_n515_), .A3(new_n520_), .A4(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT99), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n519_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT99), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n598_), .A2(new_n599_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n597_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n590_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n259_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n332_), .B(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(G229gat), .A3(G233gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n332_), .A2(new_n226_), .A3(new_n231_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT80), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n332_), .A2(new_n604_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n608_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n606_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G113gat), .B(G141gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(new_n432_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(new_n351_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n618_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n603_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n347_), .A2(KEYINPUT79), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n348_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(G1gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n627_), .A3(new_n555_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT38), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n268_), .A2(new_n275_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n603_), .A2(new_n630_), .ZN(new_n631_));
  OR4_X1    g430(.A1(KEYINPUT100), .A2(new_n320_), .A3(new_n622_), .A4(new_n346_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n320_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n621_), .A3(new_n345_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT100), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n631_), .A2(new_n632_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n627_), .B1(new_n636_), .B2(new_n555_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT101), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n629_), .A2(new_n638_), .ZN(G1324gat));
  OR3_X1    g438(.A1(new_n625_), .A2(G8gat), .A3(new_n598_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(KEYINPUT102), .A2(KEYINPUT39), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n631_), .A2(new_n632_), .A3(new_n635_), .ZN(new_n642_));
  OAI211_X1 g441(.A(G8gat), .B(new_n641_), .C1(new_n642_), .C2(new_n598_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(KEYINPUT102), .A2(KEYINPUT39), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n636_), .A2(new_n521_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n644_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n646_), .A2(G8gat), .A3(new_n641_), .A4(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n640_), .A2(new_n645_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT103), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n640_), .A2(new_n651_), .A3(new_n648_), .A4(new_n645_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n650_), .A2(KEYINPUT40), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT40), .B1(new_n650_), .B2(new_n652_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1325gat));
  INV_X1    g454(.A(new_n578_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n326_), .B1(new_n636_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT41), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n626_), .A2(new_n326_), .A3(new_n656_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT104), .ZN(G1326gat));
  XNOR2_X1  g460(.A(new_n425_), .B(KEYINPUT105), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G22gat), .B1(new_n642_), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT42), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n626_), .A2(new_n327_), .A3(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1327gat));
  AND2_X1   g466(.A1(new_n602_), .A2(new_n630_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n320_), .A2(new_n622_), .A3(new_n345_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n594_), .A2(G29gat), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT108), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n602_), .A2(new_n674_), .A3(new_n287_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n602_), .B2(new_n287_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n669_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT106), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n680_), .B(new_n669_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n678_), .A2(new_n679_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n678_), .A2(KEYINPUT107), .A3(new_n679_), .A4(new_n681_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n675_), .A2(new_n676_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(KEYINPUT44), .A3(new_n669_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n686_), .A2(new_n555_), .A3(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n673_), .B1(new_n689_), .B2(new_n215_), .ZN(G1328gat));
  NAND4_X1  g489(.A1(new_n684_), .A2(new_n521_), .A3(new_n688_), .A4(new_n685_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G36gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n670_), .A2(new_n216_), .A3(new_n521_), .ZN(new_n693_));
  XOR2_X1   g492(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n692_), .A2(KEYINPUT46), .A3(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1329gat));
  XNOR2_X1  g499(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n684_), .A2(new_n656_), .A3(new_n688_), .A4(new_n685_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G43gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n670_), .A2(new_n214_), .A3(new_n656_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n701_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n701_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n704_), .ZN(new_n707_));
  AOI211_X1 g506(.A(new_n706_), .B(new_n707_), .C1(new_n702_), .C2(G43gat), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n705_), .A2(new_n708_), .ZN(G1330gat));
  NAND4_X1  g508(.A1(new_n686_), .A2(KEYINPUT111), .A3(new_n426_), .A4(new_n688_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n684_), .A2(new_n426_), .A3(new_n688_), .A4(new_n685_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT111), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n710_), .A2(G50gat), .A3(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n670_), .A2(new_n209_), .A3(new_n662_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1331gat));
  NAND2_X1  g515(.A1(new_n320_), .A2(new_n622_), .ZN(new_n717_));
  NOR4_X1   g516(.A1(new_n603_), .A2(new_n717_), .A3(new_n287_), .A4(new_n346_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT112), .ZN(new_n719_));
  AOI21_X1  g518(.A(G57gat), .B1(new_n719_), .B2(new_n555_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n621_), .A2(new_n346_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR4_X1   g521(.A1(new_n603_), .A2(new_n633_), .A3(new_n630_), .A4(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n594_), .A2(new_n547_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(G1332gat));
  INV_X1    g524(.A(G64gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n723_), .B2(new_n521_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT48), .Z(new_n728_));
  NAND3_X1  g527(.A1(new_n719_), .A2(new_n726_), .A3(new_n521_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1333gat));
  INV_X1    g529(.A(G71gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n723_), .B2(new_n656_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT49), .Z(new_n733_));
  NAND3_X1  g532(.A1(new_n719_), .A2(new_n731_), .A3(new_n656_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT113), .ZN(G1334gat));
  INV_X1    g535(.A(G78gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n723_), .B2(new_n662_), .ZN(new_n738_));
  XOR2_X1   g537(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n719_), .A2(new_n737_), .A3(new_n662_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1335gat));
  NOR2_X1   g541(.A1(new_n717_), .A2(new_n345_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n668_), .A2(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G85gat), .B1(new_n744_), .B2(new_n555_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT115), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n687_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n687_), .A2(new_n746_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n743_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n555_), .A2(G85gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n745_), .B1(new_n749_), .B2(new_n750_), .ZN(G1336gat));
  AOI21_X1  g550(.A(G92gat), .B1(new_n744_), .B2(new_n521_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT116), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n747_), .A2(new_n748_), .A3(new_n743_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n521_), .A2(G92gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n753_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n756_), .B(new_n757_), .ZN(G1337gat));
  OAI21_X1  g557(.A(G99gat), .B1(new_n754_), .B2(new_n578_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n744_), .A2(new_n235_), .A3(new_n656_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g561(.A1(new_n687_), .A2(new_n426_), .A3(new_n743_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(G106gat), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT52), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n744_), .A2(new_n236_), .A3(new_n426_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT118), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g568(.A1(new_n521_), .A2(new_n594_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n595_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n287_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT119), .B1(new_n633_), .B2(new_n721_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n320_), .A2(new_n722_), .A3(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n772_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT54), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT120), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n315_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n304_), .B1(new_n297_), .B2(new_n302_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT55), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n305_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n297_), .A2(new_n302_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(KEYINPUT55), .A3(new_n303_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n786_), .A2(KEYINPUT56), .A3(new_n312_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT56), .B1(new_n786_), .B2(new_n312_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n780_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n605_), .A2(new_n613_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n618_), .B(new_n790_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n619_), .A2(new_n791_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n792_), .A2(new_n317_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n789_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n778_), .B(new_n779_), .C1(new_n794_), .C2(new_n630_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n630_), .B1(new_n789_), .B2(new_n793_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT57), .B1(new_n796_), .B2(KEYINPUT120), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n787_), .A2(new_n788_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n792_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n798_), .A2(KEYINPUT58), .A3(new_n314_), .A4(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n799_), .B(new_n314_), .C1(new_n788_), .C2(new_n787_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(new_n803_), .A3(new_n287_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n795_), .A2(new_n797_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n346_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n771_), .B1(new_n777_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G113gat), .B1(new_n807_), .B2(new_n621_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n776_), .B(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n806_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT59), .B1(new_n812_), .B2(new_n771_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT121), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n806_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n805_), .A2(KEYINPUT121), .A3(new_n346_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n777_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  INV_X1    g617(.A(new_n771_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n813_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n621_), .A2(G113gat), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT122), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n808_), .B1(new_n821_), .B2(new_n823_), .ZN(G1340gat));
  INV_X1    g623(.A(KEYINPUT60), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n633_), .B2(G120gat), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n807_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n813_), .A2(new_n820_), .A3(new_n827_), .A4(new_n320_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(G120gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(KEYINPUT60), .B2(new_n827_), .ZN(G1341gat));
  AOI21_X1  g629(.A(G127gat), .B1(new_n807_), .B2(new_n345_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n346_), .A2(new_n522_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n821_), .B2(new_n832_), .ZN(G1342gat));
  OAI211_X1 g632(.A(new_n630_), .B(new_n819_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n834_), .A2(KEYINPUT123), .A3(new_n523_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT123), .B1(new_n834_), .B2(new_n523_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT124), .B(G134gat), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n813_), .A2(new_n820_), .A3(new_n287_), .A4(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1343gat));
  NOR3_X1   g639(.A1(new_n812_), .A2(new_n656_), .A3(new_n425_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(new_n621_), .A3(new_n770_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g642(.A1(new_n841_), .A2(new_n320_), .A3(new_n770_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT125), .B(G148gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1345gat));
  NAND3_X1  g645(.A1(new_n841_), .A2(new_n345_), .A3(new_n770_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT61), .B(G155gat), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1346gat));
  AND2_X1   g648(.A1(new_n841_), .A2(new_n770_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n287_), .A2(G162gat), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n841_), .A2(new_n630_), .A3(new_n770_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n850_), .A2(new_n852_), .B1(new_n853_), .B2(new_n204_), .ZN(G1347gat));
  NOR2_X1   g653(.A1(new_n598_), .A2(new_n555_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n656_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n817_), .A2(new_n621_), .A3(new_n663_), .A4(new_n857_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n858_), .A2(G169gat), .ZN(new_n859_));
  INV_X1    g658(.A(new_n460_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT62), .B1(new_n859_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n858_), .A2(G169gat), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(G1348gat));
  AND3_X1   g665(.A1(new_n817_), .A2(new_n663_), .A3(new_n857_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n320_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n812_), .A2(new_n426_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n633_), .A2(new_n433_), .A3(new_n856_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n868_), .A2(new_n459_), .B1(new_n869_), .B2(new_n870_), .ZN(G1349gat));
  NAND3_X1  g670(.A1(new_n869_), .A2(new_n345_), .A3(new_n857_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n346_), .A2(new_n441_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n872_), .A2(new_n453_), .B1(new_n867_), .B2(new_n873_), .ZN(G1350gat));
  OAI21_X1  g673(.A(new_n630_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT126), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n867_), .A2(new_n876_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n867_), .A2(new_n287_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n454_), .ZN(G1351gat));
  AOI21_X1  g678(.A(new_n425_), .B1(new_n777_), .B2(new_n806_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(new_n578_), .A3(new_n855_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n622_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(new_n351_), .ZN(G1352gat));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n633_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(new_n349_), .ZN(G1353gat));
  NOR2_X1   g684(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n886_));
  AND2_X1   g685(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n887_));
  NOR4_X1   g686(.A1(new_n881_), .A2(new_n346_), .A3(new_n886_), .A4(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n886_), .B1(new_n881_), .B2(new_n346_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT127), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT127), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n891_), .B(new_n886_), .C1(new_n881_), .C2(new_n346_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n888_), .B1(new_n890_), .B2(new_n892_), .ZN(G1354gat));
  NOR3_X1   g692(.A1(new_n881_), .A2(new_n358_), .A3(new_n772_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n841_), .A2(new_n630_), .A3(new_n855_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n358_), .ZN(G1355gat));
endmodule


