//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n587_,
    new_n588_, new_n589_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT76), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT75), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G190gat), .B(G218gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G134gat), .B(G162gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT36), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT74), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G92gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G85gat), .ZN(new_n212_));
  OR3_X1    g011(.A1(new_n211_), .A2(KEYINPUT9), .A3(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G85gat), .B(G92gat), .Z(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT6), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n213_), .A2(new_n215_), .A3(new_n218_), .A4(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR3_X1   g024(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n223_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT7), .ZN(new_n228_));
  INV_X1    g027(.A(G99gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n217_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(KEYINPUT65), .A3(new_n224_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(new_n220_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n214_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n232_), .A2(KEYINPUT66), .A3(new_n214_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(KEYINPUT8), .A3(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n220_), .A2(new_n224_), .A3(new_n230_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT8), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(new_n214_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n222_), .B1(new_n237_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G29gat), .B(G36gat), .ZN(new_n242_));
  INV_X1    g041(.A(G50gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT71), .B(G43gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT73), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G232gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT34), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n248_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n246_), .B(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n247_), .B(new_n254_), .C1(new_n241_), .C2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n251_), .A2(new_n253_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n258_), .A2(new_n259_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n204_), .B(new_n209_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n257_), .A2(new_n241_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n259_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(new_n247_), .A4(new_n254_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n258_), .A2(new_n259_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT36), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .A4(new_n207_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n262_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n266_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n204_), .B1(new_n270_), .B2(new_n209_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT37), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n208_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT37), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n274_), .A3(new_n268_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n203_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n271_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(new_n268_), .A3(new_n262_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT76), .B1(new_n278_), .B2(KEYINPUT37), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G71gat), .B(G78gat), .Z(new_n281_));
  INV_X1    g080(.A(G57gat), .ZN(new_n282_));
  INV_X1    g081(.A(G64gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT11), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G57gat), .A2(G64gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n281_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n281_), .B2(new_n287_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n284_), .A2(new_n286_), .ZN(new_n292_));
  OAI22_X1  g091(.A1(new_n290_), .A2(new_n291_), .B1(new_n285_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n291_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n292_), .A2(new_n285_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n289_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G231gat), .A2(G233gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G8gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT77), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G15gat), .ZN(new_n303_));
  INV_X1    g102(.A(G22gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G15gat), .A2(G22gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G1gat), .A2(G8gat), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n305_), .A2(new_n306_), .B1(KEYINPUT14), .B2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n302_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n299_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT17), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G127gat), .B(G155gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT79), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT78), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G183gat), .B(G211gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT16), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n315_), .B(new_n317_), .ZN(new_n318_));
  OR3_X1    g117(.A1(new_n311_), .A2(new_n312_), .A3(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(KEYINPUT17), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n311_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n280_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT80), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT12), .ZN(new_n325_));
  INV_X1    g124(.A(new_n297_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n325_), .B1(new_n241_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G230gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n241_), .B2(new_n326_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n240_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n239_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n331_), .B1(new_n332_), .B2(new_n236_), .ZN(new_n333_));
  OAI211_X1 g132(.A(KEYINPUT12), .B(new_n297_), .C1(new_n333_), .C2(new_n222_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n327_), .A2(new_n330_), .A3(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n241_), .A2(new_n326_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n232_), .A2(KEYINPUT66), .A3(new_n214_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT66), .B1(new_n232_), .B2(new_n214_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n239_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n221_), .B(new_n326_), .C1(new_n339_), .C2(new_n331_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n241_), .A2(KEYINPUT68), .A3(new_n326_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n336_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n335_), .B1(new_n344_), .B2(new_n328_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G120gat), .B(G148gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(G204gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT5), .B(G176gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n345_), .A2(new_n350_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n335_), .B(new_n349_), .C1(new_n344_), .C2(new_n328_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT13), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(KEYINPUT69), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n354_), .A2(KEYINPUT69), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n353_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(KEYINPUT81), .B1(new_n324_), .B2(new_n359_), .ZN(new_n360_));
  OR2_X1    g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362_));
  INV_X1    g161(.A(G141gat), .ZN(new_n363_));
  INV_X1    g162(.A(G148gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT3), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT88), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT89), .B1(G141gat), .B2(G148gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT2), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n369_), .A2(KEYINPUT87), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n367_), .B(new_n372_), .C1(new_n371_), .C2(new_n370_), .ZN(new_n373_));
  OAI22_X1  g172(.A1(new_n366_), .A2(KEYINPUT88), .B1(KEYINPUT87), .B2(new_n369_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n361_), .B(new_n362_), .C1(new_n373_), .C2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n362_), .B(KEYINPUT1), .Z(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n361_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n365_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n380_), .A2(KEYINPUT95), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G127gat), .B(G134gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G113gat), .B(G120gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n381_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n381_), .A2(new_n385_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n386_), .A2(KEYINPUT4), .A3(new_n387_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n389_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n380_), .ZN(new_n393_));
  OR3_X1    g192(.A1(new_n393_), .A2(KEYINPUT4), .A3(new_n384_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n391_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(new_n212_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n400_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n390_), .A2(new_n395_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(G197gat), .B(G204gat), .Z(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT21), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G211gat), .B(G218gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT91), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n405_), .A2(KEYINPUT21), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(G169gat), .A2(G176gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G169gat), .A2(G176gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(KEYINPUT24), .A3(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT83), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G183gat), .A2(G190gat), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n417_), .B(KEYINPUT23), .Z(new_n418_));
  NOR2_X1   g217(.A1(new_n413_), .A2(KEYINPUT24), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT25), .B(G183gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT26), .B(G190gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n416_), .A2(new_n420_), .A3(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(KEYINPUT22), .B(G169gat), .Z(new_n425_));
  NOR2_X1   g224(.A1(G183gat), .A2(G190gat), .ZN(new_n426_));
  OAI221_X1 g225(.A(new_n414_), .B1(new_n425_), .B2(G176gat), .C1(new_n418_), .C2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT20), .B1(new_n412_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT92), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n423_), .A2(new_n415_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT93), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n420_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n427_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n412_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n429_), .A2(new_n430_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n431_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G226gat), .A2(G233gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT19), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n412_), .A2(new_n436_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT20), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n412_), .A2(new_n428_), .ZN(new_n445_));
  OR3_X1    g244(.A1(new_n444_), .A2(new_n441_), .A3(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(KEYINPUT94), .B(KEYINPUT18), .Z(new_n447_));
  XNOR2_X1  g246(.A(G8gat), .B(G36gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G64gat), .B(G92gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT32), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n442_), .A2(new_n446_), .A3(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n439_), .A2(new_n441_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n441_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT97), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n445_), .B1(new_n444_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n443_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n456_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(KEYINPUT32), .B(new_n452_), .C1(new_n455_), .C2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n404_), .A2(new_n454_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT98), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT98), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n404_), .A2(new_n464_), .A3(new_n454_), .A4(new_n461_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n442_), .A2(new_n446_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(new_n452_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n403_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT96), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n468_), .B1(new_n469_), .B2(KEYINPUT33), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n388_), .A2(new_n392_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n391_), .A2(new_n389_), .A3(new_n394_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n400_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(new_n470_), .A3(new_n473_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT33), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n463_), .B(new_n465_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(KEYINPUT29), .A2(new_n380_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT28), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G22gat), .B(G50gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT28), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n477_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n479_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G228gat), .A2(G233gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n487_), .B(KEYINPUT90), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT29), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n393_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G78gat), .B(G106gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n485_), .A2(new_n488_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n490_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n494_), .B1(new_n490_), .B2(new_n495_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT30), .B(G15gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n428_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT85), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G227gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n500_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G71gat), .B(G99gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(G43gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n384_), .B(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(new_n508_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n509_), .A2(KEYINPUT86), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT86), .B1(new_n509_), .B2(new_n510_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n498_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n476_), .A2(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n509_), .A2(new_n510_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n490_), .A2(new_n495_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n494_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n490_), .A2(new_n495_), .A3(new_n494_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n513_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n404_), .B(KEYINPUT99), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n442_), .A2(new_n446_), .A3(new_n452_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT100), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n451_), .B1(new_n455_), .B2(new_n460_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n526_), .A2(KEYINPUT100), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT27), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT27), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n467_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n524_), .A2(new_n525_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n516_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n246_), .A2(new_n309_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n537_), .B(new_n538_), .C1(new_n257_), .C2(new_n309_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n246_), .B(new_n309_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(G229gat), .A3(G233gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G113gat), .B(G141gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(G197gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT82), .B(G169gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n539_), .A2(new_n541_), .A3(new_n546_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n536_), .A2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n360_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n324_), .A2(KEYINPUT81), .A3(new_n359_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT101), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(KEYINPUT101), .A3(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n525_), .A2(G1gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n202_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n556_), .A2(KEYINPUT38), .A3(new_n557_), .A4(new_n559_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n359_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n550_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n536_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n273_), .A2(new_n268_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n322_), .A2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n525_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(G1gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT102), .Z(new_n574_));
  NAND3_X1  g373(.A1(new_n561_), .A2(new_n562_), .A3(new_n574_), .ZN(G1324gat));
  INV_X1    g374(.A(new_n534_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n570_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(G8gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT39), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n534_), .A2(G8gat), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n556_), .A2(new_n557_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT40), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n579_), .A2(new_n581_), .A3(KEYINPUT40), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(G1325gat));
  AOI21_X1  g385(.A(new_n303_), .B1(new_n570_), .B2(new_n514_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT41), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n514_), .A2(new_n303_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n588_), .B1(new_n558_), .B2(new_n589_), .ZN(G1326gat));
  AOI21_X1  g389(.A(new_n304_), .B1(new_n570_), .B2(new_n498_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT42), .Z(new_n592_));
  NAND2_X1  g391(.A1(new_n498_), .A2(new_n304_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT103), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n556_), .A2(new_n557_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT104), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT104), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(new_n595_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(G1327gat));
  INV_X1    g399(.A(new_n322_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n601_), .A2(new_n567_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n566_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(G29gat), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n571_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n536_), .A2(new_n280_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT43), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT43), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n536_), .A2(new_n608_), .A3(new_n280_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n565_), .A2(new_n322_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT44), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT44), .ZN(new_n614_));
  AOI211_X1 g413(.A(new_n614_), .B(new_n611_), .C1(new_n607_), .C2(new_n609_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n613_), .A2(new_n615_), .A3(new_n525_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT105), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G29gat), .B1(new_n616_), .B2(new_n617_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n605_), .B1(new_n618_), .B2(new_n619_), .ZN(G1328gat));
  INV_X1    g419(.A(G36gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n534_), .B(KEYINPUT106), .Z(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n603_), .A2(new_n621_), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT45), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n613_), .A2(new_n615_), .A3(new_n534_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n625_), .B1(new_n621_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT46), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n625_), .B(KEYINPUT46), .C1(new_n626_), .C2(new_n621_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1329gat));
  AOI21_X1  g430(.A(G43gat), .B1(new_n603_), .B2(new_n514_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT108), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT107), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n613_), .A2(new_n615_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n517_), .A2(G43gat), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n634_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  NOR4_X1   g437(.A1(new_n613_), .A2(new_n615_), .A3(KEYINPUT107), .A4(new_n636_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n633_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT47), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT47), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n633_), .B(new_n642_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(G1330gat));
  NAND3_X1  g443(.A1(new_n603_), .A2(new_n243_), .A3(new_n498_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n635_), .A2(new_n498_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n646_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT109), .B1(new_n646_), .B2(G50gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n645_), .B1(new_n647_), .B2(new_n648_), .ZN(G1331gat));
  NOR2_X1   g448(.A1(new_n359_), .A2(new_n550_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n516_), .B2(new_n535_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n569_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n653_), .A2(new_n282_), .A3(new_n525_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n324_), .A2(new_n652_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n571_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n654_), .B1(new_n657_), .B2(new_n282_), .ZN(G1332gat));
  OAI21_X1  g457(.A(G64gat), .B1(new_n653_), .B2(new_n622_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT48), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n656_), .A2(new_n283_), .A3(new_n623_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1333gat));
  OAI21_X1  g461(.A(G71gat), .B1(new_n653_), .B2(new_n513_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT49), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n513_), .A2(G71gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n655_), .B2(new_n665_), .ZN(G1334gat));
  INV_X1    g465(.A(new_n498_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G78gat), .B1(new_n653_), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT50), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n667_), .A2(G78gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n655_), .B2(new_n670_), .ZN(G1335gat));
  NAND2_X1  g470(.A1(new_n652_), .A2(new_n602_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT110), .Z(new_n673_));
  AOI21_X1  g472(.A(G85gat), .B1(new_n673_), .B2(new_n571_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT111), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n651_), .A2(new_n601_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n610_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n525_), .A2(new_n212_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT112), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n675_), .B1(new_n677_), .B2(new_n679_), .ZN(G1336gat));
  AOI21_X1  g479(.A(G92gat), .B1(new_n673_), .B2(new_n576_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n622_), .A2(new_n211_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n677_), .B2(new_n682_), .ZN(G1337gat));
  INV_X1    g482(.A(new_n677_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G99gat), .B1(new_n684_), .B2(new_n513_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n517_), .A2(new_n216_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT113), .ZN(new_n687_));
  AOI22_X1  g486(.A1(new_n673_), .A2(new_n686_), .B1(new_n687_), .B2(KEYINPUT51), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n687_), .A2(KEYINPUT51), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1338gat));
  NAND3_X1  g490(.A1(new_n673_), .A2(new_n217_), .A3(new_n498_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT52), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n677_), .A2(new_n498_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(G106gat), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT52), .B(new_n217_), .C1(new_n677_), .C2(new_n498_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT53), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT53), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n699_), .B(new_n692_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1339gat));
  INV_X1    g500(.A(KEYINPUT116), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT115), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n546_), .B1(new_n540_), .B2(new_n537_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n538_), .B1(new_n257_), .B2(new_n309_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(new_n537_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n549_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n703_), .B1(new_n353_), .B2(new_n708_), .ZN(new_n709_));
  AOI211_X1 g508(.A(KEYINPUT115), .B(new_n707_), .C1(new_n351_), .C2(new_n352_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT114), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n550_), .A2(new_n352_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT68), .B1(new_n241_), .B2(new_n326_), .ZN(new_n714_));
  NOR4_X1   g513(.A1(new_n333_), .A2(new_n341_), .A3(new_n222_), .A4(new_n297_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n327_), .A2(new_n334_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n329_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n327_), .A2(new_n330_), .A3(KEYINPUT55), .A4(new_n334_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT55), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n335_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n718_), .A2(new_n719_), .A3(new_n721_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n722_), .A2(KEYINPUT56), .A3(new_n350_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT56), .B1(new_n722_), .B2(new_n350_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n712_), .B(new_n713_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n711_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n722_), .A2(new_n350_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT56), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n722_), .A2(KEYINPUT56), .A3(new_n350_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n712_), .B1(new_n731_), .B2(new_n713_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n567_), .B1(new_n726_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT57), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n708_), .A2(new_n352_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT58), .B1(new_n731_), .B2(new_n735_), .ZN(new_n736_));
  OAI211_X1 g535(.A(KEYINPUT58), .B(new_n735_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n733_), .A2(new_n734_), .B1(new_n739_), .B2(new_n280_), .ZN(new_n740_));
  OAI211_X1 g539(.A(KEYINPUT57), .B(new_n567_), .C1(new_n726_), .C2(new_n732_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n601_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n550_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n601_), .B(new_n743_), .C1(new_n276_), .C2(new_n279_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT54), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n702_), .B1(new_n742_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n733_), .A2(new_n734_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n739_), .A2(new_n280_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n741_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n322_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n744_), .B(KEYINPUT54), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(KEYINPUT116), .A3(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n576_), .A2(new_n518_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n747_), .A2(new_n753_), .A3(new_n571_), .A4(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT59), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n742_), .A2(new_n746_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n525_), .A2(KEYINPUT59), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n754_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n751_), .A2(new_n752_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n762_), .A2(KEYINPUT117), .A3(new_n754_), .A4(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n756_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(G113gat), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n564_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n755_), .A2(new_n564_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(new_n768_), .ZN(G1340gat));
  OAI21_X1  g568(.A(KEYINPUT118), .B1(new_n765_), .B2(new_n359_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(G120gat), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n765_), .A2(KEYINPUT118), .A3(new_n359_), .ZN(new_n772_));
  INV_X1    g571(.A(G120gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n773_), .B1(new_n359_), .B2(KEYINPUT60), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(KEYINPUT60), .B2(new_n773_), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n771_), .A2(new_n772_), .B1(new_n755_), .B2(new_n775_), .ZN(G1341gat));
  NAND4_X1  g575(.A1(new_n756_), .A2(G127gat), .A3(new_n764_), .A4(new_n601_), .ZN(new_n777_));
  INV_X1    g576(.A(G127gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(new_n755_), .B2(new_n322_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT119), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(G1342gat));
  NAND2_X1  g581(.A1(new_n280_), .A2(G134gat), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n755_), .A2(new_n567_), .ZN(new_n784_));
  OAI22_X1  g583(.A1(new_n765_), .A2(new_n783_), .B1(G134gat), .B2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT120), .ZN(G1343gat));
  NOR2_X1   g585(.A1(new_n623_), .A2(new_n523_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n747_), .A2(new_n753_), .A3(new_n571_), .A4(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT121), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n789_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n564_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(new_n363_), .ZN(G1344gat));
  AOI21_X1  g592(.A(new_n359_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(new_n364_), .ZN(G1345gat));
  NAND2_X1  g594(.A1(new_n790_), .A2(new_n791_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT61), .B(G155gat), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n796_), .A2(new_n601_), .A3(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n796_), .B2(new_n601_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(G1346gat));
  AOI21_X1  g599(.A(G162gat), .B1(new_n796_), .B2(new_n568_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n280_), .A2(G162gat), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT122), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n801_), .B1(new_n796_), .B2(new_n803_), .ZN(G1347gat));
  NAND3_X1  g603(.A1(new_n623_), .A2(new_n514_), .A3(new_n525_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n758_), .A2(new_n498_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n550_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n807_), .A2(G169gat), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n808_), .A2(KEYINPUT62), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(KEYINPUT62), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n809_), .B(new_n810_), .C1(new_n425_), .C2(new_n807_), .ZN(G1348gat));
  INV_X1    g610(.A(G176gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n747_), .A2(new_n753_), .A3(new_n667_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT123), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT123), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n747_), .A2(new_n753_), .A3(new_n815_), .A4(new_n667_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n805_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n812_), .B1(new_n817_), .B2(new_n563_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n806_), .A2(new_n812_), .A3(new_n563_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT124), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT124), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n359_), .B(new_n805_), .C1(new_n814_), .C2(new_n816_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n822_), .B(new_n819_), .C1(new_n823_), .C2(new_n812_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n821_), .A2(new_n824_), .ZN(G1349gat));
  AOI21_X1  g624(.A(G183gat), .B1(new_n817_), .B2(new_n601_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n322_), .A2(new_n421_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n806_), .B2(new_n827_), .ZN(G1350gat));
  NAND2_X1  g627(.A1(new_n806_), .A2(new_n280_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n568_), .A2(new_n422_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n829_), .A2(G190gat), .B1(new_n806_), .B2(new_n830_), .ZN(new_n831_));
  XOR2_X1   g630(.A(new_n831_), .B(KEYINPUT125), .Z(G1351gat));
  NAND2_X1  g631(.A1(new_n747_), .A2(new_n753_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n571_), .A2(new_n523_), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT126), .Z(new_n835_));
  NOR3_X1   g634(.A1(new_n833_), .A2(new_n622_), .A3(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n550_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n563_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g639(.A1(new_n836_), .A2(new_n601_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT63), .B(G211gat), .Z(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n841_), .B2(new_n843_), .ZN(G1354gat));
  XNOR2_X1  g643(.A(KEYINPUT127), .B(G218gat), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(new_n836_), .B2(new_n568_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n280_), .A2(new_n845_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n836_), .B2(new_n847_), .ZN(G1355gat));
endmodule


