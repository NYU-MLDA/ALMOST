//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_;
  INV_X1    g000(.A(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(G8gat), .ZN(new_n203_));
  INV_X1    g002(.A(G36gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G8gat), .A2(G36gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT18), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G64gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n207_), .A2(new_n208_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n211_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n202_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n215_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G92gat), .A3(new_n213_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n218_), .A3(KEYINPUT32), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G226gat), .A2(G233gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT19), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT25), .B(G183gat), .ZN(new_n222_));
  INV_X1    g021(.A(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT26), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT82), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G190gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n225_), .B1(new_n224_), .B2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G183gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT23), .B1(new_n232_), .B2(new_n223_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(G183gat), .A3(G190gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(KEYINPUT24), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT24), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n236_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n231_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT87), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n233_), .A2(new_n245_), .A3(new_n235_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n232_), .A2(new_n223_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n234_), .A2(KEYINPUT87), .A3(G183gat), .A4(G190gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n249_), .A2(new_n239_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT84), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT83), .B(G169gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT22), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n251_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT86), .B(G176gat), .Z(new_n255_));
  INV_X1    g054(.A(KEYINPUT83), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(G169gat), .ZN(new_n257_));
  INV_X1    g056(.A(G169gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(KEYINPUT83), .ZN(new_n259_));
  OAI211_X1 g058(.A(KEYINPUT84), .B(KEYINPUT22), .C1(new_n257_), .C2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(KEYINPUT85), .B2(new_n253_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(KEYINPUT85), .B2(new_n253_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n254_), .A2(new_n255_), .A3(new_n260_), .A4(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n244_), .B1(new_n250_), .B2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G197gat), .B(G204gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n265_), .B1(KEYINPUT21), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(KEYINPUT21), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT20), .B1(new_n264_), .B2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n246_), .A2(new_n248_), .A3(new_n242_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT95), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n224_), .A2(new_n229_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n222_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n274_), .A2(new_n240_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT95), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n246_), .A2(new_n276_), .A3(new_n248_), .A4(new_n242_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n272_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n236_), .A2(new_n247_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT22), .B(G169gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT96), .ZN(new_n281_));
  INV_X1    g080(.A(new_n255_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n239_), .B(new_n279_), .C1(new_n281_), .C2(new_n282_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n278_), .A2(new_n269_), .A3(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n221_), .B1(new_n270_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT20), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(new_n264_), .B2(new_n269_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n278_), .A2(new_n283_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n269_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n221_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n287_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n219_), .B1(new_n285_), .B2(new_n292_), .ZN(new_n293_));
  NOR3_X1   g092(.A1(new_n270_), .A2(new_n284_), .A3(new_n221_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n291_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT101), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n219_), .B(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n293_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n300_), .B(KEYINPUT98), .Z(new_n301_));
  NAND2_X1  g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT90), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT2), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT2), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n307_));
  OAI22_X1  g106(.A1(KEYINPUT89), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .A4(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n302_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n318_), .A2(new_n319_), .A3(new_n309_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n313_), .A2(new_n317_), .A3(new_n314_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n316_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT91), .ZN(new_n324_));
  XOR2_X1   g123(.A(G127gat), .B(G134gat), .Z(new_n325_));
  XOR2_X1   g124(.A(G113gat), .B(G120gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n312_), .A2(new_n315_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT91), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n324_), .A2(new_n328_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n327_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n301_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(KEYINPUT4), .A3(new_n333_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n329_), .B(KEYINPUT91), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT99), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n327_), .A2(KEYINPUT4), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n324_), .A2(new_n331_), .A3(new_n338_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT99), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n335_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n334_), .B1(new_n342_), .B2(new_n301_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G57gat), .B(G85gat), .Z(new_n344_));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n343_), .A2(new_n349_), .ZN(new_n350_));
  AOI211_X1 g149(.A(new_n348_), .B(new_n334_), .C1(new_n342_), .C2(new_n301_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n299_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT102), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n216_), .A2(new_n218_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT97), .ZN(new_n356_));
  INV_X1    g155(.A(new_n244_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n263_), .A2(new_n239_), .A3(new_n249_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT20), .B1(new_n359_), .B2(new_n289_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n269_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n221_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n354_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n286_), .B1(new_n359_), .B2(new_n289_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n278_), .A2(new_n269_), .A3(new_n283_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n291_), .A3(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n362_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n355_), .A2(new_n356_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n296_), .A2(KEYINPUT97), .A3(new_n363_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n342_), .A2(new_n301_), .ZN(new_n371_));
  OAI211_X1 g170(.A(KEYINPUT33), .B(new_n348_), .C1(new_n371_), .C2(new_n334_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n332_), .A2(new_n333_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n348_), .B1(new_n373_), .B2(new_n301_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n374_), .B1(new_n301_), .B2(new_n342_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT33), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n343_), .B2(new_n349_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n370_), .A2(new_n372_), .A3(new_n375_), .A4(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT102), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n299_), .B(new_n379_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n353_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n327_), .B(KEYINPUT31), .Z(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT30), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n359_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n264_), .A2(KEYINPUT30), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G15gat), .B(G43gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(new_n386_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n389_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n357_), .A2(new_n358_), .A3(KEYINPUT30), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT30), .B1(new_n357_), .B2(new_n358_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n391_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G71gat), .B(G99gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n390_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT88), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n395_), .B1(new_n390_), .B2(new_n394_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n383_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n399_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n401_), .A2(new_n397_), .A3(new_n396_), .A4(new_n382_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n405_));
  OR3_X1    g204(.A1(new_n329_), .A2(KEYINPUT94), .A3(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT94), .B1(new_n329_), .B2(new_n405_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n289_), .A3(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n324_), .A2(KEYINPUT29), .A3(new_n331_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n269_), .A2(new_n409_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n408_), .A2(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n336_), .B2(KEYINPUT29), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n324_), .A2(new_n331_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT29), .ZN(new_n416_));
  INV_X1    g215(.A(new_n413_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n414_), .A2(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n412_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G78gat), .B(G106gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G22gat), .B(G50gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n412_), .A2(new_n419_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n420_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n423_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n412_), .A2(new_n419_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n412_), .A2(new_n419_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n404_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n381_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n403_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n425_), .A2(new_n429_), .A3(new_n400_), .A4(new_n402_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n350_), .A2(new_n351_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT27), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n368_), .A2(new_n437_), .A3(new_n369_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n285_), .A2(new_n292_), .ZN(new_n439_));
  OAI211_X1 g238(.A(KEYINPUT27), .B(new_n367_), .C1(new_n439_), .C2(new_n363_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n436_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n432_), .A2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT75), .B(G1gat), .Z(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT76), .B(G8gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT14), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G15gat), .B(G22gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G1gat), .B(G8gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT77), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n449_), .B(KEYINPUT77), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G29gat), .B(G36gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G43gat), .B(G50gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT79), .B1(new_n455_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT79), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n452_), .A2(new_n454_), .A3(new_n461_), .A4(new_n458_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n455_), .A2(new_n459_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G229gat), .A2(G233gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT15), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n458_), .A2(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n456_), .A2(new_n457_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n456_), .A2(new_n457_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(KEYINPUT15), .A3(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n467_), .B1(new_n474_), .B2(new_n455_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n463_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT80), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT80), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n463_), .A2(new_n478_), .A3(new_n475_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n468_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G113gat), .B(G141gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(G169gat), .ZN(new_n482_));
  INV_X1    g281(.A(G197gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT81), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n480_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n468_), .A2(new_n477_), .A3(new_n488_), .A4(new_n479_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n443_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT103), .ZN(new_n492_));
  INV_X1    g291(.A(new_n436_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G190gat), .B(G218gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(G134gat), .B(G162gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n498_), .A2(new_n499_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G232gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT34), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT35), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G85gat), .A2(G92gat), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n515_), .A2(KEYINPUT9), .ZN(new_n516_));
  OR2_X1    g315(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n517_));
  INV_X1    g316(.A(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(G85gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n202_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(KEYINPUT9), .A3(new_n515_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n514_), .A2(new_n516_), .A3(new_n520_), .A4(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT8), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT66), .ZN(new_n526_));
  AND2_X1   g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527_));
  NOR2_X1   g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n522_), .A2(KEYINPUT66), .A3(new_n515_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT7), .ZN(new_n532_));
  INV_X1    g331(.A(G99gat), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n518_), .A4(KEYINPUT65), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT65), .ZN(new_n535_));
  OAI22_X1  g334(.A1(new_n535_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n534_), .A2(new_n536_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n525_), .B1(new_n531_), .B2(new_n537_), .ZN(new_n538_));
  AND4_X1   g337(.A1(new_n525_), .A2(new_n537_), .A3(new_n529_), .A4(new_n530_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n524_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n474_), .A2(new_n540_), .A3(KEYINPUT71), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT71), .ZN(new_n542_));
  INV_X1    g341(.A(new_n524_), .ZN(new_n543_));
  AND4_X1   g342(.A1(new_n512_), .A2(new_n534_), .A3(new_n513_), .A4(new_n536_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n529_), .A2(new_n530_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT8), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n531_), .A2(new_n525_), .A3(new_n537_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n543_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n470_), .A2(new_n473_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n542_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n541_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n509_), .B1(new_n551_), .B2(KEYINPUT72), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n548_), .A2(new_n458_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n506_), .A2(new_n507_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n541_), .A2(new_n550_), .B1(new_n458_), .B2(new_n548_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT72), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n541_), .B2(new_n550_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n557_), .A2(new_n559_), .A3(new_n509_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n501_), .B(new_n503_), .C1(new_n556_), .C2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n557_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n552_), .A2(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n557_), .B(new_n554_), .C1(new_n559_), .C2(new_n509_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n563_), .A2(new_n564_), .A3(new_n499_), .A4(new_n498_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n561_), .A2(KEYINPUT37), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT37), .B1(new_n561_), .B2(new_n565_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G230gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT64), .ZN(new_n570_));
  XOR2_X1   g369(.A(G71gat), .B(G78gat), .Z(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G57gat), .B(G64gat), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(KEYINPUT11), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(KEYINPUT11), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT11), .ZN(new_n576_));
  INV_X1    g375(.A(G57gat), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n577_), .A2(G64gat), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n211_), .A2(G57gat), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n576_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n575_), .A2(new_n580_), .A3(new_n571_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n574_), .A2(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n524_), .B(new_n582_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n570_), .B1(new_n584_), .B2(KEYINPUT67), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT67), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n548_), .B2(new_n582_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n584_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT12), .ZN(new_n589_));
  INV_X1    g388(.A(new_n582_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n540_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT12), .B1(new_n548_), .B2(new_n582_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n583_), .A2(new_n570_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT68), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n583_), .A2(KEYINPUT68), .A3(new_n570_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n593_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n588_), .A2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(G176gat), .B(G204gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(G120gat), .B(G148gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n599_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n588_), .A2(new_n598_), .A3(new_n604_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT13), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(KEYINPUT70), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n610_), .B1(new_n608_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n568_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n582_), .B(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(new_n455_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G127gat), .B(G155gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT17), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n622_), .A2(KEYINPUT17), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n617_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n617_), .A2(new_n623_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n614_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n492_), .A2(new_n493_), .A3(new_n444_), .A4(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT104), .B1(new_n613_), .B2(new_n490_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n613_), .A2(KEYINPUT104), .A3(new_n490_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n634_), .A2(new_n627_), .A3(new_n635_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n381_), .A2(new_n431_), .B1(new_n435_), .B2(new_n441_), .ZN(new_n637_));
  AOI211_X1 g436(.A(new_n500_), .B(new_n502_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n565_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n636_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n436_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n630_), .A2(new_n631_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n632_), .A2(new_n643_), .A3(new_n644_), .ZN(G1324gat));
  INV_X1    g444(.A(KEYINPUT106), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n438_), .A2(new_n440_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n636_), .A2(new_n641_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n203_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n636_), .A2(new_n641_), .A3(KEYINPUT105), .A4(new_n648_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n646_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n651_), .A2(new_n652_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(KEYINPUT106), .B2(new_n656_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n492_), .A2(new_n648_), .A3(new_n445_), .A4(new_n629_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n653_), .A2(new_n654_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n657_), .A2(KEYINPUT40), .A3(new_n658_), .A4(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n656_), .A2(KEYINPUT106), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n662_), .A2(new_n654_), .A3(new_n653_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n659_), .A2(new_n658_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n660_), .A2(new_n665_), .ZN(G1325gat));
  OAI21_X1  g465(.A(G15gat), .B1(new_n642_), .B2(new_n403_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT41), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n492_), .A2(new_n629_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n669_), .A2(G15gat), .A3(new_n403_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n668_), .A2(new_n670_), .ZN(G1326gat));
  INV_X1    g470(.A(new_n430_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G22gat), .B1(new_n642_), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT42), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n672_), .A2(G22gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n669_), .B2(new_n675_), .ZN(G1327gat));
  INV_X1    g475(.A(new_n613_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n640_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n677_), .A2(new_n627_), .A3(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n492_), .A2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n493_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n634_), .A2(new_n628_), .A3(new_n635_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n684_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT37), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n561_), .A2(KEYINPUT37), .A3(new_n565_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(KEYINPUT107), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n685_), .A2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT43), .B1(new_n637_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n687_), .A2(new_n688_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n443_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n683_), .B1(new_n691_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n682_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  AOI211_X1 g498(.A(KEYINPUT108), .B(new_n683_), .C1(new_n691_), .C2(new_n696_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT109), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n694_), .B1(new_n432_), .B2(new_n442_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n685_), .A2(new_n689_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n443_), .A2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n702_), .B1(new_n704_), .B2(KEYINPUT43), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT108), .B1(new_n705_), .B2(new_n683_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n697_), .A2(new_n698_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n682_), .A4(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n701_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n697_), .A2(KEYINPUT44), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n711_), .A2(G29gat), .A3(new_n493_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n681_), .B1(new_n710_), .B2(new_n712_), .ZN(G1328gat));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n648_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n204_), .B1(new_n710_), .B2(new_n716_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n492_), .A2(new_n204_), .A3(new_n648_), .A4(new_n679_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n714_), .B1(new_n717_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n718_), .B(KEYINPUT45), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n715_), .B1(new_n701_), .B2(new_n709_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n722_), .B(KEYINPUT46), .C1(new_n723_), .C2(new_n204_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(G1329gat));
  NAND3_X1  g524(.A1(new_n711_), .A2(G43gat), .A3(new_n404_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n701_), .B2(new_n709_), .ZN(new_n727_));
  XOR2_X1   g526(.A(KEYINPUT110), .B(G43gat), .Z(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n680_), .B2(new_n404_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OR3_X1    g530(.A1(new_n727_), .A2(new_n729_), .A3(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1330gat));
  AOI21_X1  g533(.A(G50gat), .B1(new_n680_), .B2(new_n430_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n711_), .A2(G50gat), .A3(new_n430_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n710_), .B2(new_n736_), .ZN(G1331gat));
  NOR3_X1   g536(.A1(new_n637_), .A2(new_n490_), .A3(new_n613_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n738_), .A2(new_n627_), .A3(new_n568_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(new_n577_), .A3(new_n493_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n487_), .A2(new_n489_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n641_), .A2(new_n741_), .A3(new_n627_), .A4(new_n677_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G57gat), .B1(new_n742_), .B2(new_n436_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n743_), .ZN(G1332gat));
  OAI21_X1  g543(.A(G64gat), .B1(new_n742_), .B2(new_n647_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT48), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n739_), .A2(new_n211_), .A3(new_n648_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1333gat));
  OAI21_X1  g547(.A(G71gat), .B1(new_n742_), .B2(new_n403_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT49), .ZN(new_n750_));
  INV_X1    g549(.A(G71gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n739_), .A2(new_n751_), .A3(new_n404_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1334gat));
  OAI21_X1  g552(.A(G78gat), .B1(new_n742_), .B2(new_n672_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT50), .ZN(new_n755_));
  INV_X1    g554(.A(G78gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n739_), .A2(new_n756_), .A3(new_n430_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1335gat));
  NAND3_X1  g557(.A1(new_n677_), .A2(new_n741_), .A3(new_n628_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n691_), .B2(new_n696_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n761_), .A2(new_n521_), .A3(new_n436_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n678_), .A2(new_n627_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n738_), .A2(KEYINPUT112), .A3(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n443_), .A2(new_n741_), .A3(new_n677_), .A4(new_n763_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G85gat), .B1(new_n768_), .B2(new_n493_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n770_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n762_), .B1(new_n771_), .B2(new_n772_), .ZN(G1336gat));
  OAI21_X1  g572(.A(G92gat), .B1(new_n761_), .B2(new_n647_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n768_), .A2(new_n202_), .A3(new_n648_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1337gat));
  AOI21_X1  g575(.A(new_n533_), .B1(new_n760_), .B2(new_n404_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n404_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n768_), .B2(new_n778_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(G106gat), .C1(new_n761_), .C2(new_n672_), .ZN(new_n782_));
  AOI211_X1 g581(.A(new_n672_), .B(new_n759_), .C1(new_n691_), .C2(new_n696_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT52), .B1(new_n783_), .B2(new_n518_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n672_), .A2(G106gat), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n764_), .B2(new_n767_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT114), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n785_), .A2(new_n792_), .A3(new_n789_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(KEYINPUT53), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n792_), .B1(new_n785_), .B2(new_n789_), .ZN(new_n796_));
  AOI211_X1 g595(.A(KEYINPUT114), .B(new_n788_), .C1(new_n782_), .C2(new_n784_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n794_), .A2(new_n798_), .ZN(G1339gat));
  NOR2_X1   g598(.A1(new_n692_), .A2(new_n677_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT115), .B1(new_n490_), .B2(new_n628_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n741_), .A2(new_n802_), .A3(new_n627_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n800_), .A2(KEYINPUT54), .A3(new_n801_), .A4(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n801_), .A2(new_n803_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n614_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n589_), .B1(new_n540_), .B2(new_n590_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n548_), .A2(KEYINPUT12), .A3(new_n582_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n583_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n570_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT116), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n584_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n570_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n813_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n598_), .A2(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n593_), .A2(new_n596_), .A3(KEYINPUT55), .A4(new_n597_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n605_), .B1(new_n817_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT56), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT56), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n824_), .B(new_n605_), .C1(new_n817_), .C2(new_n821_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n823_), .A2(new_n490_), .A3(new_n607_), .A4(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n480_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n460_), .A2(new_n462_), .B1(new_n455_), .B2(new_n459_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n485_), .B1(new_n828_), .B2(new_n467_), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n829_), .A2(KEYINPUT117), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n466_), .B1(new_n474_), .B2(new_n455_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n829_), .A2(KEYINPUT117), .B1(new_n463_), .B2(new_n831_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n484_), .A2(new_n827_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n608_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n826_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n678_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n640_), .B1(new_n826_), .B2(new_n834_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT57), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n823_), .A2(new_n833_), .A3(new_n607_), .A4(new_n825_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n607_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n822_), .B2(KEYINPUT56), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n845_), .A2(KEYINPUT58), .A3(new_n833_), .A4(new_n825_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(new_n692_), .A3(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n838_), .A2(new_n840_), .A3(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n808_), .B1(new_n848_), .B2(new_n628_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n434_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n647_), .A3(new_n493_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n852_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT59), .B1(new_n849_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n843_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n846_), .A2(new_n692_), .ZN(new_n858_));
  OAI22_X1  g657(.A1(new_n857_), .A2(new_n858_), .B1(new_n839_), .B2(KEYINPUT57), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n839_), .A2(KEYINPUT57), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n628_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n808_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864_));
  INV_X1    g663(.A(new_n855_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n856_), .A2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(G113gat), .B1(new_n867_), .B2(new_n741_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n863_), .A2(new_n865_), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n741_), .A2(G113gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(G1340gat));
  NAND3_X1  g670(.A1(new_n856_), .A2(new_n866_), .A3(new_n677_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G120gat), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n874_));
  AOI21_X1  g673(.A(G120gat), .B1(new_n677_), .B2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n874_), .B2(G120gat), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT119), .B1(new_n869_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n863_), .A2(new_n879_), .A3(new_n865_), .A4(new_n876_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n873_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n873_), .A2(new_n881_), .A3(KEYINPUT120), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1341gat));
  OAI21_X1  g685(.A(G127gat), .B1(new_n867_), .B2(new_n628_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n628_), .A2(G127gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n869_), .B2(new_n888_), .ZN(G1342gat));
  OAI21_X1  g688(.A(G134gat), .B1(new_n867_), .B2(new_n568_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n678_), .A2(G134gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n869_), .B2(new_n891_), .ZN(G1343gat));
  NOR3_X1   g691(.A1(new_n648_), .A2(new_n436_), .A3(new_n433_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n490_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n677_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n895_), .B2(new_n627_), .ZN(new_n901_));
  NOR4_X1   g700(.A1(new_n849_), .A2(KEYINPUT121), .A3(new_n628_), .A4(new_n894_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT61), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n863_), .A2(new_n627_), .A3(new_n893_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT121), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n895_), .A2(new_n900_), .A3(new_n627_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n903_), .A2(G155gat), .A3(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(G155gat), .B1(new_n903_), .B2(new_n908_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1346gat));
  AOI21_X1  g710(.A(G162gat), .B1(new_n895_), .B2(new_n640_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n703_), .A2(G162gat), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n895_), .B2(new_n913_), .ZN(G1347gat));
  NOR2_X1   g713(.A1(new_n647_), .A2(new_n493_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n863_), .A2(new_n850_), .A3(new_n490_), .A4(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n916_), .A2(new_n917_), .A3(G169gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n917_), .B1(new_n916_), .B2(G169gat), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n918_), .A2(new_n919_), .ZN(new_n922_));
  OAI221_X1 g721(.A(new_n920_), .B1(new_n281_), .B2(new_n916_), .C1(new_n921_), .C2(new_n922_), .ZN(G1348gat));
  AND3_X1   g722(.A1(new_n863_), .A2(new_n850_), .A3(new_n915_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n924_), .A2(new_n925_), .A3(G176gat), .A4(new_n677_), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n863_), .A2(new_n850_), .A3(new_n677_), .A4(new_n915_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n255_), .ZN(new_n928_));
  INV_X1    g727(.A(G176gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(KEYINPUT124), .B1(new_n927_), .B2(new_n929_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n926_), .A2(new_n928_), .A3(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n926_), .A2(KEYINPUT125), .A3(new_n930_), .A4(new_n928_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1349gat));
  NAND2_X1  g734(.A1(new_n924_), .A2(new_n627_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(G183gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n222_), .B1(KEYINPUT126), .B2(G183gat), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n936_), .B2(new_n939_), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n924_), .A2(new_n273_), .A3(new_n640_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n863_), .A2(new_n915_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n942_), .A2(new_n434_), .A3(new_n568_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n941_), .B1(new_n943_), .B2(new_n223_), .ZN(G1351gat));
  NOR2_X1   g743(.A1(new_n942_), .A2(new_n433_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n490_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n677_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n950_));
  INV_X1    g749(.A(G211gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n627_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n952_));
  XOR2_X1   g751(.A(new_n952_), .B(KEYINPUT127), .Z(new_n953_));
  NAND2_X1  g752(.A1(new_n945_), .A2(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n950_), .A2(new_n951_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n954_), .B(new_n955_), .ZN(G1354gat));
  INV_X1    g755(.A(G218gat), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n945_), .A2(new_n957_), .A3(new_n640_), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n942_), .A2(new_n433_), .A3(new_n568_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n959_), .B2(new_n957_), .ZN(G1355gat));
endmodule


