//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_;
  AND2_X1   g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT83), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  INV_X1    g004(.A(G204gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G197gat), .A2(G204gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(KEYINPUT21), .A3(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212_));
  INV_X1    g011(.A(new_n208_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G197gat), .A2(G204gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G155gat), .ZN(new_n219_));
  INV_X1    g018(.A(G162gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT80), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT80), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(G155gat), .B2(G162gat), .ZN(new_n223_));
  AOI22_X1  g022(.A1(new_n221_), .A2(new_n223_), .B1(G155gat), .B2(G162gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT2), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n228_));
  NOR3_X1   g027(.A1(KEYINPUT81), .A2(G141gat), .A3(G148gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n227_), .B(new_n228_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G141gat), .A2(G148gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT81), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(KEYINPUT3), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n224_), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G141gat), .B(G148gat), .Z(new_n237_));
  NOR3_X1   g036(.A1(new_n222_), .A2(G155gat), .A3(G162gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT80), .B1(new_n219_), .B2(new_n220_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT1), .B1(new_n219_), .B2(new_n220_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(G155gat), .A3(G162gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n237_), .B1(new_n240_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n236_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n218_), .B1(KEYINPUT29), .B2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n202_), .A2(new_n203_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n247_), .A2(new_n249_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n204_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G22gat), .B(G50gat), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT29), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n236_), .A2(new_n245_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT28), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT82), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n236_), .A2(new_n245_), .A3(new_n259_), .A4(new_n255_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n257_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n258_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n254_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n234_), .A2(KEYINPUT3), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n229_), .A2(new_n230_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n241_), .B(new_n243_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n266_), .A2(new_n224_), .B1(new_n267_), .B2(new_n237_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n259_), .B1(new_n268_), .B2(new_n255_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n260_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT82), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n257_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n253_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n263_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT84), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n252_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G78gat), .B(G106gat), .Z(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n263_), .A2(new_n273_), .A3(KEYINPUT84), .A4(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n263_), .A2(KEYINPUT84), .A3(new_n273_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n277_), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n276_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n274_), .A2(new_n275_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n252_), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n281_), .A2(new_n279_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G127gat), .B(G134gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G113gat), .B(G120gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n268_), .A2(new_n291_), .A3(KEYINPUT93), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n236_), .A2(new_n245_), .A3(KEYINPUT93), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n290_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n287_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT96), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n246_), .A2(new_n291_), .A3(new_n287_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OR3_X1    g098(.A1(new_n295_), .A2(new_n296_), .A3(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n296_), .B1(new_n295_), .B2(new_n299_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G1gat), .B(G29gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G57gat), .B(G85gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n292_), .A2(new_n294_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n298_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n300_), .A2(new_n301_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n291_), .B1(new_n268_), .B2(KEYINPUT93), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n293_), .A2(new_n290_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n298_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n297_), .A2(new_n308_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n313_), .B(new_n306_), .C1(new_n295_), .C2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT95), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n315_), .A2(new_n316_), .A3(KEYINPUT33), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT33), .B1(new_n315_), .B2(new_n316_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n310_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT89), .ZN(new_n320_));
  INV_X1    g119(.A(G183gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT25), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G183gat), .ZN(new_n324_));
  INV_X1    g123(.A(G190gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT26), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT26), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G190gat), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n322_), .A2(new_n324_), .A3(new_n326_), .A4(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT24), .ZN(new_n330_));
  INV_X1    g129(.A(G169gat), .ZN(new_n331_));
  INV_X1    g130(.A(G176gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT23), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(G183gat), .A3(G190gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n331_), .A2(new_n332_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(KEYINPUT24), .A3(new_n340_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n329_), .A2(new_n333_), .A3(new_n338_), .A4(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT85), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n346_), .A2(new_n340_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n347_), .A2(KEYINPUT85), .A3(new_n333_), .A4(new_n329_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n331_), .A2(KEYINPUT22), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT22), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G169gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n352_), .A3(new_n332_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n340_), .A2(KEYINPUT78), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(G169gat), .A3(G176gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n353_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT87), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n334_), .A2(new_n336_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n321_), .A2(new_n325_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT87), .B1(G183gat), .B2(G190gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n361_), .A2(new_n365_), .B1(new_n338_), .B2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n360_), .A2(new_n368_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n349_), .A2(new_n369_), .A3(new_n217_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n346_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n371_), .A2(new_n329_), .A3(new_n333_), .A4(new_n338_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n365_), .A2(new_n353_), .A3(new_n354_), .A4(new_n356_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n217_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT19), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(KEYINPUT20), .A3(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n320_), .B1(new_n370_), .B2(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n360_), .A2(new_n368_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n381_), .A2(new_n218_), .A3(new_n344_), .A4(new_n348_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n374_), .B2(new_n217_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n382_), .A2(KEYINPUT89), .A3(new_n378_), .A4(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n217_), .B1(new_n349_), .B2(new_n369_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n372_), .A2(new_n373_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n383_), .B1(new_n389_), .B2(new_n218_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n387_), .B1(new_n391_), .B2(new_n377_), .ZN(new_n392_));
  AOI211_X1 g191(.A(KEYINPUT88), .B(new_n378_), .C1(new_n388_), .C2(new_n390_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n386_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT91), .ZN(new_n396_));
  XOR2_X1   g195(.A(KEYINPUT90), .B(KEYINPUT18), .Z(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G8gat), .B(G36gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n394_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n400_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n386_), .B(new_n402_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(KEYINPUT92), .A3(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n392_), .A2(new_n393_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT92), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n402_), .A4(new_n386_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n319_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT32), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n400_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n394_), .A2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n313_), .B1(new_n295_), .B2(new_n314_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n306_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n315_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n381_), .A2(new_n218_), .A3(new_n342_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n384_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n377_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n419_), .B1(new_n377_), .B2(new_n391_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n420_), .A2(new_n410_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n411_), .A2(new_n416_), .A3(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n286_), .B1(new_n408_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n281_), .A2(new_n279_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n283_), .A2(new_n284_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n276_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT27), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n404_), .A2(new_n429_), .A3(new_n407_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n420_), .A2(new_n400_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n403_), .A2(new_n431_), .A3(KEYINPUT27), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n428_), .A2(new_n430_), .A3(new_n416_), .A4(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n423_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G71gat), .B(G99gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G43gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n389_), .B(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G227gat), .A2(G233gat), .ZN(new_n438_));
  INV_X1    g237(.A(G15gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT30), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT31), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n437_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT79), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n444_), .A2(new_n291_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n291_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n434_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT97), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n447_), .A2(new_n415_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n430_), .A2(new_n432_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n286_), .A3(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n434_), .A2(KEYINPUT97), .A3(new_n447_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n450_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT70), .B(G8gat), .ZN(new_n456_));
  INV_X1    g255(.A(G1gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT14), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G15gat), .B(G22gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT71), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G1gat), .B(G8gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n460_), .B(KEYINPUT71), .ZN(new_n465_));
  INV_X1    g264(.A(new_n463_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G43gat), .B(G50gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n464_), .A2(new_n467_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n470_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n472_));
  OAI211_X1 g271(.A(G229gat), .B(G233gat), .C1(new_n471_), .C2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n464_), .A2(new_n467_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n470_), .B(KEYINPUT15), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT76), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n464_), .A2(new_n467_), .A3(new_n470_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G229gat), .A2(G233gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT75), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .A4(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n473_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n476_), .A2(new_n478_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n480_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT76), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G113gat), .B(G141gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G169gat), .B(G197gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n486_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n485_), .A2(new_n473_), .A3(new_n481_), .A4(new_n489_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(KEYINPUT77), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT77), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G190gat), .B(G218gat), .Z(new_n499_));
  XNOR2_X1  g298(.A(G134gat), .B(G162gat), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n500_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n501_), .A2(KEYINPUT36), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT36), .B1(new_n501_), .B2(new_n502_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n505_), .B(KEYINPUT68), .Z(new_n506_));
  XOR2_X1   g305(.A(KEYINPUT10), .B(G99gat), .Z(new_n507_));
  INV_X1    g306(.A(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G85gat), .B(G92gat), .Z(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT9), .ZN(new_n511_));
  INV_X1    g310(.A(G85gat), .ZN(new_n512_));
  INV_X1    g311(.A(G92gat), .ZN(new_n513_));
  OR3_X1    g312(.A1(new_n512_), .A2(new_n513_), .A3(KEYINPUT9), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT6), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n509_), .A2(new_n511_), .A3(new_n514_), .A4(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT7), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT6), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n515_), .B(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n510_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT8), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT64), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n523_), .A2(new_n525_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n517_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n475_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT66), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G232gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT34), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT35), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AND4_X1   g336(.A1(new_n514_), .A2(new_n509_), .A3(new_n511_), .A4(new_n516_), .ZN(new_n538_));
  OAI221_X1 g337(.A(new_n510_), .B1(KEYINPUT64), .B2(new_n524_), .C1(new_n520_), .C2(new_n522_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n523_), .A2(new_n525_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n541_), .A2(new_n470_), .B1(new_n535_), .B2(new_n534_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n531_), .A2(new_n537_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n537_), .B1(new_n531_), .B2(new_n542_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n506_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n545_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n504_), .B(KEYINPUT67), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n543_), .A3(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n546_), .A2(new_n549_), .A3(KEYINPUT37), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT69), .B1(new_n544_), .B2(new_n545_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT69), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n547_), .A2(new_n553_), .A3(new_n543_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n554_), .A3(new_n505_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n549_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT37), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n551_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT11), .ZN(new_n560_));
  XOR2_X1   g359(.A(G71gat), .B(G78gat), .Z(new_n561_));
  OR2_X1    g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n559_), .A2(KEYINPUT11), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n561_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT72), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n474_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n569_), .A2(new_n570_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  OR3_X1    g378(.A1(new_n571_), .A2(new_n572_), .A3(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n577_), .A2(new_n578_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT74), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n558_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n541_), .A2(new_n565_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n517_), .B(new_n565_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OAI22_X1  g387(.A1(new_n586_), .A2(new_n588_), .B1(KEYINPUT12), .B2(new_n565_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G230gat), .A2(G233gat), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT65), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n564_), .A2(new_n563_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n528_), .A2(new_n562_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n591_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n594_), .B1(new_n541_), .B2(new_n565_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(KEYINPUT65), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n589_), .B(new_n590_), .C1(new_n595_), .C2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n590_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n599_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G120gat), .B(G148gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT5), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G176gat), .B(G204gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n598_), .A2(new_n600_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n605_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT13), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n585_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n455_), .A2(new_n498_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n455_), .A2(new_n612_), .A3(KEYINPUT98), .A4(new_n498_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n416_), .A2(G1gat), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n455_), .A2(new_n556_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n610_), .A2(new_n493_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(new_n583_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G1gat), .B1(new_n624_), .B2(new_n416_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT100), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n620_), .A2(new_n628_), .A3(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(G1324gat));
  INV_X1    g429(.A(new_n452_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n631_), .A2(new_n456_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n615_), .A2(new_n616_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n455_), .A2(new_n631_), .A3(new_n556_), .A4(new_n623_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(G8gat), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n637_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  AOI211_X1 g439(.A(KEYINPUT102), .B(KEYINPUT39), .C1(new_n636_), .C2(G8gat), .ZN(new_n641_));
  OAI22_X1  g440(.A1(new_n640_), .A2(new_n641_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n635_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT40), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n635_), .A2(KEYINPUT40), .A3(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1325gat));
  OAI21_X1  g446(.A(G15gat), .B1(new_n624_), .B2(new_n447_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT41), .Z(new_n649_));
  AND2_X1   g448(.A1(new_n445_), .A2(new_n446_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n439_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n613_), .B2(new_n651_), .ZN(G1326gat));
  OAI21_X1  g451(.A(G22gat), .B1(new_n624_), .B2(new_n286_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT42), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n286_), .A2(G22gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n613_), .B2(new_n655_), .ZN(G1327gat));
  NOR3_X1   g455(.A1(new_n584_), .A2(new_n611_), .A3(new_n556_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n455_), .A2(new_n657_), .A3(new_n498_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(G29gat), .B1(new_n659_), .B2(new_n415_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n558_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n454_), .A2(new_n453_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT97), .B1(new_n434_), .B2(new_n447_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n661_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT43), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n455_), .A2(new_n666_), .A3(new_n661_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n622_), .A2(new_n584_), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT44), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  INV_X1    g470(.A(new_n669_), .ZN(new_n672_));
  AOI211_X1 g471(.A(new_n671_), .B(new_n672_), .C1(new_n665_), .C2(new_n667_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n670_), .A2(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n415_), .A2(G29gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n660_), .B1(new_n674_), .B2(new_n675_), .ZN(G1328gat));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  INV_X1    g476(.A(G36gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n674_), .B2(new_n631_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n631_), .A2(new_n678_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT103), .Z(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OR3_X1    g482(.A1(new_n658_), .A2(new_n680_), .A3(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n658_), .B2(new_n680_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n677_), .B1(new_n679_), .B2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n664_), .A2(KEYINPUT43), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n666_), .B1(new_n455_), .B2(new_n661_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n669_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n671_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n668_), .A2(KEYINPUT44), .A3(new_n669_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(new_n631_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G36gat), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n694_), .A2(KEYINPUT46), .A3(new_n684_), .A4(new_n685_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n687_), .A2(new_n695_), .ZN(G1329gat));
  NAND4_X1  g495(.A1(new_n691_), .A2(G43gat), .A3(new_n650_), .A4(new_n692_), .ZN(new_n697_));
  INV_X1    g496(.A(G43gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n698_), .B1(new_n658_), .B2(new_n447_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT105), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT47), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n697_), .A2(new_n703_), .A3(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1330gat));
  OR3_X1    g504(.A1(new_n658_), .A2(G50gat), .A3(new_n286_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n674_), .A2(KEYINPUT106), .A3(new_n428_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(G50gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT106), .B1(new_n674_), .B2(new_n428_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n706_), .B1(new_n708_), .B2(new_n709_), .ZN(G1331gat));
  INV_X1    g509(.A(new_n493_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n455_), .A2(new_n711_), .ZN(new_n712_));
  AND4_X1   g511(.A1(new_n611_), .A2(new_n712_), .A3(new_n584_), .A4(new_n558_), .ZN(new_n713_));
  INV_X1    g512(.A(G57gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n415_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n584_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n498_), .A2(new_n716_), .A3(new_n610_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n621_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n621_), .A2(KEYINPUT107), .A3(new_n717_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(new_n415_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n715_), .B1(new_n723_), .B2(new_n714_), .ZN(G1332gat));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n713_), .A2(new_n725_), .A3(new_n631_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n720_), .A2(new_n631_), .A3(new_n721_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(G64gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G64gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(G1333gat));
  INV_X1    g530(.A(G71gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n713_), .A2(new_n732_), .A3(new_n650_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n720_), .A2(new_n650_), .A3(new_n721_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT49), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(G71gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n734_), .B2(G71gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(G1334gat));
  INV_X1    g537(.A(G78gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n713_), .A2(new_n739_), .A3(new_n428_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n720_), .A2(new_n428_), .A3(new_n721_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(G78gat), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n741_), .B2(G78gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1335gat));
  INV_X1    g544(.A(new_n556_), .ZN(new_n746_));
  AND4_X1   g545(.A1(new_n746_), .A2(new_n712_), .A3(new_n611_), .A4(new_n716_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n512_), .A3(new_n415_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n611_), .A2(new_n716_), .A3(new_n711_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT109), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n750_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT110), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(new_n415_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n748_), .B1(new_n753_), .B2(new_n512_), .ZN(G1336gat));
  NAND3_X1  g553(.A1(new_n747_), .A2(new_n513_), .A3(new_n631_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n752_), .A2(new_n631_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(new_n513_), .ZN(G1337gat));
  AND2_X1   g556(.A1(new_n650_), .A2(new_n507_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n668_), .A2(new_n650_), .A3(new_n750_), .ZN(new_n759_));
  AOI22_X1  g558(.A1(new_n747_), .A2(new_n758_), .B1(new_n759_), .B2(G99gat), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g560(.A1(new_n747_), .A2(new_n508_), .A3(new_n428_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n668_), .A2(new_n428_), .A3(new_n750_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(G106gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G106gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT53), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n769_), .B(new_n762_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1339gat));
  NAND4_X1  g570(.A1(new_n558_), .A2(new_n497_), .A3(new_n610_), .A4(new_n584_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n775_), .A2(KEYINPUT56), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n778_));
  XOR2_X1   g577(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n779_));
  NAND3_X1  g578(.A1(new_n598_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n589_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n599_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n593_), .A2(new_n591_), .A3(new_n594_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n596_), .A2(KEYINPUT65), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n786_), .A2(KEYINPUT55), .A3(new_n590_), .A4(new_n589_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n783_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n778_), .B1(new_n598_), .B2(new_n779_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n781_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n777_), .B1(new_n790_), .B2(new_n605_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n598_), .A2(new_n779_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT112), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n793_), .A2(new_n780_), .A3(new_n787_), .A4(new_n783_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(new_n604_), .A3(new_n776_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n489_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n796_));
  AND4_X1   g595(.A1(new_n485_), .A2(new_n473_), .A3(new_n481_), .A4(new_n489_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n606_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n791_), .A2(new_n795_), .A3(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n480_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n490_), .C1(new_n483_), .C2(new_n480_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n492_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT114), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n492_), .A2(new_n805_), .A3(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n609_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n746_), .B1(new_n800_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT115), .B1(new_n809_), .B2(KEYINPUT57), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n794_), .A2(new_n604_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n798_), .B1(new_n813_), .B2(new_n777_), .ZN(new_n814_));
  AOI22_X1  g613(.A1(new_n814_), .A2(new_n795_), .B1(new_n609_), .B2(new_n807_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n811_), .B(new_n812_), .C1(new_n815_), .C2(new_n746_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n809_), .A2(KEYINPUT57), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n813_), .A2(KEYINPUT56), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n607_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n794_), .A2(new_n820_), .A3(new_n604_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n819_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n818_), .A2(new_n819_), .A3(KEYINPUT58), .A4(new_n821_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n661_), .A3(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n810_), .A2(new_n816_), .A3(new_n817_), .A4(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n774_), .B1(new_n827_), .B2(new_n583_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n650_), .A2(new_n452_), .A3(new_n415_), .A4(new_n286_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT116), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT59), .B1(new_n828_), .B2(new_n831_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n558_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n834_), .A2(new_n825_), .B1(new_n809_), .B2(KEYINPUT57), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n812_), .B1(new_n815_), .B2(new_n746_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n584_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n830_), .B(new_n833_), .C1(new_n837_), .C2(new_n774_), .ZN(new_n838_));
  XOR2_X1   g637(.A(KEYINPUT118), .B(G113gat), .Z(new_n839_));
  NAND2_X1  g638(.A1(new_n498_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n832_), .A2(new_n838_), .A3(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n828_), .A2(new_n831_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G113gat), .B1(new_n843_), .B2(new_n493_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT119), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(G113gat), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n827_), .A2(new_n583_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n774_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n830_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n846_), .B1(new_n850_), .B2(new_n711_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n832_), .A2(new_n838_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n851_), .B(new_n852_), .C1(new_n853_), .C2(new_n840_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n845_), .A2(new_n854_), .ZN(G1340gat));
  OAI21_X1  g654(.A(G120gat), .B1(new_n853_), .B2(new_n610_), .ZN(new_n856_));
  INV_X1    g655(.A(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n610_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(KEYINPUT60), .B2(new_n857_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n850_), .B2(new_n859_), .ZN(G1341gat));
  AOI21_X1  g659(.A(G127gat), .B1(new_n843_), .B2(new_n584_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n853_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT120), .B(G127gat), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n583_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n861_), .B1(new_n862_), .B2(new_n864_), .ZN(G1342gat));
  AOI21_X1  g664(.A(G134gat), .B1(new_n843_), .B2(new_n746_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n661_), .A2(G134gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT121), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n862_), .B2(new_n868_), .ZN(G1343gat));
  NOR4_X1   g668(.A1(new_n631_), .A2(new_n416_), .A3(new_n650_), .A4(new_n286_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n849_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n493_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g673(.A1(new_n871_), .A2(new_n610_), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT122), .B(G148gat), .Z(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1345gat));
  NOR2_X1   g676(.A1(new_n871_), .A2(new_n716_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT61), .B(G155gat), .Z(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  OAI21_X1  g679(.A(G162gat), .B1(new_n871_), .B2(new_n558_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n746_), .A2(new_n220_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n871_), .B2(new_n882_), .ZN(G1347gat));
  NAND2_X1  g682(.A1(new_n451_), .A2(new_n631_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n428_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n837_), .B2(new_n774_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n887_), .A2(new_n350_), .A3(new_n352_), .A4(new_n493_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n884_), .A2(new_n711_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(KEYINPUT123), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n889_), .A2(KEYINPUT123), .ZN(new_n891_));
  OAI221_X1 g690(.A(new_n286_), .B1(new_n890_), .B2(new_n891_), .C1(new_n837_), .C2(new_n774_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n331_), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n892_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n893_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n888_), .B1(new_n896_), .B2(new_n897_), .ZN(G1348gat));
  NOR2_X1   g697(.A1(new_n828_), .A2(new_n428_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n884_), .A2(new_n610_), .A3(new_n332_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n332_), .B1(new_n886_), .B2(new_n610_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT125), .ZN(G1349gat));
  NAND4_X1  g703(.A1(new_n899_), .A2(new_n631_), .A3(new_n451_), .A4(new_n584_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n583_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n905_), .A2(new_n321_), .B1(new_n887_), .B2(new_n906_), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n886_), .B2(new_n558_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n746_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n909_));
  XOR2_X1   g708(.A(new_n909_), .B(KEYINPUT126), .Z(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n886_), .B2(new_n910_), .ZN(G1351gat));
  NAND4_X1  g710(.A1(new_n631_), .A2(new_n416_), .A3(new_n447_), .A4(new_n428_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n828_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n493_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n611_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g716(.A(new_n583_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT127), .Z(new_n919_));
  NAND2_X1  g718(.A1(new_n913_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n920_), .B(new_n921_), .Z(G1354gat));
  INV_X1    g721(.A(G218gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n913_), .A2(new_n923_), .A3(new_n746_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n828_), .A2(new_n558_), .A3(new_n912_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n923_), .ZN(G1355gat));
endmodule


