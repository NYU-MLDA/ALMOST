//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n960_, new_n961_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n972_, new_n973_,
    new_n974_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_, new_n985_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT64), .Z(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G92gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n207_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  AND3_X1   g012(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT67), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n220_));
  NAND3_X1  g019(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT10), .B(G99gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(G106gat), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n216_), .B(new_n222_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n213_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NOR3_X1   g027(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n219_), .A2(KEYINPUT68), .A3(new_n221_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT68), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n230_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G85gat), .B(G92gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT8), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n230_), .A2(new_n216_), .A3(new_n222_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n235_), .A2(KEYINPUT8), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n226_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G57gat), .B(G64gat), .ZN(new_n243_));
  INV_X1    g042(.A(G78gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G71gat), .ZN(new_n245_));
  INV_X1    g044(.A(G71gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G78gat), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n243_), .A2(KEYINPUT11), .A3(new_n245_), .A4(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G64gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G57gat), .ZN(new_n250_));
  INV_X1    g049(.A(G57gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G64gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n252_), .A3(KEYINPUT11), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n245_), .A2(new_n247_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n243_), .A2(KEYINPUT11), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n248_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(KEYINPUT69), .B(new_n248_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n204_), .B1(new_n242_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G92gat), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n212_), .ZN(new_n265_));
  OAI22_X1  g064(.A1(new_n264_), .A2(new_n265_), .B1(new_n206_), .B2(new_n205_), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n223_), .A2(new_n224_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n266_), .A2(new_n267_), .A3(new_n216_), .A4(new_n222_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n239_), .A2(new_n240_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT8), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n268_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT12), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n259_), .A2(new_n260_), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n257_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n273_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n262_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT70), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n242_), .A2(new_n261_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n272_), .A2(new_n274_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n204_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n283_), .B(new_n262_), .C1(new_n275_), .C2(new_n277_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n279_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G120gat), .B(G148gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT5), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G176gat), .B(G204gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n287_), .B(new_n288_), .Z(new_n289_));
  NAND2_X1  g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n289_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n279_), .A2(new_n282_), .A3(new_n284_), .A4(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT13), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n290_), .A2(KEYINPUT13), .A3(new_n292_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT71), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n296_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n298_), .A2(new_n301_), .A3(KEYINPUT72), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT15), .ZN(new_n307_));
  XOR2_X1   g106(.A(G29gat), .B(G36gat), .Z(new_n308_));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G29gat), .B(G36gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT73), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G43gat), .B(G50gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n313_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n307_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n316_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(KEYINPUT15), .A3(new_n314_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n272_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G232gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT34), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT35), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT68), .B1(new_n219_), .B2(new_n221_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT7), .ZN(new_n327_));
  INV_X1    g126(.A(G99gat), .ZN(new_n328_));
  INV_X1    g127(.A(G106gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n227_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n326_), .A2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n235_), .B1(new_n332_), .B2(new_n231_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n241_), .B1(new_n333_), .B2(new_n270_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n318_), .A2(new_n314_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n268_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n320_), .A2(new_n325_), .A3(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n323_), .A2(new_n324_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n338_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n320_), .A2(new_n340_), .A3(new_n325_), .A4(new_n336_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G190gat), .B(G218gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G134gat), .B(G162gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT36), .Z(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n345_), .A2(KEYINPUT36), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n339_), .A2(new_n341_), .A3(new_n348_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n347_), .A2(KEYINPUT37), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT74), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n342_), .A2(KEYINPUT74), .A3(new_n346_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(new_n353_), .A3(new_n349_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT37), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n350_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G1gat), .B(G8gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT75), .ZN(new_n359_));
  INV_X1    g158(.A(G15gat), .ZN(new_n360_));
  INV_X1    g159(.A(G22gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G15gat), .A2(G22gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G1gat), .A2(G8gat), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n362_), .A2(new_n363_), .B1(KEYINPUT14), .B2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n359_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT76), .ZN(new_n367_));
  AND2_X1   g166(.A1(G231gat), .A2(G233gat), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n367_), .A2(new_n368_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n257_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n367_), .A2(new_n368_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n368_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n276_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G127gat), .B(G155gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT16), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G183gat), .B(G211gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT17), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n371_), .A2(new_n374_), .A3(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n274_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n372_), .A2(new_n373_), .A3(new_n261_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n378_), .B(KEYINPUT17), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n381_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n357_), .A2(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n306_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G197gat), .B(G204gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT88), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G211gat), .B(G218gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT21), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n389_), .B(KEYINPUT21), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n392_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT87), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT87), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n396_), .A2(new_n399_), .A3(new_n392_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n395_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(G169gat), .A2(G176gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G169gat), .A2(G176gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT24), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n404_), .B2(KEYINPUT91), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(KEYINPUT91), .B2(new_n404_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G183gat), .A2(G190gat), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n407_), .A2(KEYINPUT23), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(KEYINPUT23), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT24), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n408_), .A2(new_n409_), .B1(new_n410_), .B2(new_n402_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT26), .B(G190gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT25), .B(G183gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n406_), .A2(new_n411_), .A3(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n407_), .B(KEYINPUT23), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(G183gat), .B2(G190gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n403_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT22), .B(G169gat), .ZN(new_n419_));
  INV_X1    g218(.A(G176gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n415_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n401_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n395_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n396_), .A2(new_n399_), .A3(new_n392_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n399_), .B1(new_n396_), .B2(new_n392_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n404_), .A2(new_n402_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT78), .ZN(new_n430_));
  XOR2_X1   g229(.A(KEYINPUT77), .B(G183gat), .Z(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT25), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT25), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(G183gat), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n430_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT77), .B(G183gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n436_), .A2(new_n433_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n412_), .B1(new_n437_), .B2(KEYINPUT78), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n411_), .B(new_n429_), .C1(new_n435_), .C2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n416_), .B1(G190gat), .B2(new_n436_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n421_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n428_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n424_), .A2(new_n443_), .A3(KEYINPUT20), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G226gat), .A2(G233gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT19), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n439_), .A2(new_n441_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n401_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n446_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n415_), .A2(new_n422_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n428_), .A2(new_n451_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n449_), .A2(KEYINPUT20), .A3(new_n450_), .A4(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n447_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G64gat), .B(G92gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT94), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT95), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n456_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G8gat), .B(G36gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n454_), .A2(KEYINPUT32), .A3(new_n461_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n461_), .A2(KEYINPUT32), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT20), .B1(new_n428_), .B2(new_n442_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n401_), .A2(new_n423_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n446_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT92), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(KEYINPUT92), .B(new_n446_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n424_), .A2(new_n443_), .A3(KEYINPUT20), .A4(new_n450_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G1gat), .B(G29gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT99), .B(G85gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT0), .B(G57gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  XNOR2_X1  g275(.A(G127gat), .B(G134gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G113gat), .B(G120gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G141gat), .A2(G148gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT83), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G155gat), .A2(G162gat), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n483_), .A2(KEYINPUT1), .ZN(new_n484_));
  NOR2_X1   g283(.A1(G155gat), .A2(G162gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(KEYINPUT1), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(G141gat), .ZN(new_n489_));
  INV_X1    g288(.A(G148gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n482_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n480_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n493_), .A2(KEYINPUT2), .B1(new_n491_), .B2(KEYINPUT3), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n491_), .A2(KEYINPUT3), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n494_), .B(new_n495_), .C1(new_n481_), .C2(KEYINPUT2), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n486_), .A2(new_n483_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n497_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n479_), .B(new_n492_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G225gat), .A2(G233gat), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n479_), .A2(KEYINPUT81), .ZN(new_n504_));
  INV_X1    g303(.A(new_n477_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n478_), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT81), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n492_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n496_), .A2(new_n498_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT84), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n510_), .B1(new_n512_), .B2(new_n499_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n502_), .B(new_n503_), .C1(new_n509_), .C2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT100), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n492_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n508_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT100), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n503_), .A4(new_n502_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(KEYINPUT98), .B(KEYINPUT4), .Z(new_n521_));
  NOR2_X1   g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n502_), .B(KEYINPUT4), .C1(new_n509_), .C2(new_n513_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT96), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n517_), .A2(KEYINPUT96), .A3(KEYINPUT4), .A4(new_n502_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n522_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n503_), .B(KEYINPUT97), .ZN(new_n528_));
  AOI211_X1 g327(.A(new_n476_), .B(new_n520_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n476_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n525_), .A2(new_n526_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n522_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n528_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n520_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n530_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  OAI221_X1 g334(.A(new_n462_), .B1(new_n463_), .B2(new_n471_), .C1(new_n529_), .C2(new_n535_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n533_), .A2(KEYINPUT33), .A3(new_n530_), .A4(new_n534_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT101), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n520_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n540_), .A2(KEYINPUT101), .A3(KEYINPUT33), .A4(new_n530_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n517_), .A2(new_n528_), .A3(new_n502_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n544_), .A2(new_n476_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n527_), .A2(KEYINPUT102), .A3(new_n503_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT102), .B1(new_n527_), .B2(new_n503_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n545_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n540_), .A2(new_n530_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT33), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n461_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n471_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n468_), .A2(new_n461_), .A3(new_n469_), .A4(new_n470_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n549_), .A2(new_n552_), .A3(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n536_), .B1(new_n543_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G227gat), .A2(G233gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n560_), .B(KEYINPUT80), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT30), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT31), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G15gat), .B(G43gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT79), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(G71gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(G99gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n566_), .B(new_n246_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n328_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n448_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n568_), .A2(new_n570_), .A3(new_n442_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n509_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n509_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n564_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n572_), .A2(new_n573_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n508_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(new_n563_), .A3(new_n574_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n577_), .A2(new_n580_), .A3(KEYINPUT82), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT82), .B1(new_n577_), .B2(new_n580_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G22gat), .B(G50gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT86), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n585_), .B1(new_n516_), .B2(KEYINPUT29), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT29), .ZN(new_n588_));
  INV_X1    g387(.A(new_n585_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n513_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n586_), .A2(new_n587_), .A3(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n587_), .B1(new_n586_), .B2(new_n590_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n428_), .B1(new_n513_), .B2(new_n588_), .ZN(new_n594_));
  INV_X1    g393(.A(G228gat), .ZN(new_n595_));
  INV_X1    g394(.A(G233gat), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  OAI221_X1 g397(.A(new_n428_), .B1(new_n595_), .B2(new_n596_), .C1(new_n513_), .C2(new_n588_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G78gat), .B(G106gat), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n598_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n593_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT89), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT89), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n593_), .B(new_n606_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n598_), .A2(new_n599_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n600_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n610_), .B1(new_n602_), .B2(KEYINPUT90), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT90), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n609_), .A2(new_n612_), .A3(new_n600_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n593_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n583_), .A2(new_n608_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n583_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n577_), .A2(new_n580_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n615_), .A2(new_n605_), .A3(new_n620_), .A4(new_n607_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT27), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n454_), .B2(new_n553_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n555_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT103), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT103), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n555_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n529_), .A2(new_n535_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n556_), .A2(new_n623_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n629_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n559_), .A2(new_n617_), .B1(new_n622_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT75), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n358_), .B(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(new_n365_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n314_), .A3(new_n318_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n366_), .A2(new_n335_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n637_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n366_), .B2(new_n335_), .ZN(new_n644_));
  AOI22_X1  g443(.A1(new_n640_), .A2(new_n642_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G113gat), .B(G141gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G169gat), .B(G197gat), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n646_), .B(new_n647_), .Z(new_n648_));
  XNOR2_X1  g447(.A(new_n645_), .B(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n634_), .A2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n388_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(G1gat), .ZN(new_n653_));
  INV_X1    g452(.A(new_n535_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n550_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n652_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT38), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n354_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n559_), .A2(new_n617_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n622_), .A2(new_n633_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n659_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n302_), .A2(new_n650_), .A3(new_n386_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G1gat), .B1(new_n664_), .B2(new_n630_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n656_), .A2(new_n657_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n658_), .A2(new_n665_), .A3(new_n666_), .ZN(G1324gat));
  AND2_X1   g466(.A1(new_n629_), .A2(new_n631_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G8gat), .B1(new_n664_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT39), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n668_), .A2(G8gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n388_), .A2(new_n651_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n388_), .A2(KEYINPUT104), .A3(new_n651_), .A4(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n670_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n670_), .B2(new_n676_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1325gat));
  OAI21_X1  g479(.A(G15gat), .B1(new_n664_), .B2(new_n583_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT41), .Z(new_n682_));
  INV_X1    g481(.A(new_n583_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n652_), .A2(new_n360_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1326gat));
  INV_X1    g484(.A(new_n618_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G22gat), .B1(new_n664_), .B2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n652_), .A2(new_n361_), .A3(new_n618_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1327gat));
  INV_X1    g490(.A(new_n386_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n302_), .A2(new_n692_), .A3(new_n354_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n651_), .A2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G29gat), .B1(new_n694_), .B2(new_n655_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n298_), .A2(new_n649_), .A3(new_n301_), .A4(new_n386_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT43), .B1(new_n634_), .B2(new_n356_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n542_), .A2(new_n552_), .A3(new_n549_), .A4(new_n557_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n616_), .B1(new_n699_), .B2(new_n536_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n632_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n698_), .B(new_n357_), .C1(new_n700_), .C2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n696_), .B1(new_n697_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT44), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n704_), .A2(G29gat), .A3(new_n655_), .ZN(new_n705_));
  XOR2_X1   g504(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n706_));
  OR2_X1    g505(.A1(new_n703_), .A2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n695_), .B1(new_n705_), .B2(new_n707_), .ZN(G1328gat));
  AOI21_X1  g507(.A(new_n668_), .B1(new_n703_), .B2(KEYINPUT44), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G36gat), .ZN(new_n711_));
  INV_X1    g510(.A(G36gat), .ZN(new_n712_));
  INV_X1    g511(.A(new_n668_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n651_), .A2(new_n712_), .A3(new_n713_), .A4(new_n693_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT45), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n711_), .A2(KEYINPUT46), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n712_), .B1(new_n707_), .B2(new_n709_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n715_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n716_), .A2(new_n720_), .ZN(G1329gat));
  NAND2_X1  g520(.A1(new_n694_), .A2(new_n683_), .ZN(new_n722_));
  XOR2_X1   g521(.A(KEYINPUT108), .B(G43gat), .Z(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n704_), .A2(G43gat), .A3(new_n620_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n703_), .A2(new_n706_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n724_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT47), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n729_), .B(new_n724_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1330gat));
  INV_X1    g530(.A(G50gat), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n618_), .A2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT110), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n694_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n686_), .B1(new_n703_), .B2(KEYINPUT44), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n707_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n738_), .B2(G50gat), .ZN(new_n739_));
  AOI211_X1 g538(.A(KEYINPUT109), .B(new_n732_), .C1(new_n707_), .C2(new_n737_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n735_), .B1(new_n739_), .B2(new_n740_), .ZN(G1331gat));
  INV_X1    g540(.A(new_n305_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT72), .B1(new_n298_), .B2(new_n301_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n386_), .A2(new_n649_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n662_), .A2(new_n744_), .A3(new_n745_), .A4(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n304_), .A2(new_n305_), .A3(new_n746_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n354_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT111), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G57gat), .B1(new_n751_), .B2(new_n630_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n634_), .A2(new_n649_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n753_), .A2(new_n302_), .A3(new_n387_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n251_), .A3(new_n655_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(G1332gat));
  NAND3_X1  g555(.A1(new_n754_), .A2(new_n249_), .A3(new_n713_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n747_), .A2(new_n750_), .A3(new_n713_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT48), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(G64gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G64gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT112), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n764_), .B(new_n757_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1333gat));
  NAND3_X1  g565(.A1(new_n754_), .A2(new_n246_), .A3(new_n683_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT49), .ZN(new_n768_));
  INV_X1    g567(.A(new_n751_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n683_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n768_), .B1(new_n770_), .B2(G71gat), .ZN(new_n771_));
  AOI211_X1 g570(.A(KEYINPUT49), .B(new_n246_), .C1(new_n769_), .C2(new_n683_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n767_), .B1(new_n771_), .B2(new_n772_), .ZN(G1334gat));
  NAND3_X1  g572(.A1(new_n754_), .A2(new_n244_), .A3(new_n618_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n769_), .A2(new_n618_), .ZN(new_n775_));
  XOR2_X1   g574(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n776_));
  AND3_X1   g575(.A1(new_n775_), .A2(G78gat), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n775_), .B2(G78gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(G1335gat));
  NOR2_X1   g578(.A1(new_n692_), .A2(new_n354_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n753_), .A2(new_n744_), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(G85gat), .B1(new_n782_), .B2(new_n655_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n692_), .A2(new_n649_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n302_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT114), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n302_), .A2(new_n787_), .A3(new_n784_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n697_), .A2(new_n702_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n630_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n783_), .B1(new_n791_), .B2(new_n792_), .ZN(G1336gat));
  NAND3_X1  g592(.A1(new_n782_), .A2(new_n263_), .A3(new_n713_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n791_), .A2(new_n713_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n263_), .ZN(G1337gat));
  INV_X1    g595(.A(new_n620_), .ZN(new_n797_));
  OR3_X1    g596(.A1(new_n781_), .A2(new_n797_), .A3(new_n223_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n789_), .A2(new_n683_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n328_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g600(.A1(new_n781_), .A2(new_n686_), .A3(new_n224_), .ZN(new_n802_));
  AOI211_X1 g601(.A(KEYINPUT52), .B(new_n329_), .C1(new_n789_), .C2(new_n618_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n697_), .A2(new_n702_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n786_), .A2(new_n788_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n618_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n804_), .B1(new_n807_), .B2(G106gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n802_), .B1(new_n803_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT53), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(new_n802_), .C1(new_n803_), .C2(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1339gat));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n356_), .A2(new_n746_), .A3(new_n296_), .A4(new_n295_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n815_), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT116), .B1(new_n815_), .B2(KEYINPUT54), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n815_), .A2(KEYINPUT54), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n816_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT12), .B1(new_n242_), .B2(new_n257_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n281_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  OAI22_X1  g623(.A1(new_n821_), .A2(new_n278_), .B1(new_n824_), .B2(new_n203_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n284_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n257_), .B1(new_n334_), .B2(new_n268_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n823_), .B1(new_n827_), .B2(new_n273_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n283_), .B1(new_n828_), .B2(new_n262_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n826_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n825_), .B1(new_n830_), .B2(new_n821_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n820_), .B(KEYINPUT56), .C1(new_n831_), .C2(new_n291_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n279_), .A2(new_n821_), .A3(new_n284_), .ZN(new_n834_));
  OAI22_X1  g633(.A1(new_n275_), .A2(new_n277_), .B1(new_n274_), .B2(new_n272_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n203_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n204_), .A2(new_n835_), .B1(new_n837_), .B2(KEYINPUT55), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n291_), .B1(new_n834_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n833_), .B1(new_n839_), .B2(KEYINPUT117), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n649_), .A2(new_n292_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n832_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n648_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n643_), .A2(new_n639_), .A3(new_n642_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n645_), .A2(new_n648_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n293_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT57), .B1(new_n847_), .B2(new_n354_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n659_), .B1(new_n842_), .B2(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT57), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n292_), .A2(new_n845_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n839_), .B2(new_n833_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT56), .B1(new_n831_), .B2(new_n291_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n356_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n853_), .A2(new_n854_), .A3(KEYINPUT58), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT118), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n853_), .A2(new_n854_), .A3(new_n860_), .A4(KEYINPUT58), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n859_), .A3(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n849_), .A2(new_n851_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n819_), .B1(new_n863_), .B2(new_n386_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n713_), .A2(new_n630_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n621_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n864_), .A2(new_n868_), .A3(new_n650_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n814_), .B1(new_n869_), .B2(G113gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT59), .B1(new_n864_), .B2(new_n868_), .ZN(new_n871_));
  INV_X1    g670(.A(G113gat), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n650_), .A2(new_n872_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n857_), .A2(new_n861_), .A3(new_n859_), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT121), .B1(new_n874_), .B2(new_n848_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n862_), .B(new_n876_), .C1(KEYINPUT57), .C2(new_n850_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(new_n851_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n819_), .B1(new_n878_), .B2(new_n386_), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n880_));
  NAND2_X1  g679(.A1(new_n867_), .A2(new_n880_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n871_), .B(new_n873_), .C1(new_n879_), .C2(new_n881_), .ZN(new_n882_));
  OR3_X1    g681(.A1(new_n816_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884_));
  AOI211_X1 g683(.A(new_n884_), .B(new_n659_), .C1(new_n842_), .C2(new_n846_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n874_), .A2(new_n848_), .A3(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n883_), .B1(new_n886_), .B2(new_n692_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n867_), .ZN(new_n888_));
  OAI211_X1 g687(.A(KEYINPUT119), .B(new_n872_), .C1(new_n888_), .C2(new_n650_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n870_), .A2(new_n882_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT122), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n870_), .A2(new_n882_), .A3(new_n892_), .A4(new_n889_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1340gat));
  INV_X1    g693(.A(G120gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n306_), .B1(new_n888_), .B2(KEYINPUT59), .ZN(new_n896_));
  INV_X1    g695(.A(new_n881_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n862_), .B1(KEYINPUT57), .B2(new_n850_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n885_), .B1(new_n898_), .B2(KEYINPUT121), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n692_), .B1(new_n899_), .B2(new_n877_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n897_), .B1(new_n900_), .B2(new_n819_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n895_), .B1(new_n896_), .B2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n895_), .A2(KEYINPUT60), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n904_));
  AOI21_X1  g703(.A(G120gat), .B1(new_n302_), .B2(new_n904_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n888_), .A2(new_n903_), .A3(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT123), .B1(new_n902_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n871_), .A2(new_n744_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n879_), .A2(new_n881_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G120gat), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911_));
  INV_X1    g710(.A(new_n906_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n907_), .A2(new_n913_), .ZN(G1341gat));
  NAND3_X1  g713(.A1(new_n901_), .A2(new_n692_), .A3(new_n871_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(G127gat), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n386_), .A2(G127gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n888_), .B2(new_n917_), .ZN(G1342gat));
  NAND3_X1  g717(.A1(new_n901_), .A2(new_n357_), .A3(new_n871_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(G134gat), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n354_), .A2(G134gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n888_), .B2(new_n921_), .ZN(G1343gat));
  NOR2_X1   g721(.A1(new_n864_), .A2(new_n619_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n865_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n650_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n489_), .ZN(G1344gat));
  NOR2_X1   g725(.A1(new_n924_), .A2(new_n306_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(new_n490_), .ZN(G1345gat));
  INV_X1    g727(.A(new_n619_), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n887_), .A2(new_n929_), .A3(new_n692_), .A4(new_n865_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n930_), .A2(KEYINPUT124), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(KEYINPUT124), .ZN(new_n932_));
  XNOR2_X1  g731(.A(KEYINPUT61), .B(G155gat), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  OR3_X1    g733(.A1(new_n931_), .A2(new_n932_), .A3(new_n934_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1346gat));
  OR3_X1    g736(.A1(new_n924_), .A2(G162gat), .A3(new_n354_), .ZN(new_n938_));
  OAI21_X1  g737(.A(G162gat), .B1(new_n924_), .B2(new_n356_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1347gat));
  NOR3_X1   g739(.A1(new_n668_), .A2(new_n655_), .A3(new_n583_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n686_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  OAI211_X1 g742(.A(new_n649_), .B(new_n943_), .C1(new_n900_), .C2(new_n819_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n945_));
  AND3_X1   g744(.A1(new_n944_), .A2(new_n945_), .A3(G169gat), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n944_), .B2(G169gat), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n943_), .B1(new_n900_), .B2(new_n819_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n649_), .A2(new_n419_), .ZN(new_n949_));
  XOR2_X1   g748(.A(new_n949_), .B(KEYINPUT125), .Z(new_n950_));
  OAI22_X1  g749(.A1(new_n946_), .A2(new_n947_), .B1(new_n948_), .B2(new_n950_), .ZN(G1348gat));
  NOR2_X1   g750(.A1(new_n879_), .A2(new_n942_), .ZN(new_n952_));
  AOI21_X1  g751(.A(G176gat), .B1(new_n952_), .B2(new_n302_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n954_), .B1(new_n864_), .B2(new_n618_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n887_), .A2(KEYINPUT126), .A3(new_n686_), .ZN(new_n956_));
  AND3_X1   g755(.A1(new_n955_), .A2(new_n956_), .A3(new_n941_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n306_), .A2(new_n420_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n953_), .B1(new_n957_), .B2(new_n958_), .ZN(G1349gat));
  NOR3_X1   g758(.A1(new_n948_), .A2(new_n413_), .A3(new_n386_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n957_), .A2(new_n692_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n960_), .B1(new_n961_), .B2(new_n431_), .ZN(G1350gat));
  INV_X1    g761(.A(G190gat), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n963_), .B1(new_n952_), .B2(new_n357_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n659_), .A2(new_n412_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n948_), .A2(new_n965_), .ZN(new_n966_));
  OAI21_X1  g765(.A(KEYINPUT127), .B1(new_n964_), .B2(new_n966_), .ZN(new_n967_));
  OAI21_X1  g766(.A(G190gat), .B1(new_n948_), .B2(new_n356_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969_));
  OAI211_X1 g768(.A(new_n968_), .B(new_n969_), .C1(new_n948_), .C2(new_n965_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n967_), .A2(new_n970_), .ZN(G1351gat));
  NOR2_X1   g770(.A1(new_n668_), .A2(new_n655_), .ZN(new_n972_));
  AND2_X1   g771(.A1(new_n923_), .A2(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n973_), .A2(new_n649_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g774(.A1(new_n973_), .A2(new_n744_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g776(.A1(new_n923_), .A2(new_n692_), .A3(new_n972_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n979_));
  AND2_X1   g778(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n980_));
  NOR3_X1   g779(.A1(new_n978_), .A2(new_n979_), .A3(new_n980_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n981_), .B1(new_n978_), .B2(new_n979_), .ZN(G1354gat));
  INV_X1    g781(.A(G218gat), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n973_), .A2(new_n983_), .A3(new_n659_), .ZN(new_n984_));
  AND2_X1   g783(.A1(new_n973_), .A2(new_n357_), .ZN(new_n985_));
  OAI21_X1  g784(.A(new_n984_), .B1(new_n985_), .B2(new_n983_), .ZN(G1355gat));
endmodule


