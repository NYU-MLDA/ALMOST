//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_;
  INV_X1    g000(.A(G228gat), .ZN(new_n202_));
  INV_X1    g001(.A(G233gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT91), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT2), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n206_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT90), .ZN(new_n211_));
  OAI22_X1  g010(.A1(new_n211_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT90), .A3(new_n214_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n208_), .A2(new_n210_), .A3(new_n212_), .A4(new_n215_), .ZN(new_n216_));
  OR3_X1    g015(.A1(KEYINPUT89), .A2(G155gat), .A3(G162gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT89), .B1(G155gat), .B2(G162gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(KEYINPUT1), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G155gat), .A3(G162gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n217_), .A2(new_n218_), .A3(new_n222_), .A4(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n213_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n226_), .A2(new_n205_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n221_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT28), .B1(new_n229_), .B2(KEYINPUT29), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n216_), .A2(new_n220_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT28), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT29), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT92), .ZN(new_n236_));
  INV_X1    g035(.A(G204gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n236_), .B1(new_n237_), .B2(G197gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(G197gat), .ZN(new_n239_));
  INV_X1    g038(.A(G197gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n238_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT93), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT93), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n238_), .A2(new_n241_), .A3(new_n244_), .A4(new_n239_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G211gat), .B(G218gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT21), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n243_), .A2(new_n245_), .A3(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n237_), .A2(G197gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n240_), .A2(G204gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT21), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n252_), .B(new_n246_), .C1(new_n242_), .C2(KEYINPUT21), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n233_), .B2(new_n231_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n235_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G22gat), .B(G50gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n230_), .A3(new_n234_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n258_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n204_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT94), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT95), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n257_), .A2(new_n259_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n258_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n204_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(new_n260_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n263_), .A2(new_n266_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n266_), .B1(new_n263_), .B2(new_n271_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G127gat), .B(G134gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G113gat), .B(G120gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT88), .B(KEYINPUT31), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G227gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(G15gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(KEYINPUT86), .B(G43gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G71gat), .B(G99gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  AND3_X1   g085(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G169gat), .ZN(new_n292_));
  INV_X1    g091(.A(G176gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT22), .B1(new_n292_), .B2(KEYINPUT85), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT22), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G169gat), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n296_), .B(new_n293_), .C1(KEYINPUT85), .C2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n291_), .A2(new_n295_), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302_));
  NOR3_X1   g101(.A1(new_n294_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT25), .B(G183gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT26), .B(G190gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT83), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n307_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n304_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n302_), .A2(new_n301_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n289_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT84), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT84), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n289_), .A2(new_n315_), .A3(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n300_), .B1(new_n311_), .B2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT30), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT87), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n320_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n286_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n286_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n280_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n277_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n229_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n231_), .A2(new_n277_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(KEYINPUT4), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT4), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n229_), .A2(new_n333_), .A3(new_n327_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n330_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n328_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G1gat), .B(G29gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G85gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT0), .B(G57gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n221_), .A2(new_n277_), .A3(new_n228_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n277_), .B1(new_n221_), .B2(new_n228_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n344_), .A2(new_n345_), .A3(new_n333_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n334_), .A2(new_n332_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n336_), .B(new_n341_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n319_), .B(KEYINPUT87), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n324_), .B(new_n279_), .C1(new_n351_), .C2(new_n286_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n326_), .A2(new_n350_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT27), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT20), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n291_), .A2(new_n295_), .A3(new_n299_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n305_), .A2(new_n306_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT83), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n303_), .B1(new_n358_), .B2(new_n308_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n289_), .A2(new_n315_), .A3(new_n312_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n315_), .B1(new_n289_), .B2(new_n312_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n356_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n249_), .A2(new_n253_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT99), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT99), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n318_), .A2(new_n366_), .A3(new_n254_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n355_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n304_), .A2(new_n357_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n373_), .A2(new_n313_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n292_), .A2(KEYINPUT22), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n298_), .A3(new_n293_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n376_), .A2(KEYINPUT97), .A3(new_n295_), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT97), .B1(new_n376_), .B2(new_n295_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n291_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT98), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  OAI211_X1 g180(.A(KEYINPUT98), .B(new_n291_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n374_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n372_), .B1(new_n383_), .B2(new_n364_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n368_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n355_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n386_), .B1(new_n383_), .B2(new_n364_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n372_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n385_), .A2(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(G8gat), .B(G36gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT18), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n385_), .A2(new_n388_), .A3(new_n393_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n396_), .A2(KEYINPUT27), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n364_), .B(new_n379_), .C1(new_n313_), .C2(new_n373_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n371_), .B1(new_n368_), .B2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n386_), .B(new_n371_), .C1(new_n383_), .C2(new_n364_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n394_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n354_), .A2(new_n397_), .B1(new_n398_), .B2(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n274_), .A2(new_n353_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n348_), .A2(KEYINPUT33), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT33), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n335_), .A2(new_n407_), .A3(new_n336_), .A4(new_n341_), .ZN(new_n408_));
  OR3_X1    g207(.A1(new_n344_), .A2(new_n345_), .A3(KEYINPUT100), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT100), .B1(new_n344_), .B2(new_n345_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n332_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n332_), .B1(new_n345_), .B2(new_n333_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n341_), .B1(new_n330_), .B2(new_n412_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n406_), .A2(new_n408_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n395_), .A2(new_n414_), .A3(new_n396_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT101), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n395_), .A2(new_n414_), .A3(KEYINPUT101), .A4(new_n396_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n393_), .A2(KEYINPUT32), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n419_), .B(KEYINPUT102), .Z(new_n420_));
  NOR2_X1   g219(.A1(new_n400_), .A2(new_n402_), .ZN(new_n421_));
  OAI221_X1 g220(.A(new_n349_), .B1(new_n389_), .B2(new_n420_), .C1(new_n421_), .C2(new_n419_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n417_), .A2(new_n418_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n274_), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n272_), .A2(new_n273_), .A3(new_n349_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n404_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n326_), .A2(new_n352_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n405_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G29gat), .B(G36gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G43gat), .B(G50gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G15gat), .B(G22gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G8gat), .ZN(new_n434_));
  INV_X1    g233(.A(G1gat), .ZN(new_n435_));
  INV_X1    g234(.A(G8gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT80), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT80), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(G8gat), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n435_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT14), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n433_), .B(new_n434_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT80), .B(G8gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT14), .B1(new_n444_), .B2(new_n435_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n434_), .B1(new_n445_), .B2(new_n433_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n432_), .B1(new_n443_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G229gat), .A2(G233gat), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n430_), .A2(new_n431_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n430_), .A2(new_n431_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT15), .ZN(new_n452_));
  INV_X1    g251(.A(new_n434_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n437_), .A2(new_n439_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n441_), .B1(new_n454_), .B2(G1gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n433_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n453_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n442_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n447_), .B(new_n448_), .C1(new_n452_), .C2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT81), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n451_), .A3(new_n442_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n447_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n448_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n460_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  AOI211_X1 g263(.A(KEYINPUT81), .B(new_n448_), .C1(new_n447_), .C2(new_n461_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n459_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G113gat), .B(G141gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G169gat), .B(G197gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n467_), .B(new_n468_), .Z(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT82), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n459_), .B(new_n469_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n466_), .A2(KEYINPUT82), .A3(new_n470_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n429_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT65), .ZN(new_n478_));
  OAI211_X1 g277(.A(G85gat), .B(G92gat), .C1(new_n478_), .C2(KEYINPUT9), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n478_), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT66), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n483_), .B1(G99gat), .B2(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G99gat), .A2(G106gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n485_), .A2(KEYINPUT6), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n482_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(KEYINPUT6), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n483_), .A2(G99gat), .A3(G106gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(KEYINPUT66), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT10), .B(G99gat), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n481_), .B(new_n491_), .C1(G106gat), .C2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G57gat), .B(G64gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n495_));
  XOR2_X1   g294(.A(G71gat), .B(G78gat), .Z(new_n496_));
  OR2_X1    g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n496_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT8), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT67), .B1(new_n484_), .B2(new_n486_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT67), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n488_), .A2(new_n489_), .A3(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n502_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G85gat), .B(G92gat), .Z(new_n510_));
  AOI21_X1  g309(.A(new_n501_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n501_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(new_n491_), .B2(new_n508_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n493_), .B(new_n500_), .C1(new_n511_), .C2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n493_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n500_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G230gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT64), .ZN(new_n522_));
  INV_X1    g321(.A(new_n493_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n490_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT66), .B1(new_n488_), .B2(new_n489_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n508_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(new_n501_), .A3(new_n510_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT69), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n509_), .A2(new_n510_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n527_), .B(new_n528_), .C1(new_n529_), .C2(new_n501_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT69), .B1(new_n511_), .B2(new_n513_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n523_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n500_), .A2(KEYINPUT70), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT70), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n497_), .B(new_n534_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT12), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n520_), .B(new_n522_), .C1(new_n532_), .C2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT68), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n519_), .A2(new_n514_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n522_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n539_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  AOI211_X1 g341(.A(KEYINPUT68), .B(new_n522_), .C1(new_n519_), .C2(new_n514_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n538_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G120gat), .B(G148gat), .Z(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G176gat), .B(G204gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n544_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n549_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n538_), .B(new_n551_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n550_), .A2(KEYINPUT73), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT73), .B1(new_n550_), .B2(new_n552_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT13), .ZN(new_n555_));
  OR3_X1    g354(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n555_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n556_), .A2(KEYINPUT74), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(KEYINPUT74), .B1(new_n556_), .B2(new_n557_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G127gat), .B(G155gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT16), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G183gat), .B(G211gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n458_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n566_), .B1(new_n500_), .B2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n500_), .B2(new_n569_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n533_), .A2(new_n536_), .ZN(new_n572_));
  AOI211_X1 g371(.A(new_n565_), .B(new_n564_), .C1(new_n572_), .C2(new_n568_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n573_), .B1(new_n572_), .B2(new_n568_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G134gat), .B(G162gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT36), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n579_), .A2(new_n580_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT34), .Z(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT75), .B(KEYINPUT35), .Z(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n517_), .A2(new_n451_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n532_), .A2(new_n452_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n591_), .B2(KEYINPUT76), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n532_), .A2(new_n452_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT76), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n587_), .B1(new_n592_), .B2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n588_), .A2(new_n589_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n591_), .A2(new_n597_), .A3(KEYINPUT77), .A4(new_n587_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT77), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n588_), .A2(new_n587_), .A3(new_n589_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n599_), .B1(new_n593_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n581_), .B(new_n582_), .C1(new_n596_), .C2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n598_), .A2(new_n601_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n595_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n597_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n586_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n604_), .A2(new_n607_), .A3(new_n580_), .A4(new_n579_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n603_), .A2(new_n608_), .A3(KEYINPUT78), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT79), .B(KEYINPUT37), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n609_), .B(new_n611_), .ZN(new_n612_));
  AND4_X1   g411(.A1(new_n477_), .A2(new_n560_), .A3(new_n576_), .A4(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n435_), .A3(new_n349_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT38), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n274_), .A2(new_n353_), .A3(new_n404_), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n423_), .A2(new_n274_), .B1(new_n425_), .B2(new_n404_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n428_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n617_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n603_), .A2(new_n608_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n556_), .A2(new_n557_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n476_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n623_), .A2(new_n576_), .A3(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n350_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n614_), .A2(new_n615_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n616_), .A2(new_n627_), .A3(new_n628_), .ZN(G1324gat));
  INV_X1    g428(.A(new_n404_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n613_), .A2(new_n444_), .A3(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT103), .Z(new_n632_));
  OAI21_X1  g431(.A(G8gat), .B1(new_n626_), .B2(new_n404_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT104), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n634_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(KEYINPUT39), .A3(new_n636_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(KEYINPUT39), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n632_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n632_), .A2(new_n637_), .A3(KEYINPUT40), .A4(new_n638_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1325gat));
  INV_X1    g442(.A(G15gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n613_), .A2(new_n644_), .A3(new_n619_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n626_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n619_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n647_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(KEYINPUT41), .B1(new_n647_), .B2(G15gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT105), .Z(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n274_), .B(KEYINPUT106), .Z(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n646_), .B2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT42), .Z(new_n655_));
  NAND3_X1  g454(.A1(new_n613_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1327gat));
  INV_X1    g456(.A(new_n624_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n476_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n659_), .A3(new_n575_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n609_), .B(new_n610_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n620_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n620_), .B2(new_n662_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT44), .B(new_n661_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n350_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n621_), .A2(new_n576_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n477_), .A2(new_n658_), .A3(new_n672_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n350_), .A2(G29gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n673_), .B2(new_n674_), .ZN(G1328gat));
  OR2_X1    g474(.A1(new_n630_), .A2(KEYINPUT108), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n630_), .A2(KEYINPUT108), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n673_), .A2(G36gat), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT45), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT43), .B1(new_n429_), .B2(new_n612_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n620_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT44), .B1(new_n684_), .B2(new_n661_), .ZN(new_n685_));
  AOI211_X1 g484(.A(new_n667_), .B(new_n660_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT107), .B1(new_n687_), .B2(new_n630_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n668_), .A2(KEYINPUT107), .A3(new_n630_), .A4(new_n669_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G36gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n681_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n691_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n697_), .B1(new_n670_), .B2(new_n404_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(G36gat), .A3(new_n689_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n699_), .A2(new_n692_), .A3(new_n693_), .A4(new_n681_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n696_), .A2(new_n700_), .ZN(G1329gat));
  NAND3_X1  g500(.A1(new_n687_), .A2(G43gat), .A3(new_n619_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n673_), .A2(new_n428_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(G43gat), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(G1330gat));
  INV_X1    g505(.A(new_n673_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G50gat), .B1(new_n707_), .B2(new_n653_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n274_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(G50gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(new_n687_), .B2(new_n710_), .ZN(G1331gat));
  NOR3_X1   g510(.A1(new_n662_), .A2(new_n658_), .A3(new_n575_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n429_), .A2(new_n659_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n715_), .A2(KEYINPUT111), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(KEYINPUT111), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n349_), .A3(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(G57gat), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n560_), .A2(new_n659_), .A3(new_n575_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n623_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT112), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n720_), .A2(KEYINPUT112), .A3(new_n623_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n350_), .A2(new_n719_), .ZN(new_n726_));
  AOI22_X1  g525(.A1(new_n718_), .A2(new_n719_), .B1(new_n725_), .B2(new_n726_), .ZN(G1332gat));
  INV_X1    g526(.A(G64gat), .ZN(new_n728_));
  INV_X1    g527(.A(new_n678_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n715_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n725_), .A2(new_n729_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(G64gat), .ZN(new_n733_));
  AOI211_X1 g532(.A(KEYINPUT48), .B(new_n728_), .C1(new_n725_), .C2(new_n729_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(G1333gat));
  OR3_X1    g534(.A1(new_n714_), .A2(G71gat), .A3(new_n428_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n723_), .A2(new_n619_), .A3(new_n724_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(G71gat), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n737_), .B2(G71gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(KEYINPUT114), .B(new_n736_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1334gat));
  INV_X1    g544(.A(G78gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n715_), .A2(new_n746_), .A3(new_n653_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n725_), .A2(new_n653_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(G78gat), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT50), .B(new_n746_), .C1(new_n725_), .C2(new_n653_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(G1335gat));
  INV_X1    g551(.A(new_n560_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n753_), .A2(new_n672_), .A3(new_n713_), .ZN(new_n754_));
  INV_X1    g553(.A(G85gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n755_), .A3(new_n349_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n624_), .A2(new_n476_), .A3(new_n575_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(new_n349_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n759_), .B2(new_n755_), .ZN(G1336gat));
  INV_X1    g559(.A(G92gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n754_), .A2(new_n761_), .A3(new_n630_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n758_), .A2(new_n729_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n761_), .ZN(G1337gat));
  NAND2_X1  g563(.A1(new_n758_), .A2(new_n619_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n428_), .A2(new_n492_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n765_), .A2(G99gat), .B1(new_n754_), .B2(new_n766_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g567(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n758_), .A2(new_n709_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(G106gat), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(KEYINPUT52), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(KEYINPUT52), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(G106gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n754_), .A2(new_n776_), .A3(new_n709_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n769_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n774_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n777_), .B(new_n769_), .C1(new_n779_), .C2(new_n772_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n778_), .A2(new_n781_), .ZN(G1339gat));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n538_), .A2(KEYINPUT117), .A3(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n520_), .B1(new_n532_), .B2(new_n537_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n541_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n783_), .B1(new_n538_), .B2(KEYINPUT117), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n549_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT56), .B(new_n549_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n552_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT116), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n473_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n447_), .B(new_n463_), .C1(new_n452_), .C2(new_n458_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n469_), .B1(new_n462_), .B2(new_n448_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT118), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n800_), .B(new_n803_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n796_), .A2(new_n802_), .A3(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(KEYINPUT57), .A3(new_n621_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT119), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n621_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n805_), .A2(new_n811_), .A3(KEYINPUT57), .A4(new_n621_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n800_), .A2(new_n552_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n793_), .A2(KEYINPUT58), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n793_), .A2(new_n813_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n662_), .A2(new_n814_), .A3(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n807_), .A2(new_n810_), .A3(new_n812_), .A4(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n575_), .ZN(new_n820_));
  AND4_X1   g619(.A1(new_n476_), .A2(new_n556_), .A3(new_n557_), .A4(new_n576_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n821_), .A2(new_n612_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n821_), .B2(new_n612_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n820_), .A2(new_n826_), .ZN(new_n827_));
  NOR4_X1   g626(.A1(new_n709_), .A2(new_n630_), .A3(new_n350_), .A4(new_n428_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(G113gat), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n659_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n829_), .B2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n827_), .A2(KEYINPUT120), .A3(KEYINPUT59), .A4(new_n828_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n476_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n832_), .B1(new_n837_), .B2(new_n831_), .ZN(G1340gat));
  INV_X1    g637(.A(G120gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n658_), .B2(KEYINPUT60), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n830_), .B(new_n840_), .C1(KEYINPUT60), .C2(new_n839_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n560_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n839_), .ZN(G1341gat));
  INV_X1    g642(.A(G127gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n829_), .B2(new_n575_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT121), .B(new_n844_), .C1(new_n829_), .C2(new_n575_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n576_), .A2(G127gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  INV_X1    g652(.A(new_n621_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n830_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n612_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n853_), .ZN(G1343gat));
  AOI21_X1  g656(.A(new_n619_), .B1(new_n820_), .B2(new_n826_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n729_), .A2(new_n350_), .A3(new_n274_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n659_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g662(.A1(new_n860_), .A2(new_n560_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT122), .B(G148gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1345gat));
  NAND2_X1  g665(.A1(new_n861_), .A2(new_n576_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1346gat));
  OR3_X1    g668(.A1(new_n860_), .A2(G162gat), .A3(new_n621_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G162gat), .B1(new_n860_), .B2(new_n612_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1347gat));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n729_), .A2(new_n353_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n653_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n827_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n476_), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT123), .B(new_n873_), .C1(new_n877_), .C2(new_n292_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(new_n375_), .A3(new_n298_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n292_), .B1(new_n880_), .B2(KEYINPUT62), .ZN(new_n881_));
  OAI221_X1 g680(.A(new_n881_), .B1(new_n880_), .B2(KEYINPUT62), .C1(new_n876_), .C2(new_n476_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n878_), .A2(new_n879_), .A3(new_n882_), .ZN(G1348gat));
  OAI21_X1  g682(.A(new_n293_), .B1(new_n876_), .B2(new_n658_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n885_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n825_), .B1(new_n819_), .B2(new_n575_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n709_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n874_), .A2(new_n560_), .A3(new_n293_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n886_), .A2(new_n887_), .B1(new_n889_), .B2(new_n890_), .ZN(G1349gat));
  NOR3_X1   g690(.A1(new_n876_), .A2(new_n305_), .A3(new_n575_), .ZN(new_n892_));
  INV_X1    g691(.A(G183gat), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n889_), .A2(new_n353_), .A3(new_n576_), .A4(new_n729_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1350gat));
  OAI21_X1  g694(.A(G190gat), .B1(new_n876_), .B2(new_n612_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n854_), .A2(new_n306_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n876_), .B2(new_n897_), .ZN(G1351gat));
  NAND2_X1  g697(.A1(new_n729_), .A2(new_n425_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n827_), .A2(new_n428_), .A3(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n858_), .A2(KEYINPUT125), .A3(new_n900_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G197gat), .B1(new_n905_), .B2(new_n659_), .ZN(new_n906_));
  AOI21_X1  g705(.A(KEYINPUT125), .B1(new_n858_), .B2(new_n900_), .ZN(new_n907_));
  NOR4_X1   g706(.A1(new_n888_), .A2(new_n902_), .A3(new_n619_), .A4(new_n899_), .ZN(new_n908_));
  OAI211_X1 g707(.A(G197gat), .B(new_n659_), .C1(new_n907_), .C2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n906_), .A2(new_n910_), .ZN(G1352gat));
  OAI21_X1  g710(.A(new_n753_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n912_), .A2(new_n913_), .A3(G204gat), .ZN(new_n914_));
  OAI221_X1 g713(.A(new_n753_), .B1(KEYINPUT126), .B2(new_n237_), .C1(new_n907_), .C2(new_n908_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1353gat));
  OR2_X1    g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n905_), .B2(new_n576_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT63), .B(G211gat), .Z(new_n919_));
  OAI211_X1 g718(.A(new_n576_), .B(new_n919_), .C1(new_n907_), .C2(new_n908_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n918_), .A2(new_n921_), .ZN(G1354gat));
  INV_X1    g721(.A(G218gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n854_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n662_), .A2(G218gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT127), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n923_), .A2(new_n924_), .B1(new_n905_), .B2(new_n926_), .ZN(G1355gat));
endmodule


