//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT76), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n206_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n209_), .A2(new_n210_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G1gat), .B(G8gat), .ZN(new_n213_));
  OR3_X1    g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n213_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n205_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n214_), .A2(new_n215_), .A3(new_n204_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G229gat), .A2(G233gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n216_), .B(new_n204_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(new_n219_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G113gat), .B(G141gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT78), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G169gat), .B(G197gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n220_), .B(new_n226_), .C1(new_n221_), .C2(new_n219_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT82), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n233_), .A2(KEYINPUT83), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(KEYINPUT83), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G113gat), .B(G120gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n234_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT31), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n232_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n243_), .B1(new_n242_), .B2(new_n241_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G71gat), .B(G99gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n244_), .B(new_n245_), .Z(new_n246_));
  INV_X1    g045(.A(KEYINPUT80), .ZN(new_n247_));
  AOI21_X1  g046(.A(G176gat), .B1(new_n247_), .B2(KEYINPUT22), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(G169gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT23), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(G183gat), .A3(G190gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n251_), .B1(G183gat), .B2(G190gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n249_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n252_), .A2(KEYINPUT79), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n252_), .A2(KEYINPUT79), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n254_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT25), .B(G183gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G190gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G169gat), .A2(G176gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT24), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(G169gat), .ZN(new_n266_));
  INV_X1    g065(.A(G176gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT24), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n262_), .B(new_n265_), .C1(new_n263_), .C2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n256_), .B1(new_n259_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G227gat), .A2(G233gat), .ZN(new_n271_));
  INV_X1    g070(.A(G15gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT30), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n270_), .B(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(KEYINPUT81), .B(G43gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n246_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n246_), .A2(new_n277_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT84), .ZN(new_n281_));
  INV_X1    g080(.A(G155gat), .ZN(new_n282_));
  INV_X1    g081(.A(G162gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT3), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT2), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n287_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G141gat), .B(G148gat), .Z(new_n293_));
  NAND2_X1  g092(.A1(new_n285_), .A2(KEYINPUT1), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n285_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(G155gat), .A3(G162gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n284_), .A2(new_n300_), .A3(new_n286_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n293_), .B1(new_n298_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT86), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OAI211_X1 g103(.A(KEYINPUT86), .B(new_n293_), .C1(new_n298_), .C2(new_n301_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n292_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT96), .B1(new_n306_), .B2(new_n241_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n292_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n284_), .A2(new_n286_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n309_), .A2(new_n300_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT86), .B1(new_n310_), .B2(new_n293_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n305_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n308_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n241_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n307_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n314_), .A3(KEYINPUT96), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(KEYINPUT4), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT4), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT99), .ZN(new_n325_));
  XOR2_X1   g124(.A(G1gat), .B(G29gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(G57gat), .B(G85gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  AOI21_X1  g129(.A(new_n323_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n324_), .A2(new_n325_), .A3(new_n330_), .A4(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n330_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n322_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(new_n331_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n331_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n325_), .B1(new_n338_), .B2(new_n330_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT28), .B1(new_n313_), .B2(KEYINPUT29), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n306_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT87), .ZN(new_n346_));
  XOR2_X1   g145(.A(G22gat), .B(G50gat), .Z(new_n347_));
  INV_X1    g146(.A(KEYINPUT87), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n341_), .A2(new_n348_), .A3(new_n344_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n346_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n347_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n341_), .A2(new_n348_), .A3(new_n344_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n348_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G78gat), .B(G106gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT91), .ZN(new_n356_));
  OR2_X1    g155(.A1(G197gat), .A2(G204gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G197gat), .A2(G204gat), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(KEYINPUT89), .A3(KEYINPUT21), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT89), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n357_), .A2(new_n358_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT21), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n364_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n360_), .A2(new_n361_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT90), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n361_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n361_), .A2(new_n368_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n369_), .A2(KEYINPUT21), .A3(new_n370_), .A4(new_n359_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n367_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(new_n306_), .B2(new_n343_), .ZN(new_n373_));
  INV_X1    g172(.A(G233gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT88), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(G228gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(G228gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n374_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n372_), .B(new_n381_), .C1(new_n306_), .C2(new_n343_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n356_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n383_), .A2(KEYINPUT92), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n380_), .A2(new_n356_), .A3(new_n382_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n383_), .B2(KEYINPUT92), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n350_), .B(new_n354_), .C1(new_n384_), .C2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n354_), .A2(new_n350_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT93), .ZN(new_n389_));
  INV_X1    g188(.A(new_n385_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(new_n383_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n388_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n389_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n387_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G226gat), .A2(G233gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT19), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT20), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n398_), .B1(new_n270_), .B2(new_n372_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n266_), .A2(new_n267_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT22), .B(G169gat), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n401_), .B2(new_n267_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(new_n259_), .B2(new_n250_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT95), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT95), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n405_), .B(new_n402_), .C1(new_n259_), .C2(new_n250_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n269_), .A2(new_n255_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n397_), .B(new_n399_), .C1(new_n408_), .C2(new_n372_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT20), .B1(new_n270_), .B2(new_n372_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n408_), .B2(new_n372_), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n396_), .B(KEYINPUT94), .Z(new_n412_));
  OAI21_X1  g211(.A(new_n409_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G8gat), .B(G36gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT18), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G64gat), .B(G92gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n418_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n409_), .B(new_n417_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n407_), .A2(new_n371_), .A3(new_n367_), .A4(new_n403_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n397_), .B1(new_n399_), .B2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n420_), .B(KEYINPUT27), .C1(new_n426_), .C2(new_n417_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n423_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n340_), .A2(new_n394_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n417_), .A2(KEYINPUT32), .ZN(new_n431_));
  MUX2_X1   g230(.A(new_n426_), .B(new_n413_), .S(new_n431_), .Z(new_n432_));
  OAI21_X1  g231(.A(new_n432_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n338_), .A2(new_n330_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n338_), .B(new_n330_), .C1(KEYINPUT98), .C2(KEYINPUT33), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n321_), .A2(new_n322_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n316_), .A2(new_n317_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n330_), .B1(new_n439_), .B2(new_n323_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n421_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n436_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n394_), .B1(new_n433_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n280_), .B1(new_n430_), .B2(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n423_), .A2(KEYINPUT100), .A3(new_n427_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT100), .B1(new_n423_), .B2(new_n427_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n394_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n280_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n448_), .A2(new_n340_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n231_), .B1(new_n444_), .B2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G190gat), .B(G218gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G134gat), .B(G162gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n455_), .B(KEYINPUT36), .Z(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(G85gat), .A2(G92gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G85gat), .A2(G92gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(KEYINPUT9), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT65), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT64), .B(G92gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT9), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(G85gat), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n460_), .B(new_n461_), .C1(new_n462_), .C2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G99gat), .ZN(new_n466_));
  INV_X1    g265(.A(G106gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT6), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(G99gat), .A3(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT10), .B(G99gat), .Z(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n467_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n465_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n460_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT65), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT8), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n468_), .A2(new_n470_), .B1(KEYINPUT66), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT66), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n481_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT67), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G99gat), .A2(G106gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NOR4_X1   g285(.A1(KEYINPUT67), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n480_), .B(new_n482_), .C1(new_n486_), .C2(new_n487_), .ZN(new_n488_));
  AND2_X1   g287(.A1(G85gat), .A2(G92gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G85gat), .A2(G92gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT68), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT68), .B1(new_n458_), .B2(new_n459_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n478_), .B1(new_n488_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n479_), .A2(KEYINPUT66), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n471_), .A2(new_n482_), .A3(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n487_), .A2(new_n486_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n494_), .B(new_n478_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n477_), .B1(new_n495_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n205_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n494_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT8), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n504_), .A2(new_n499_), .B1(new_n476_), .B2(new_n474_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n204_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n502_), .A2(new_n506_), .A3(KEYINPUT73), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G232gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT34), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT72), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT35), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n502_), .A2(new_n506_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n507_), .B(new_n512_), .C1(new_n513_), .C2(new_n509_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(KEYINPUT73), .A3(new_n511_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n457_), .B1(new_n516_), .B2(KEYINPUT75), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(KEYINPUT75), .B2(new_n516_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT37), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n455_), .A2(KEYINPUT36), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n514_), .A2(new_n520_), .A3(new_n515_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n518_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n516_), .A2(new_n456_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT37), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT74), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT74), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n524_), .A2(new_n527_), .A3(KEYINPUT37), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n522_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT71), .ZN(new_n531_));
  XOR2_X1   g330(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n532_));
  XNOR2_X1  g331(.A(G57gat), .B(G64gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT11), .ZN(new_n534_));
  XOR2_X1   g333(.A(G71gat), .B(G78gat), .Z(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n534_), .A2(new_n535_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n533_), .A2(KEYINPUT11), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n536_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n532_), .B1(new_n505_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n501_), .A2(KEYINPUT12), .A3(new_n540_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G230gat), .A2(G233gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n504_), .A2(new_n499_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(new_n541_), .A3(new_n477_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .A4(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n544_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n546_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n505_), .A2(new_n541_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(G120gat), .B(G148gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G176gat), .B(G204gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n547_), .A2(new_n551_), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n531_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n547_), .A2(new_n551_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n556_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n547_), .A2(new_n551_), .A3(new_n556_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(KEYINPUT71), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n559_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(KEYINPUT13), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(KEYINPUT13), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n541_), .B(new_n216_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G127gat), .B(G155gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT17), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n573_), .A2(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n578_), .A2(KEYINPUT17), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n573_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n530_), .A2(new_n570_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n452_), .A2(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n585_), .A2(G1gat), .A3(new_n340_), .ZN(new_n586_));
  XOR2_X1   g385(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n587_));
  AND2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n586_), .A2(new_n587_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n518_), .A2(new_n521_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n444_), .B2(new_n451_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n570_), .A2(new_n231_), .A3(new_n583_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n340_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n207_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n588_), .A2(new_n589_), .A3(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT102), .ZN(G1324gat));
  INV_X1    g397(.A(new_n585_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(new_n208_), .A3(new_n447_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT103), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n592_), .A2(new_n593_), .A3(new_n602_), .A4(new_n447_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n603_), .A2(G8gat), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n592_), .A2(new_n447_), .A3(new_n593_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT103), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n601_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  AND4_X1   g406(.A1(new_n601_), .A2(new_n606_), .A3(G8gat), .A4(new_n603_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n600_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT40), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(G1325gat));
  AOI21_X1  g410(.A(new_n272_), .B1(new_n594_), .B2(new_n450_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT41), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n599_), .A2(new_n272_), .A3(new_n450_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1326gat));
  INV_X1    g414(.A(G22gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n394_), .B(KEYINPUT104), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n616_), .B1(new_n594_), .B2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT42), .Z(new_n619_));
  NAND3_X1  g418(.A1(new_n599_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1327gat));
  INV_X1    g420(.A(new_n583_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n590_), .A2(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n623_), .A2(new_n569_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n452_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(G29gat), .B1(new_n625_), .B2(new_n595_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n569_), .A2(new_n230_), .A3(new_n583_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT105), .Z(new_n628_));
  INV_X1    g427(.A(KEYINPUT43), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n444_), .A2(new_n451_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n530_), .ZN(new_n631_));
  AOI211_X1 g430(.A(KEYINPUT43), .B(new_n529_), .C1(new_n444_), .C2(new_n451_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT106), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT44), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n628_), .B(KEYINPUT106), .C1(new_n631_), .C2(new_n632_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n628_), .B(KEYINPUT44), .C1(new_n631_), .C2(new_n632_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n639_), .A2(G29gat), .A3(new_n595_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n626_), .B1(new_n638_), .B2(new_n640_), .ZN(G1328gat));
  INV_X1    g440(.A(KEYINPUT46), .ZN(new_n642_));
  INV_X1    g441(.A(G36gat), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n447_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n643_), .B1(new_n638_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT45), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n448_), .A2(G36gat), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n452_), .A2(new_n624_), .A3(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(KEYINPUT107), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(KEYINPUT107), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n647_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n649_), .A2(KEYINPUT107), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n649_), .A2(KEYINPUT107), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(KEYINPUT45), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n642_), .B1(new_n646_), .B2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n652_), .A2(new_n655_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT44), .B1(new_n633_), .B2(new_n634_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n644_), .B1(new_n659_), .B2(new_n637_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n658_), .B(KEYINPUT46), .C1(new_n660_), .C2(new_n643_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n657_), .A2(new_n661_), .ZN(G1329gat));
  AOI21_X1  g461(.A(G43gat), .B1(new_n625_), .B2(new_n450_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n639_), .A2(G43gat), .A3(new_n450_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n638_), .B2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(KEYINPUT47), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT47), .ZN(new_n667_));
  AOI211_X1 g466(.A(new_n667_), .B(new_n663_), .C1(new_n638_), .C2(new_n664_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1330gat));
  AOI21_X1  g468(.A(G50gat), .B1(new_n625_), .B2(new_n617_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n639_), .A2(G50gat), .A3(new_n394_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n638_), .B2(new_n671_), .ZN(G1331gat));
  NOR2_X1   g471(.A1(new_n569_), .A2(new_n230_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n630_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n530_), .A2(new_n583_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n676_), .A2(G57gat), .A3(new_n340_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n592_), .A2(new_n622_), .A3(new_n673_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n595_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n677_), .B1(G57gat), .B2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT108), .ZN(G1332gat));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n447_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G64gat), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n448_), .A2(G64gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n676_), .B2(new_n686_), .ZN(G1333gat));
  INV_X1    g486(.A(G71gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n678_), .B2(new_n450_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT49), .Z(new_n690_));
  INV_X1    g489(.A(new_n676_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(new_n688_), .A3(new_n450_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1334gat));
  INV_X1    g492(.A(G78gat), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n617_), .A2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT110), .Z(new_n696_));
  NAND2_X1  g495(.A1(new_n691_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n694_), .B1(new_n678_), .B2(new_n617_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT50), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n698_), .A2(new_n699_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT111), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT111), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n704_), .B(new_n697_), .C1(new_n700_), .C2(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1335gat));
  INV_X1    g505(.A(KEYINPUT113), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n529_), .B1(new_n444_), .B2(new_n451_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(new_n629_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n569_), .A2(new_n230_), .A3(new_n622_), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT112), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n707_), .B1(new_n711_), .B2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n709_), .A2(KEYINPUT112), .A3(new_n710_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n712_), .A2(new_n713_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n717_), .A3(KEYINPUT113), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n715_), .A2(new_n595_), .A3(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G85gat), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n674_), .A2(new_n623_), .ZN(new_n721_));
  OR3_X1    g520(.A1(new_n721_), .A2(G85gat), .A3(new_n340_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1336gat));
  INV_X1    g522(.A(new_n721_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G92gat), .B1(new_n724_), .B2(new_n447_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n715_), .A2(new_n718_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n448_), .A2(new_n462_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT114), .Z(new_n728_));
  AOI21_X1  g527(.A(new_n725_), .B1(new_n726_), .B2(new_n728_), .ZN(G1337gat));
  NAND3_X1  g528(.A1(new_n724_), .A2(new_n450_), .A3(new_n472_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n280_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(new_n466_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT51), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n734_), .B(new_n730_), .C1(new_n731_), .C2(new_n466_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1338gat));
  NAND3_X1  g535(.A1(new_n724_), .A2(new_n467_), .A3(new_n394_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n394_), .B(new_n710_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(G106gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G106gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n230_), .A2(new_n744_), .A3(new_n563_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n230_), .B2(new_n563_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n547_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT116), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT116), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n547_), .A2(new_n751_), .A3(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n544_), .A2(new_n748_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n542_), .A2(new_n543_), .A3(new_n546_), .A4(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n548_), .A2(KEYINPUT117), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n755_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n542_), .A2(new_n543_), .A3(new_n546_), .A4(new_n757_), .ZN(new_n758_));
  AOI22_X1  g557(.A1(new_n750_), .A2(new_n752_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT56), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n556_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n759_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n756_), .A2(new_n758_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n547_), .A2(new_n751_), .A3(new_n748_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n751_), .B1(new_n547_), .B2(new_n748_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT56), .B1(new_n767_), .B2(new_n561_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n747_), .B1(new_n763_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n219_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n217_), .A2(new_n218_), .A3(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n227_), .C1(new_n221_), .C2(new_n770_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n229_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n565_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT118), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n565_), .A2(new_n777_), .A3(new_n774_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n769_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(KEYINPUT57), .A3(new_n590_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n777_), .B1(new_n565_), .B2(new_n774_), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT118), .B(new_n773_), .C1(new_n559_), .C2(new_n564_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n591_), .B1(new_n783_), .B2(new_n769_), .ZN(new_n784_));
  XOR2_X1   g583(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n785_));
  OAI21_X1  g584(.A(new_n780_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n760_), .B1(new_n759_), .B2(new_n556_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT120), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n767_), .A2(KEYINPUT120), .A3(new_n761_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n557_), .A2(new_n773_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n791_), .A2(KEYINPUT58), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT58), .B1(new_n791_), .B2(new_n792_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n529_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT121), .B1(new_n786_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n791_), .A2(new_n792_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n791_), .A2(KEYINPUT58), .A3(new_n792_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n530_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n779_), .A2(new_n590_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n785_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT121), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n801_), .A2(new_n804_), .A3(new_n805_), .A4(new_n780_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n796_), .A2(new_n583_), .A3(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n529_), .A2(new_n231_), .A3(new_n569_), .A4(new_n622_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT54), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  NOR4_X1   g609(.A1(new_n447_), .A2(new_n340_), .A3(new_n394_), .A4(new_n280_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT59), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n583_), .B1(new_n786_), .B2(new_n795_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n809_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n811_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n816_), .A2(KEYINPUT59), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n813_), .A2(new_n230_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G113gat), .ZN(new_n820_));
  OR3_X1    g619(.A1(new_n812_), .A2(G113gat), .A3(new_n231_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1340gat));
  AOI21_X1  g621(.A(new_n569_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n816_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT123), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT123), .B(new_n823_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(G120gat), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT60), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT122), .B1(new_n831_), .B2(G120gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(G120gat), .B1(new_n570_), .B2(new_n831_), .ZN(new_n833_));
  MUX2_X1   g632(.A(new_n832_), .B(KEYINPUT122), .S(new_n833_), .Z(new_n834_));
  NAND2_X1  g633(.A1(new_n824_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n830_), .A2(new_n835_), .ZN(G1341gat));
  NAND3_X1  g635(.A1(new_n813_), .A2(new_n622_), .A3(new_n818_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(G127gat), .ZN(new_n838_));
  OR3_X1    g637(.A1(new_n812_), .A2(G127gat), .A3(new_n583_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1342gat));
  NAND3_X1  g639(.A1(new_n813_), .A2(new_n530_), .A3(new_n818_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(G134gat), .ZN(new_n842_));
  OR3_X1    g641(.A1(new_n812_), .A2(G134gat), .A3(new_n590_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1343gat));
  NOR4_X1   g643(.A1(new_n449_), .A2(new_n447_), .A3(new_n340_), .A4(new_n450_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n810_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n230_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n570_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g649(.A1(new_n810_), .A2(new_n845_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n583_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT61), .B(G155gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1346gat));
  NAND3_X1  g653(.A1(new_n846_), .A2(new_n283_), .A3(new_n591_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G162gat), .B1(new_n851_), .B2(new_n529_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1347gat));
  INV_X1    g656(.A(new_n815_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(new_n617_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n448_), .A2(new_n595_), .A3(new_n280_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n859_), .A2(new_n401_), .A3(new_n230_), .A4(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n230_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT124), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n859_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n862_), .B1(new_n865_), .B2(G169gat), .ZN(new_n866_));
  AOI211_X1 g665(.A(KEYINPUT62), .B(new_n266_), .C1(new_n859_), .C2(new_n864_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n861_), .B1(new_n866_), .B2(new_n867_), .ZN(G1348gat));
  NAND3_X1  g667(.A1(new_n859_), .A2(new_n570_), .A3(new_n860_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n394_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n860_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n871_), .A2(new_n569_), .A3(new_n267_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n869_), .A2(new_n267_), .B1(new_n870_), .B2(new_n872_), .ZN(G1349gat));
  NOR2_X1   g672(.A1(new_n871_), .A2(new_n583_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G183gat), .B1(new_n870_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n260_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n622_), .A2(new_n876_), .ZN(new_n877_));
  NOR4_X1   g676(.A1(new_n858_), .A2(new_n617_), .A3(new_n871_), .A4(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT125), .ZN(new_n879_));
  OR3_X1    g678(.A1(new_n875_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n875_), .B2(new_n878_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1350gat));
  NAND4_X1  g681(.A1(new_n859_), .A2(new_n261_), .A3(new_n591_), .A4(new_n860_), .ZN(new_n883_));
  INV_X1    g682(.A(G190gat), .ZN(new_n884_));
  NOR4_X1   g683(.A1(new_n858_), .A2(new_n529_), .A3(new_n617_), .A4(new_n871_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1351gat));
  NAND3_X1  g685(.A1(new_n340_), .A2(new_n394_), .A3(new_n280_), .ZN(new_n887_));
  XOR2_X1   g686(.A(new_n887_), .B(KEYINPUT126), .Z(new_n888_));
  AOI211_X1 g687(.A(new_n448_), .B(new_n888_), .C1(new_n807_), .C2(new_n809_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n230_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n570_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g692(.A(new_n583_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n889_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT127), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n895_), .B(new_n897_), .ZN(G1354gat));
  INV_X1    g697(.A(G218gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n889_), .A2(new_n899_), .A3(new_n591_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n889_), .A2(new_n530_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(G1355gat));
endmodule


