//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n929_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT36), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT6), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT10), .B(G99gat), .Z(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n209_), .B2(G106gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G85gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G92gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  AOI22_X1  g013(.A1(new_n212_), .A2(new_n213_), .B1(KEYINPUT9), .B2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT7), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT7), .ZN(new_n223_));
  OAI211_X1 g022(.A(KEYINPUT66), .B(new_n222_), .C1(new_n223_), .C2(new_n221_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n207_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n221_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(KEYINPUT65), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n219_), .A2(KEYINPUT7), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n226_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT66), .B1(new_n230_), .B2(new_n222_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n218_), .B1(new_n225_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n227_), .A2(KEYINPUT65), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n221_), .B1(new_n220_), .B2(new_n236_), .ZN(new_n237_));
  AOI211_X1 g036(.A(G99gat), .B(G106gat), .C1(new_n219_), .C2(KEYINPUT7), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n235_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(new_n207_), .A3(new_n224_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(KEYINPUT67), .A3(new_n218_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n234_), .A2(KEYINPUT8), .A3(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n230_), .A2(new_n207_), .A3(new_n222_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT8), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n218_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n216_), .B1(new_n242_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G29gat), .B(G36gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G43gat), .B(G50gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT15), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT71), .B1(new_n246_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n253_));
  INV_X1    g052(.A(new_n245_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT67), .B1(new_n240_), .B2(new_n218_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(new_n244_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n254_), .B1(new_n256_), .B2(new_n241_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n253_), .B(new_n250_), .C1(new_n257_), .C2(new_n216_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G232gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT34), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT35), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n263_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT72), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n259_), .A2(new_n265_), .A3(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n265_), .B1(new_n259_), .B2(new_n268_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n205_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n216_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n240_), .A2(KEYINPUT67), .A3(new_n218_), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n273_), .A2(new_n255_), .A3(new_n244_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n272_), .B1(new_n274_), .B2(new_n254_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n253_), .B1(new_n275_), .B2(new_n250_), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n246_), .A2(KEYINPUT71), .A3(new_n251_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n268_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n264_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n259_), .A2(new_n265_), .A3(new_n268_), .ZN(new_n280_));
  XOR2_X1   g079(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n281_));
  NAND2_X1  g080(.A1(new_n204_), .A2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n282_), .B(KEYINPUT74), .Z(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n271_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n285_), .A2(KEYINPUT37), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n271_), .A2(KEYINPUT76), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(KEYINPUT75), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT76), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n289_), .B(new_n205_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT75), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n279_), .A2(new_n291_), .A3(new_n280_), .A4(new_n283_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n287_), .A2(new_n288_), .A3(new_n290_), .A4(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n286_), .B1(new_n293_), .B2(KEYINPUT37), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G57gat), .B(G64gat), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n295_), .A2(KEYINPUT11), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(KEYINPUT11), .ZN(new_n297_));
  XOR2_X1   g096(.A(G71gat), .B(G78gat), .Z(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n297_), .A2(new_n298_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G231gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT77), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G15gat), .B(G22gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G1gat), .A2(G8gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT14), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G1gat), .B(G8gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n308_), .B(new_n309_), .Z(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n304_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G183gat), .B(G211gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT79), .ZN(new_n314_));
  XOR2_X1   g113(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G127gat), .B(G155gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT17), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n312_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT17), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n312_), .B1(new_n321_), .B2(new_n318_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n294_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT80), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT12), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT68), .ZN(new_n329_));
  INV_X1    g128(.A(new_n301_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n275_), .A2(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n246_), .A2(new_n301_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n329_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G230gat), .A2(G233gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G120gat), .B(G148gat), .Z(new_n341_));
  XNOR2_X1  g140(.A(G176gat), .B(G204gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT69), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n340_), .B(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT13), .ZN(new_n348_));
  INV_X1    g147(.A(new_n346_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n340_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT13), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n310_), .B(new_n249_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(G229gat), .A3(G233gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n250_), .A2(new_n311_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n310_), .A2(new_n249_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G229gat), .A2(G233gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n358_), .B(KEYINPUT81), .Z(new_n359_));
  NAND3_X1  g158(.A1(new_n356_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G113gat), .B(G141gat), .Z(new_n362_));
  XNOR2_X1  g161(.A(G169gat), .B(G197gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n361_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n353_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G78gat), .B(G106gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G211gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n369_), .A2(G218gat), .ZN(new_n370_));
  INV_X1    g169(.A(G218gat), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n371_), .A2(G211gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT87), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(G197gat), .A2(G204gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G197gat), .A2(G204gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(KEYINPUT21), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT21), .ZN(new_n378_));
  INV_X1    g177(.A(new_n376_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n378_), .B1(new_n379_), .B2(new_n374_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n371_), .A2(G211gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n369_), .A2(G218gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT87), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n373_), .A2(new_n377_), .A3(new_n380_), .A4(new_n384_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n379_), .A2(new_n374_), .A3(new_n378_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n383_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n386_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(G228gat), .ZN(new_n391_));
  INV_X1    g190(.A(G233gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G141gat), .A2(G148gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT85), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT2), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT2), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n394_), .A2(KEYINPUT85), .A3(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n396_), .A2(new_n398_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(G155gat), .B(G162gat), .Z(new_n404_));
  NAND2_X1  g203(.A1(G155gat), .A2(G162gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT1), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT1), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(G155gat), .A3(G162gat), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n406_), .B(new_n408_), .C1(G155gat), .C2(G162gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n399_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n410_), .A2(new_n394_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n403_), .A2(new_n404_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT29), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n393_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT88), .B(KEYINPUT29), .Z(new_n417_));
  OAI21_X1  g216(.A(new_n390_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n391_), .A2(new_n392_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(KEYINPUT89), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT89), .B1(new_n418_), .B2(new_n419_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n368_), .B(new_n416_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT91), .ZN(new_n425_));
  XOR2_X1   g224(.A(G22gat), .B(G50gat), .Z(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n403_), .A2(new_n404_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n409_), .A2(new_n411_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT28), .B1(new_n430_), .B2(KEYINPUT29), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT86), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT28), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n412_), .A2(new_n433_), .A3(new_n413_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n432_), .B1(new_n431_), .B2(new_n434_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n427_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n437_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n426_), .A3(new_n435_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n424_), .A2(new_n425_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n416_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n367_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT90), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n443_), .A2(new_n444_), .B1(KEYINPUT91), .B2(new_n423_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n441_), .B(new_n445_), .C1(new_n444_), .C2(new_n443_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n423_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(new_n440_), .A3(new_n438_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G8gat), .B(G36gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT18), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G64gat), .B(G92gat), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n451_), .B(new_n452_), .Z(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G226gat), .A2(G233gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT93), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G183gat), .A2(G190gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G183gat), .A2(G190gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT82), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT82), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(G183gat), .A3(G190gat), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT23), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT23), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(G183gat), .B2(G190gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n461_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT95), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(KEYINPUT95), .B(new_n461_), .C1(new_n466_), .C2(new_n468_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT22), .B(G169gat), .ZN(new_n473_));
  INV_X1    g272(.A(G176gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G169gat), .A2(G176gat), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n471_), .A2(new_n472_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n463_), .A2(new_n465_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n480_), .B1(new_n481_), .B2(new_n467_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT25), .B(G183gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT26), .B(G190gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(G169gat), .A2(G176gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n487_), .A2(KEYINPUT24), .A3(new_n476_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT24), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n485_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n482_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n478_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT96), .B1(new_n493_), .B2(new_n390_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT96), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n385_), .A2(new_n389_), .ZN(new_n496_));
  AOI211_X1 g295(.A(new_n495_), .B(new_n496_), .C1(new_n478_), .C2(new_n492_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n483_), .A2(new_n484_), .B1(new_n489_), .B2(new_n486_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n499_), .B(new_n488_), .C1(new_n468_), .C2(new_n466_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n480_), .B(new_n461_), .C1(new_n481_), .C2(new_n467_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n477_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n496_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT20), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT94), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT94), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n463_), .A2(new_n465_), .ZN(new_n507_));
  AOI211_X1 g306(.A(new_n479_), .B(new_n460_), .C1(new_n507_), .C2(KEYINPUT23), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n475_), .A2(new_n476_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n466_), .A2(new_n468_), .ZN(new_n510_));
  OAI22_X1  g309(.A1(new_n508_), .A2(new_n509_), .B1(new_n491_), .B2(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n506_), .B(KEYINPUT20), .C1(new_n511_), .C2(new_n390_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n505_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n459_), .B1(new_n498_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n478_), .A2(new_n496_), .A3(new_n492_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n515_), .A2(KEYINPUT20), .A3(new_n457_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n390_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT97), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT97), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n511_), .A2(new_n519_), .A3(new_n390_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n454_), .B1(new_n514_), .B2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n482_), .A2(new_n491_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n509_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n525_), .B1(new_n526_), .B2(new_n472_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n495_), .B1(new_n527_), .B2(new_n496_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n493_), .A2(KEYINPUT96), .A3(new_n390_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n512_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n506_), .B1(new_n503_), .B2(KEYINPUT20), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n528_), .B(new_n529_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n458_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(new_n453_), .A3(new_n522_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n524_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT27), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(KEYINPUT27), .ZN(new_n538_));
  INV_X1    g337(.A(new_n457_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT102), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT101), .B(KEYINPUT20), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n515_), .A2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n521_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n541_), .B1(new_n527_), .B2(new_n496_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(KEYINPUT102), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n539_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n498_), .A2(new_n513_), .A3(new_n459_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n453_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n538_), .A2(new_n549_), .A3(KEYINPUT103), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT103), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n532_), .A2(new_n458_), .B1(new_n521_), .B2(new_n516_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n536_), .B1(new_n552_), .B2(new_n453_), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n545_), .A2(KEYINPUT102), .B1(new_n518_), .B2(new_n520_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n543_), .A2(new_n540_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n457_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n532_), .A2(new_n458_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n454_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n551_), .B1(new_n553_), .B2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n537_), .B1(new_n550_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT104), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT103), .B1(new_n538_), .B2(new_n549_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n553_), .A2(new_n558_), .A3(new_n551_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT104), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n565_), .A3(new_n537_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n449_), .B1(new_n561_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT83), .ZN(new_n568_));
  XOR2_X1   g367(.A(G127gat), .B(G134gat), .Z(new_n569_));
  XOR2_X1   g368(.A(G113gat), .B(G120gat), .Z(new_n570_));
  AOI21_X1  g369(.A(new_n568_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n570_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G127gat), .B(G134gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G113gat), .B(G120gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n571_), .B1(new_n576_), .B2(new_n568_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT4), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n430_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT98), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G225gat), .A2(G233gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT98), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n577_), .A2(new_n430_), .A3(new_n583_), .A4(new_n578_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n428_), .A2(new_n576_), .A3(new_n429_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n573_), .A2(new_n574_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n573_), .A2(new_n574_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n568_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n571_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n585_), .B(KEYINPUT4), .C1(new_n590_), .C2(new_n412_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n580_), .A2(new_n582_), .A3(new_n584_), .A4(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n577_), .A2(new_n430_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT99), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n593_), .A2(new_n596_), .A3(new_n581_), .A4(new_n585_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n592_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G1gat), .B(G29gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(G85gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT0), .B(G57gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n592_), .A2(new_n602_), .A3(new_n595_), .A4(new_n597_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G71gat), .B(G99gat), .ZN(new_n607_));
  INV_X1    g406(.A(G43gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n511_), .B(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G227gat), .A2(G233gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(G15gat), .Z(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT30), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT31), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n610_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT84), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n616_), .A2(new_n577_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n577_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n606_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  AND4_X1   g418(.A1(new_n581_), .A2(new_n580_), .A3(new_n584_), .A4(new_n591_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n593_), .A2(new_n582_), .A3(new_n585_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n603_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT33), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n605_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n605_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n524_), .A2(new_n624_), .A3(new_n626_), .A4(new_n534_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n605_), .A2(new_n625_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n605_), .B2(new_n623_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n631_), .A2(KEYINPUT100), .A3(new_n534_), .A4(new_n524_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n453_), .A2(KEYINPUT32), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n552_), .A2(new_n633_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n634_));
  OAI211_X1 g433(.A(KEYINPUT32), .B(new_n453_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n629_), .A2(new_n632_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n449_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n606_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n564_), .A2(new_n537_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n617_), .A2(new_n618_), .ZN(new_n643_));
  AOI22_X1  g442(.A1(new_n567_), .A2(new_n619_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n366_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n327_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n327_), .A2(KEYINPUT105), .A3(new_n645_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n606_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(G1gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n649_), .A3(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n285_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n324_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n645_), .A2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n658_), .B2(new_n650_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n648_), .A2(new_n649_), .A3(new_n651_), .A4(new_n653_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n655_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n655_), .A2(KEYINPUT107), .A3(new_n659_), .A4(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1324gat));
  NOR2_X1   g464(.A1(new_n560_), .A2(KEYINPUT104), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n565_), .B1(new_n564_), .B2(new_n537_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G8gat), .B1(new_n658_), .B2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT39), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n648_), .A2(new_n649_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n669_), .A2(G8gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n671_), .B(KEYINPUT40), .C1(new_n672_), .C2(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1325gat));
  OAI21_X1  g478(.A(G15gat), .B1(new_n658_), .B2(new_n643_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT41), .Z(new_n681_));
  OR2_X1    g480(.A1(new_n643_), .A2(G15gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n672_), .B2(new_n682_), .ZN(G1326gat));
  OAI21_X1  g482(.A(G22gat), .B1(new_n658_), .B2(new_n638_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT42), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n638_), .A2(G22gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n672_), .B2(new_n686_), .ZN(G1327gat));
  OAI211_X1 g486(.A(new_n638_), .B(new_n619_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n641_), .ZN(new_n689_));
  AOI22_X1  g488(.A1(new_n627_), .A2(new_n628_), .B1(new_n635_), .B2(new_n634_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n449_), .B1(new_n690_), .B2(new_n632_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n643_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n688_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n294_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n293_), .A2(KEYINPUT37), .ZN(new_n698_));
  INV_X1    g497(.A(new_n286_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT43), .B1(new_n644_), .B2(new_n700_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n693_), .A2(KEYINPUT108), .A3(new_n694_), .A4(new_n294_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n697_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n366_), .A2(new_n323_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(KEYINPUT44), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT44), .B1(new_n703_), .B2(new_n704_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(new_n650_), .ZN(new_n708_));
  INV_X1    g507(.A(G29gat), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n285_), .A2(new_n323_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n645_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n606_), .A2(new_n709_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT109), .ZN(new_n713_));
  OAI22_X1  g512(.A1(new_n708_), .A2(new_n709_), .B1(new_n711_), .B2(new_n713_), .ZN(G1328gat));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  INV_X1    g514(.A(G36gat), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n703_), .A2(new_n704_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n669_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n716_), .B1(new_n719_), .B2(new_n705_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n711_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n716_), .A3(new_n668_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n715_), .B1(new_n720_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n723_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n722_), .B(new_n726_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n706_), .A2(new_n707_), .A3(new_n669_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n727_), .B(KEYINPUT46), .C1(new_n728_), .C2(new_n716_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n725_), .A2(new_n729_), .ZN(G1329gat));
  NAND2_X1  g529(.A1(new_n717_), .A2(new_n718_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n643_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n731_), .A2(G43gat), .A3(new_n732_), .A4(new_n705_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n608_), .B1(new_n711_), .B2(new_n643_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT47), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n733_), .A2(new_n737_), .A3(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1330gat));
  AOI21_X1  g538(.A(G50gat), .B1(new_n721_), .B2(new_n449_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n731_), .A2(G50gat), .A3(new_n449_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(new_n705_), .ZN(G1331gat));
  NOR3_X1   g541(.A1(new_n644_), .A2(new_n365_), .A3(new_n353_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(new_n657_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G57gat), .B1(new_n745_), .B2(new_n650_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n327_), .A2(new_n743_), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n650_), .A2(G57gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n747_), .B2(new_n748_), .ZN(G1332gat));
  INV_X1    g548(.A(G64gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n744_), .B2(new_n668_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT48), .Z(new_n752_));
  INV_X1    g551(.A(new_n747_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n750_), .A3(new_n668_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1333gat));
  INV_X1    g554(.A(G71gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n744_), .B2(new_n732_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT49), .Z(new_n758_));
  NAND3_X1  g557(.A1(new_n753_), .A2(new_n756_), .A3(new_n732_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1334gat));
  OAI21_X1  g559(.A(G78gat), .B1(new_n745_), .B2(new_n638_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n638_), .A2(G78gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n747_), .B2(new_n764_), .ZN(G1335gat));
  AND2_X1   g564(.A1(new_n743_), .A2(new_n710_), .ZN(new_n766_));
  AOI21_X1  g565(.A(G85gat), .B1(new_n766_), .B2(new_n606_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n353_), .A2(new_n365_), .A3(new_n323_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n703_), .A2(new_n768_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n606_), .A2(new_n211_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n767_), .B1(new_n769_), .B2(new_n770_), .ZN(G1336gat));
  NAND3_X1  g570(.A1(new_n703_), .A2(new_n668_), .A3(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G92gat), .ZN(new_n773_));
  INV_X1    g572(.A(G92gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n766_), .A2(new_n774_), .A3(new_n668_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT112), .Z(G1337gat));
  NAND3_X1  g576(.A1(new_n703_), .A2(new_n732_), .A3(new_n768_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G99gat), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n643_), .A2(new_n209_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n743_), .A2(new_n710_), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT114), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n779_), .A2(new_n788_), .A3(new_n782_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n784_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n788_), .B1(new_n779_), .B2(new_n782_), .ZN(new_n791_));
  AOI211_X1 g590(.A(KEYINPUT114), .B(new_n781_), .C1(new_n778_), .C2(G99gat), .ZN(new_n792_));
  OAI22_X1  g591(.A1(new_n791_), .A2(new_n792_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(G1338gat));
  XNOR2_X1  g593(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n701_), .A2(new_n702_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n700_), .B1(new_n692_), .B2(new_n688_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT108), .B1(new_n797_), .B2(new_n694_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n449_), .B(new_n768_), .C1(new_n796_), .C2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G106gat), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT52), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n802_), .A3(G106gat), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(G106gat), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n766_), .A2(new_n805_), .A3(new_n449_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n795_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n799_), .A2(new_n802_), .A3(G106gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n802_), .B1(new_n799_), .B2(G106gat), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n806_), .B(new_n795_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n807_), .A2(new_n811_), .ZN(G1339gat));
  NAND2_X1  g611(.A1(new_n275_), .A2(new_n330_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n246_), .A2(new_n301_), .ZN(new_n814_));
  AOI22_X1  g613(.A1(new_n813_), .A2(new_n814_), .B1(KEYINPUT68), .B2(new_n328_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n332_), .A2(new_n334_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n815_), .A2(new_n338_), .A3(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n338_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(KEYINPUT55), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  NOR4_X1   g619(.A1(new_n815_), .A2(new_n816_), .A3(new_n820_), .A4(new_n338_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n345_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT56), .ZN(new_n823_));
  INV_X1    g622(.A(new_n345_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n337_), .A2(new_n339_), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n359_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n356_), .A2(new_n357_), .A3(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n364_), .B1(new_n354_), .B2(new_n359_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n361_), .A2(new_n364_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n825_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT119), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n825_), .A2(new_n832_), .A3(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n336_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n337_), .B1(new_n835_), .B2(new_n820_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n821_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n824_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT56), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n823_), .A2(new_n834_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n823_), .A2(new_n834_), .A3(new_n840_), .A4(KEYINPUT58), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n294_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n825_), .A2(new_n365_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n822_), .A2(new_n849_), .A3(KEYINPUT56), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n839_), .B1(new_n838_), .B2(KEYINPUT118), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n848_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n350_), .A2(new_n829_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n656_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n845_), .B1(new_n854_), .B2(KEYINPUT57), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n856_), .B(new_n656_), .C1(new_n852_), .C2(new_n853_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n324_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n365_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n325_), .A2(new_n859_), .A3(new_n353_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n858_), .A2(new_n862_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n567_), .A2(new_n606_), .A3(new_n732_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(G113gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n365_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n865_), .A2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n863_), .A2(KEYINPUT59), .A3(new_n864_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n859_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n868_), .B1(new_n872_), .B2(new_n867_), .ZN(G1340gat));
  XOR2_X1   g672(.A(KEYINPUT120), .B(G120gat), .Z(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n353_), .B2(KEYINPUT60), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n866_), .B(new_n875_), .C1(KEYINPUT60), .C2(new_n874_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n353_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n874_), .ZN(G1341gat));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n863_), .A2(new_n323_), .A3(new_n864_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(G127gat), .ZN(new_n881_));
  INV_X1    g680(.A(G127gat), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT121), .B(new_n882_), .C1(new_n865_), .C2(new_n324_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n870_), .A2(new_n871_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n324_), .A2(new_n882_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n881_), .A2(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1342gat));
  AND3_X1   g685(.A1(new_n863_), .A2(new_n656_), .A3(new_n864_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT122), .B1(new_n887_), .B2(G134gat), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889_));
  INV_X1    g688(.A(G134gat), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n889_), .B(new_n890_), .C1(new_n865_), .C2(new_n285_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n700_), .A2(new_n890_), .ZN(new_n892_));
  AOI22_X1  g691(.A1(new_n888_), .A2(new_n891_), .B1(new_n884_), .B2(new_n892_), .ZN(G1343gat));
  NAND2_X1  g692(.A1(new_n643_), .A2(new_n606_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n668_), .A2(new_n638_), .A3(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n365_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g698(.A1(new_n348_), .A2(new_n352_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n897_), .A2(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g701(.A(KEYINPUT61), .B(G155gat), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n897_), .A2(new_n905_), .A3(new_n323_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n897_), .B2(new_n323_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n904_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n863_), .A2(new_n323_), .A3(new_n895_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT123), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(new_n906_), .A3(new_n903_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n912_), .ZN(G1346gat));
  AOI21_X1  g712(.A(G162gat), .B1(new_n897_), .B2(new_n656_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n294_), .A2(G162gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT124), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n897_), .B2(new_n916_), .ZN(G1347gat));
  AND2_X1   g716(.A1(new_n619_), .A2(new_n638_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n863_), .A2(new_n668_), .A3(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919_), .B2(new_n859_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  OAI211_X1 g721(.A(KEYINPUT62), .B(G169gat), .C1(new_n919_), .C2(new_n859_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n919_), .A2(new_n859_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n473_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n922_), .A2(new_n923_), .A3(new_n925_), .ZN(G1348gat));
  NAND4_X1  g725(.A1(new_n863_), .A2(new_n900_), .A3(new_n668_), .A4(new_n918_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G176gat), .ZN(G1349gat));
  NAND4_X1  g727(.A1(new_n863_), .A2(new_n668_), .A3(new_n323_), .A4(new_n918_), .ZN(new_n929_));
  MUX2_X1   g728(.A(new_n483_), .B(G183gat), .S(new_n929_), .Z(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n919_), .B2(new_n700_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n656_), .A2(new_n484_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n919_), .B2(new_n932_), .ZN(G1351gat));
  NAND2_X1  g732(.A1(new_n643_), .A2(new_n640_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(KEYINPUT125), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n863_), .A2(new_n365_), .A3(new_n668_), .A4(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(G197gat), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n936_), .A2(KEYINPUT126), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(KEYINPUT126), .B1(new_n936_), .B2(new_n937_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n936_), .A2(new_n937_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n938_), .A2(new_n939_), .A3(new_n940_), .ZN(G1352gat));
  AND3_X1   g740(.A1(new_n863_), .A2(new_n668_), .A3(new_n935_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n900_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(G204gat), .ZN(new_n944_));
  INV_X1    g743(.A(G204gat), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n942_), .A2(new_n945_), .A3(new_n900_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n944_), .A2(new_n946_), .ZN(G1353gat));
  NAND4_X1  g746(.A1(new_n863_), .A2(new_n668_), .A3(new_n323_), .A4(new_n935_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n949_));
  AND2_X1   g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n948_), .A2(new_n949_), .A3(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n951_), .B1(new_n948_), .B2(new_n949_), .ZN(G1354gat));
  NAND2_X1  g751(.A1(new_n942_), .A2(new_n656_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n294_), .A2(G218gat), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(KEYINPUT127), .ZN(new_n955_));
  AOI22_X1  g754(.A1(new_n953_), .A2(new_n371_), .B1(new_n942_), .B2(new_n955_), .ZN(G1355gat));
endmodule


