//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n902_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G15gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G71gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT83), .B(G99gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT82), .B(G43gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT84), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT23), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(G169gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  AND2_X1   g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n235_), .A2(new_n224_), .ZN(new_n236_));
  AOI22_X1  g035(.A1(new_n231_), .A2(new_n234_), .B1(new_n236_), .B2(KEYINPUT24), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n227_), .B1(new_n237_), .B2(KEYINPUT80), .ZN(new_n238_));
  AND2_X1   g037(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n239_));
  AND2_X1   g038(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n241_));
  OAI22_X1  g040(.A1(new_n228_), .A2(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n224_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G169gat), .A2(G176gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(KEYINPUT24), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT80), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT81), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n212_), .A2(new_n248_), .A3(KEYINPUT23), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n248_), .B1(new_n212_), .B2(KEYINPUT23), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n246_), .A2(new_n247_), .B1(new_n251_), .B2(new_n215_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n223_), .B1(new_n238_), .B2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT30), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n210_), .B1(new_n211_), .B2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n211_), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  OR2_X1    g056(.A1(G113gat), .A2(G120gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G113gat), .A2(G120gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  OR2_X1    g059(.A1(G127gat), .A2(G134gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G127gat), .A2(G134gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT85), .B1(new_n260_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n263_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n258_), .A2(new_n261_), .A3(new_n262_), .A4(new_n259_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n264_), .B1(new_n267_), .B2(KEYINPUT85), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT31), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n257_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n216_), .A2(new_n226_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n237_), .A2(new_n279_), .A3(KEYINPUT90), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT90), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(new_n246_), .B2(new_n278_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n250_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n212_), .A2(new_n248_), .A3(KEYINPUT23), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n215_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n218_), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n280_), .A2(new_n282_), .B1(new_n221_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT21), .ZN(new_n288_));
  INV_X1    g087(.A(G197gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G204gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT88), .B(G204gat), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n288_), .B(new_n290_), .C1(new_n291_), .C2(new_n289_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G197gat), .A2(G204gat), .ZN(new_n293_));
  OAI211_X1 g092(.A(KEYINPUT21), .B(new_n293_), .C1(new_n291_), .C2(G197gat), .ZN(new_n294_));
  AND2_X1   g093(.A1(G211gat), .A2(G218gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G211gat), .A2(G218gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n292_), .A2(new_n294_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(KEYINPUT89), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT89), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n288_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n290_), .B1(new_n291_), .B2(new_n289_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n299_), .A2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT20), .B1(new_n287_), .B2(new_n305_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n229_), .A2(new_n230_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n235_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n247_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n242_), .A2(new_n245_), .A3(KEYINPUT80), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n309_), .A2(new_n285_), .A3(new_n226_), .A4(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n222_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n299_), .A2(new_n304_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT19), .ZN(new_n316_));
  NOR3_X1   g115(.A1(new_n306_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n316_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT20), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n286_), .A2(new_n221_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n305_), .B(new_n321_), .C1(new_n246_), .C2(new_n278_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n318_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n277_), .B1(new_n317_), .B2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT90), .B1(new_n237_), .B2(new_n279_), .ZN(new_n325_));
  NOR3_X1   g124(.A1(new_n246_), .A2(new_n278_), .A3(new_n281_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n321_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n318_), .B1(new_n327_), .B2(new_n313_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT20), .B1(new_n253_), .B2(new_n305_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT91), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n316_), .B1(new_n306_), .B2(new_n314_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n316_), .B1(new_n287_), .B2(new_n305_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT91), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n320_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n330_), .A2(new_n331_), .A3(new_n334_), .A4(new_n276_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n324_), .A2(new_n335_), .A3(KEYINPUT97), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT97), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n337_), .B(new_n277_), .C1(new_n317_), .C2(new_n323_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT27), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n330_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n277_), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT27), .B1(new_n342_), .B2(new_n335_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(G85gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT0), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n348_), .B(G57gat), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT94), .ZN(new_n351_));
  AND2_X1   g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT87), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT2), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT2), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(KEYINPUT87), .A3(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n360_));
  OR3_X1    g159(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n357_), .A2(new_n359_), .A3(new_n360_), .A4(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT1), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n353_), .B1(new_n352_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT1), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT86), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT86), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(new_n368_), .A3(KEYINPUT1), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n364_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G141gat), .B(G148gat), .Z(new_n371_));
  AOI22_X1  g170(.A1(new_n354_), .A2(new_n362_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n351_), .B1(new_n372_), .B2(new_n267_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n362_), .A2(new_n354_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(new_n371_), .ZN(new_n375_));
  AND4_X1   g174(.A1(new_n351_), .A2(new_n374_), .A3(new_n375_), .A4(new_n267_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n375_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n268_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n377_), .A2(KEYINPUT95), .A3(KEYINPUT4), .A4(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n267_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT94), .B1(new_n378_), .B2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n374_), .A2(new_n375_), .A3(new_n351_), .A4(new_n267_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n382_), .A2(KEYINPUT4), .A3(new_n379_), .A4(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT95), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n379_), .A2(KEYINPUT4), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n380_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n350_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  AOI211_X1 g193(.A(new_n349_), .B(new_n392_), .C1(new_n388_), .C2(new_n390_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n313_), .B1(new_n372_), .B2(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n398_), .A2(G50gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(G50gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G78gat), .B(G106gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n402_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n399_), .A2(new_n404_), .A3(new_n400_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  OR3_X1    g205(.A1(new_n378_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT28), .B1(new_n378_), .B2(KEYINPUT29), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(G22gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n409_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n412_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n406_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n403_), .A2(new_n413_), .A3(new_n414_), .A4(new_n405_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n396_), .A2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT98), .B1(new_n345_), .B2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n343_), .B1(new_n339_), .B2(KEYINPUT27), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT98), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n396_), .A4(new_n418_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n342_), .A2(new_n335_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT93), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n342_), .A2(KEYINPUT93), .A3(new_n335_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OR3_X1    g228(.A1(new_n388_), .A2(KEYINPUT96), .A3(new_n390_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n377_), .A2(new_n390_), .A3(new_n379_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT96), .B1(new_n388_), .B2(new_n390_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n430_), .A2(new_n350_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n392_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n434_), .B1(new_n435_), .B2(new_n350_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n394_), .A2(KEYINPUT33), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n429_), .A2(new_n433_), .A3(new_n436_), .A4(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n276_), .A2(KEYINPUT32), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(new_n317_), .B2(new_n323_), .ZN(new_n441_));
  OAI221_X1 g240(.A(new_n441_), .B1(new_n341_), .B2(new_n440_), .C1(new_n394_), .C2(new_n395_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n418_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n271_), .B1(new_n424_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT99), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n271_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n345_), .A2(new_n418_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n396_), .A3(new_n448_), .ZN(new_n449_));
  OAI211_X1 g248(.A(KEYINPUT99), .B(new_n271_), .C1(new_n424_), .C2(new_n443_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(G85gat), .A2(G92gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(G85gat), .A2(G92gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(G99gat), .A2(G106gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT7), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G99gat), .A2(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n454_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT67), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT8), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(KEYINPUT8), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n464_), .B(new_n454_), .C1(new_n457_), .C2(new_n460_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n467_));
  NAND2_X1  g266(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n467_), .B(new_n468_), .C1(G85gat), .C2(G92gat), .ZN(new_n469_));
  OR2_X1    g268(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(G92gat), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n452_), .A2(KEYINPUT9), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n460_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT10), .B(G99gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n476_), .A2(G106gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT66), .B1(new_n475_), .B2(new_n478_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n469_), .A2(new_n472_), .B1(KEYINPUT9), .B2(new_n452_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT66), .ZN(new_n481_));
  NOR4_X1   g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n460_), .A4(new_n477_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n466_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G57gat), .B(G64gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT11), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G71gat), .B(G78gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G71gat), .B(G78gat), .Z(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(KEYINPUT11), .A3(new_n484_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n484_), .A2(KEYINPUT11), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n487_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT68), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT68), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n487_), .A2(new_n489_), .A3(new_n490_), .A4(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n483_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT12), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G230gat), .A2(G233gat), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n495_), .B(new_n466_), .C1(new_n479_), .C2(new_n482_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n483_), .A2(KEYINPUT12), .A3(new_n491_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .A4(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(new_n501_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n500_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G120gat), .B(G148gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT5), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(G176gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(G204gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n503_), .A2(new_n506_), .A3(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n511_), .A2(KEYINPUT69), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(KEYINPUT69), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n503_), .A2(new_n506_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n510_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT70), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(KEYINPUT13), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(KEYINPUT13), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n519_), .A2(KEYINPUT13), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n514_), .B(new_n517_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT15), .ZN(new_n526_));
  OR2_X1    g325(.A1(G29gat), .A2(G36gat), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT71), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n528_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n532_));
  OAI21_X1  g331(.A(G43gat), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n527_), .A2(new_n529_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT71), .ZN(new_n535_));
  INV_X1    g334(.A(G43gat), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n536_), .A3(new_n530_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(G50gat), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(G50gat), .B1(new_n533_), .B2(new_n537_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n526_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n533_), .A2(new_n537_), .ZN(new_n542_));
  INV_X1    g341(.A(G50gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(KEYINPUT15), .A3(new_n538_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT76), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT75), .B(G15gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(G22gat), .ZN(new_n549_));
  INV_X1    g348(.A(G1gat), .ZN(new_n550_));
  INV_X1    g349(.A(G8gat), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT14), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n547_), .B1(new_n549_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G1gat), .B(G8gat), .Z(new_n555_));
  NAND3_X1  g354(.A1(new_n549_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n555_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n556_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n558_), .B1(new_n559_), .B2(new_n553_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n546_), .A2(new_n557_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n557_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n544_), .A2(new_n538_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n561_), .A2(new_n562_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n562_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n564_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(new_n557_), .A3(new_n560_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n568_), .B1(new_n560_), .B2(new_n557_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n567_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574_));
  INV_X1    g373(.A(G169gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(new_n289_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n577_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n566_), .A2(new_n572_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n525_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n451_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n483_), .A2(new_n541_), .A3(new_n545_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT73), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT34), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(KEYINPUT35), .A3(new_n588_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n564_), .B(new_n466_), .C1(new_n479_), .C2(new_n482_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT72), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n473_), .A2(new_n474_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n460_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n594_), .A3(new_n478_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n481_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n475_), .A2(KEYINPUT66), .A3(new_n478_), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n596_), .A2(new_n597_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(KEYINPUT72), .A3(new_n564_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n592_), .A2(new_n599_), .A3(new_n585_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n589_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n588_), .A2(KEYINPUT35), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT35), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n585_), .B2(KEYINPUT73), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n602_), .B1(new_n604_), .B2(new_n588_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n601_), .B1(new_n605_), .B2(new_n600_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(G134gat), .ZN(new_n609_));
  INV_X1    g408(.A(G162gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n607_), .A2(KEYINPUT36), .A3(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(KEYINPUT36), .ZN(new_n614_));
  INV_X1    g413(.A(new_n602_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n600_), .B1(new_n589_), .B2(new_n615_), .ZN(new_n616_));
  AOI22_X1  g415(.A1(new_n546_), .A2(new_n483_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n617_), .A2(new_n599_), .B1(new_n604_), .B2(new_n588_), .ZN(new_n618_));
  OAI211_X1 g417(.A(KEYINPUT74), .B(new_n614_), .C1(new_n616_), .C2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n614_), .B1(new_n606_), .B2(KEYINPUT74), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n613_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n563_), .B(new_n626_), .Z(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(new_n491_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n491_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n625_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G183gat), .B(G211gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G127gat), .B(G155gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n630_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT79), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT79), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n630_), .A2(new_n638_), .A3(new_n635_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n627_), .B(new_n495_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n635_), .B(KEYINPUT17), .Z(new_n641_));
  AOI22_X1  g440(.A1(new_n637_), .A2(new_n639_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n584_), .A2(new_n624_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G1gat), .B1(new_n645_), .B2(new_n396_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n584_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT37), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n622_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n613_), .B(KEYINPUT37), .C1(new_n620_), .C2(new_n621_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n651_), .A2(new_n642_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n647_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT100), .ZN(new_n654_));
  INV_X1    g453(.A(new_n396_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n550_), .A3(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n656_), .A2(new_n658_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n646_), .B1(new_n659_), .B2(new_n660_), .ZN(G1324gat));
  INV_X1    g460(.A(KEYINPUT40), .ZN(new_n662_));
  OAI21_X1  g461(.A(G8gat), .B1(new_n645_), .B2(new_n421_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n654_), .A2(new_n551_), .A3(new_n345_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n662_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n663_), .B(KEYINPUT39), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(KEYINPUT40), .A3(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(G1325gat));
  INV_X1    g470(.A(new_n653_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n203_), .A3(new_n447_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n644_), .A2(new_n447_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n674_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT41), .B1(new_n674_), .B2(G15gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT103), .Z(G1326gat));
  AOI21_X1  g477(.A(new_n411_), .B1(new_n644_), .B2(new_n418_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT42), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n672_), .A2(new_n411_), .A3(new_n418_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1327gat));
  INV_X1    g481(.A(new_n622_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n584_), .A2(new_n683_), .A3(new_n642_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n655_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n583_), .B1(KEYINPUT105), .B2(KEYINPUT44), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(new_n642_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  INV_X1    g487(.A(new_n651_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n451_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n451_), .B2(new_n689_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT105), .B1(new_n693_), .B2(KEYINPUT44), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n694_), .B(new_n687_), .C1(new_n690_), .C2(new_n691_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n396_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n685_), .B1(new_n698_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g498(.A(G36gat), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n642_), .A2(new_n683_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n451_), .A2(new_n700_), .A3(new_n583_), .A4(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(new_n421_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT45), .Z(new_n704_));
  AOI21_X1  g503(.A(new_n421_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(new_n700_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(KEYINPUT46), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT46), .B1(new_n706_), .B2(new_n707_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  NAND2_X1  g509(.A1(new_n696_), .A2(new_n697_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(G43gat), .A3(new_n447_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n684_), .A2(new_n447_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(KEYINPUT107), .A2(G43gat), .ZN(new_n714_));
  OR2_X1    g513(.A1(KEYINPUT107), .A2(G43gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n713_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n712_), .A2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g517(.A1(new_n684_), .A2(new_n543_), .A3(new_n418_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n418_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n721_), .B2(new_n543_), .ZN(G1331gat));
  NOR2_X1   g521(.A1(new_n524_), .A2(new_n581_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n451_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n725_), .A2(new_n624_), .A3(new_n643_), .ZN(new_n726_));
  XOR2_X1   g525(.A(KEYINPUT108), .B(G57gat), .Z(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n655_), .A3(new_n727_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT109), .Z(new_n729_));
  AND2_X1   g528(.A1(new_n724_), .A2(new_n652_), .ZN(new_n730_));
  AOI21_X1  g529(.A(G57gat), .B1(new_n730_), .B2(new_n655_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1332gat));
  INV_X1    g531(.A(G64gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n726_), .B2(new_n345_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT48), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n730_), .A2(new_n733_), .A3(new_n345_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1333gat));
  AOI21_X1  g536(.A(new_n205_), .B1(new_n726_), .B2(new_n447_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT49), .Z(new_n739_));
  NAND3_X1  g538(.A1(new_n730_), .A2(new_n205_), .A3(new_n447_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1334gat));
  INV_X1    g540(.A(G78gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n726_), .B2(new_n418_), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n730_), .A2(new_n742_), .A3(new_n418_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1335gat));
  AND2_X1   g546(.A1(new_n724_), .A2(new_n701_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G85gat), .B1(new_n748_), .B2(new_n655_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n643_), .B(new_n723_), .C1(new_n690_), .C2(new_n691_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT111), .Z(new_n751_));
  NAND3_X1  g550(.A1(new_n655_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT112), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n749_), .B1(new_n751_), .B2(new_n753_), .ZN(G1336gat));
  AOI21_X1  g553(.A(G92gat), .B1(new_n748_), .B2(new_n345_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n751_), .A2(new_n345_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g556(.A(G99gat), .B1(new_n750_), .B2(new_n271_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n476_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n748_), .A2(new_n759_), .A3(new_n447_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g561(.A(G106gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n748_), .A2(new_n763_), .A3(new_n418_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n750_), .A2(new_n720_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G106gat), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n765_), .B(G106gat), .C1(new_n750_), .C2(new_n720_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n772_), .B(new_n764_), .C1(new_n767_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1339gat));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n491_), .A2(KEYINPUT12), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n501_), .B1(new_n598_), .B2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT12), .B1(new_n483_), .B2(new_n496_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n505_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT55), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n505_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n503_), .A2(KEYINPUT114), .A3(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(new_n782_), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n786_), .A3(new_n516_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(new_n514_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n567_), .B1(new_n565_), .B2(new_n569_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(new_n579_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n562_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(KEYINPUT116), .A3(new_n577_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n561_), .A2(new_n567_), .A3(new_n565_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n580_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n785_), .A2(new_n516_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(KEYINPUT56), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT58), .B1(new_n788_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n775_), .B1(new_n651_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(KEYINPUT56), .ZN(new_n801_));
  INV_X1    g600(.A(new_n796_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n801_), .A2(new_n514_), .A3(new_n802_), .A4(new_n787_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n805_), .A2(KEYINPUT117), .A3(new_n649_), .A4(new_n650_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n788_), .A2(new_n798_), .A3(KEYINPUT58), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n800_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n797_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n785_), .A2(KEYINPUT115), .A3(new_n786_), .A4(new_n516_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n512_), .A2(new_n513_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n801_), .A2(new_n810_), .A3(new_n811_), .A4(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n518_), .A2(new_n802_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT57), .B1(new_n815_), .B2(new_n683_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  AOI211_X1 g616(.A(new_n817_), .B(new_n622_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n808_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n643_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n581_), .B1(new_n520_), .B2(new_n523_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n823_), .A2(KEYINPUT113), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(KEYINPUT113), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n652_), .A2(new_n822_), .A3(new_n824_), .A4(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n822_), .A2(new_n651_), .A3(new_n642_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(KEYINPUT113), .A3(new_n823_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n396_), .B1(new_n821_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n448_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n831_), .A2(new_n582_), .A3(new_n271_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n833_));
  OR3_X1    g632(.A1(new_n832_), .A2(new_n833_), .A3(G113gat), .ZN(new_n834_));
  OR3_X1    g633(.A1(new_n831_), .A2(KEYINPUT59), .A3(new_n271_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT59), .B1(new_n831_), .B2(new_n271_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n835_), .A2(G113gat), .A3(new_n581_), .A4(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n833_), .B1(new_n832_), .B2(G113gat), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n834_), .A2(new_n837_), .A3(new_n838_), .ZN(G1340gat));
  NOR2_X1   g638(.A1(new_n831_), .A2(new_n271_), .ZN(new_n840_));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n524_), .B2(KEYINPUT60), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n841_), .A2(KEYINPUT60), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT119), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n835_), .A2(new_n525_), .A3(new_n836_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G120gat), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1341gat));
  AOI21_X1  g647(.A(G127gat), .B1(new_n840_), .B2(new_n642_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n835_), .A2(new_n836_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n642_), .A2(G127gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT120), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n849_), .B1(new_n850_), .B2(new_n852_), .ZN(G1342gat));
  AOI21_X1  g652(.A(G134gat), .B1(new_n840_), .B2(new_n624_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n689_), .A2(G134gat), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n855_), .B(KEYINPUT121), .Z(new_n856_));
  AOI21_X1  g655(.A(new_n854_), .B1(new_n850_), .B2(new_n856_), .ZN(G1343gat));
  AOI21_X1  g656(.A(new_n642_), .B1(new_n808_), .B2(new_n819_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n826_), .A2(new_n828_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n655_), .B(new_n271_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n345_), .A2(new_n720_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n581_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n525_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT122), .B(G148gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1345gat));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n863_), .B2(new_n642_), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n860_), .A2(KEYINPUT123), .A3(new_n643_), .A4(new_n862_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT61), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n830_), .A2(new_n271_), .A3(new_n642_), .A4(new_n861_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT123), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n863_), .A2(new_n869_), .A3(new_n642_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT61), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n872_), .A2(G155gat), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(G155gat), .B1(new_n872_), .B2(new_n877_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1346gat));
  AOI21_X1  g679(.A(G162gat), .B1(new_n863_), .B2(new_n624_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n651_), .A2(new_n610_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n863_), .B2(new_n882_), .ZN(G1347gat));
  NAND2_X1  g682(.A1(new_n821_), .A2(new_n829_), .ZN(new_n884_));
  NOR4_X1   g683(.A1(new_n271_), .A2(new_n655_), .A3(new_n418_), .A4(new_n421_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n581_), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n884_), .A2(KEYINPUT124), .A3(new_n581_), .A4(new_n885_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(G169gat), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT125), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n888_), .A2(new_n892_), .A3(G169gat), .A4(new_n889_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n891_), .A2(KEYINPUT62), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n890_), .A2(KEYINPUT125), .A3(new_n895_), .ZN(new_n896_));
  XOR2_X1   g695(.A(KEYINPUT22), .B(G169gat), .Z(new_n897_));
  OAI211_X1 g696(.A(new_n894_), .B(new_n896_), .C1(new_n886_), .C2(new_n897_), .ZN(G1348gat));
  AND2_X1   g697(.A1(new_n884_), .A2(new_n885_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n525_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n642_), .ZN(new_n902_));
  MUX2_X1   g701(.A(new_n231_), .B(G183gat), .S(new_n902_), .Z(G1350gat));
  NAND2_X1  g702(.A1(new_n899_), .A2(new_n689_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(G190gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n899_), .A2(new_n234_), .A3(new_n624_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1351gat));
  NOR2_X1   g706(.A1(new_n447_), .A2(new_n421_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n884_), .A2(new_n396_), .A3(new_n418_), .A4(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n582_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(new_n289_), .ZN(G1352gat));
  INV_X1    g710(.A(new_n909_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n525_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G204gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n914_), .B1(new_n291_), .B2(new_n913_), .ZN(G1353gat));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n916_));
  INV_X1    g715(.A(G211gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n642_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT126), .Z(new_n919_));
  OR3_X1    g718(.A1(new_n909_), .A2(KEYINPUT127), .A3(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT127), .B1(new_n909_), .B2(new_n919_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n916_), .A2(new_n917_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1354gat));
  INV_X1    g723(.A(G218gat), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n909_), .A2(new_n925_), .A3(new_n651_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n912_), .A2(new_n624_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n926_), .B1(new_n925_), .B2(new_n927_), .ZN(G1355gat));
endmodule


