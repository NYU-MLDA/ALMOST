//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT24), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT24), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n206_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT84), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT84), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G183gat), .A3(G190gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT23), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n210_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT26), .B(G190gat), .ZN(new_n219_));
  INV_X1    g018(.A(G183gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT25), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G183gat), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n221_), .A2(new_n223_), .A3(KEYINPUT92), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT92), .B1(new_n221_), .B2(new_n223_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n219_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n218_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(G169gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n204_), .A2(KEYINPUT22), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT93), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n204_), .A2(KEYINPUT22), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(G169gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT93), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n231_), .A2(new_n205_), .A3(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n212_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n237_));
  INV_X1    g036(.A(G190gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n220_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n236_), .A2(new_n207_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n227_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G211gat), .B(G218gat), .ZN(new_n244_));
  INV_X1    g043(.A(G197gat), .ZN(new_n245_));
  INV_X1    g044(.A(G204gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G197gat), .A2(G204gat), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(KEYINPUT21), .B(new_n244_), .C1(new_n249_), .C2(KEYINPUT89), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT21), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT89), .B1(new_n247_), .B2(new_n248_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G211gat), .B(G218gat), .Z(new_n253_));
  OAI21_X1  g052(.A(new_n251_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n247_), .A2(new_n248_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n250_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n243_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n210_), .ZN(new_n260_));
  OR3_X1    g059(.A1(new_n220_), .A2(KEYINPUT83), .A3(KEYINPUT25), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT25), .B1(new_n220_), .B2(KEYINPUT83), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n219_), .A3(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n260_), .A2(new_n263_), .A3(new_n237_), .A4(new_n240_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n215_), .A2(new_n217_), .B1(new_n220_), .B2(new_n238_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT22), .B(G169gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT85), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n266_), .A2(new_n267_), .A3(new_n205_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n267_), .B1(new_n266_), .B2(new_n205_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n207_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n257_), .B(new_n264_), .C1(new_n265_), .C2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n259_), .A2(KEYINPUT20), .A3(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G226gat), .A2(G233gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G8gat), .B(G36gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT18), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT95), .ZN(new_n280_));
  XOR2_X1   g079(.A(G64gat), .B(G92gat), .Z(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n264_), .B1(new_n270_), .B2(new_n265_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(new_n258_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n257_), .A2(new_n227_), .A3(new_n242_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n285_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n277_), .B(new_n282_), .C1(new_n276_), .C2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT100), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n281_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n280_), .B(new_n290_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n276_), .A4(new_n285_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT20), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n243_), .B2(new_n258_), .ZN(new_n294_));
  AOI211_X1 g093(.A(KEYINPUT94), .B(new_n276_), .C1(new_n294_), .C2(new_n271_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT94), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n291_), .B(new_n292_), .C1(new_n295_), .C2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT27), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n289_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n292_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n272_), .A2(new_n275_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT94), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n272_), .A2(new_n296_), .A3(new_n275_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n302_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT96), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(new_n291_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n292_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT96), .B1(new_n309_), .B2(new_n282_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n298_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n308_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n301_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT87), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT87), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G155gat), .A3(G162gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n319_), .A3(KEYINPUT1), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT1), .B1(new_n317_), .B2(new_n319_), .ZN(new_n322_));
  OAI22_X1  g121(.A1(new_n321_), .A2(new_n322_), .B1(G155gat), .B2(G162gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G141gat), .A2(G148gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G141gat), .A2(G148gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(KEYINPUT88), .A2(KEYINPUT3), .ZN(new_n328_));
  NOR2_X1   g127(.A1(KEYINPUT88), .A2(KEYINPUT3), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n328_), .B1(new_n326_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(KEYINPUT2), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G141gat), .A3(G148gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(KEYINPUT88), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n330_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n337_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n323_), .A2(new_n327_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT29), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n258_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G228gat), .A2(G233gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n258_), .B(new_n342_), .C1(new_n339_), .C2(new_n340_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G78gat), .B(G106gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n344_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT90), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT28), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n339_), .A2(new_n350_), .A3(new_n340_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n336_), .A2(new_n338_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n318_), .B1(G155gat), .B2(G162gat), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n316_), .A2(KEYINPUT87), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n337_), .B1(new_n356_), .B2(new_n320_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n327_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n352_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT28), .B1(new_n359_), .B2(KEYINPUT29), .ZN(new_n360_));
  XOR2_X1   g159(.A(G22gat), .B(G50gat), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n351_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n362_), .B1(new_n351_), .B2(new_n360_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n348_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n347_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n349_), .B(new_n366_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n344_), .A2(new_n345_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n346_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n365_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n363_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n371_), .B(new_n348_), .C1(new_n373_), .C2(KEYINPUT90), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n369_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n315_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G127gat), .B(G134gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G113gat), .B(G120gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n359_), .A2(new_n380_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n352_), .B(new_n379_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(KEYINPUT4), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n359_), .A2(new_n384_), .A3(new_n380_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT97), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n383_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT0), .ZN(new_n390_));
  INV_X1    g189(.A(G57gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G85gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n381_), .A2(new_n382_), .A3(new_n386_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n388_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n388_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT99), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n388_), .A2(new_n394_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n393_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT99), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n388_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n397_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n283_), .B(KEYINPUT30), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(G15gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G71gat), .B(G99gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(KEYINPUT86), .B(G43gat), .Z(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n405_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT31), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n413_), .A2(new_n379_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n379_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n376_), .A2(new_n404_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n289_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n419_));
  AND4_X1   g218(.A1(new_n397_), .A2(new_n403_), .A3(new_n369_), .A4(new_n374_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n298_), .A2(KEYINPUT96), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n307_), .B1(new_n306_), .B2(new_n291_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(new_n298_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n419_), .B(new_n420_), .C1(new_n423_), .C2(new_n313_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT102), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n312_), .A2(new_n314_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT102), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n419_), .A4(new_n420_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n291_), .A2(KEYINPUT32), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n429_), .B(new_n277_), .C1(new_n276_), .C2(new_n286_), .ZN(new_n430_));
  OAI221_X1 g229(.A(new_n430_), .B1(new_n396_), .B2(new_n395_), .C1(new_n309_), .C2(new_n429_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT33), .B1(new_n395_), .B2(KEYINPUT98), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n383_), .A2(new_n386_), .A3(new_n385_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n381_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n399_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT98), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT33), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n402_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n432_), .A2(new_n435_), .A3(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n431_), .B1(new_n312_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n375_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n425_), .A2(new_n428_), .A3(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n442_), .A2(KEYINPUT103), .A3(new_n416_), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT103), .B1(new_n442_), .B2(new_n416_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n418_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G230gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G57gat), .B(G64gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT11), .ZN(new_n448_));
  XOR2_X1   g247(.A(G71gat), .B(G78gat), .Z(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n449_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n447_), .A2(KEYINPUT11), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G99gat), .A2(G106gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT6), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n457_));
  OR3_X1    g256(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G85gat), .B(G92gat), .Z(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(KEYINPUT8), .A3(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(KEYINPUT10), .B(G99gat), .Z(new_n462_));
  INV_X1    g261(.A(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n460_), .A2(KEYINPUT9), .ZN(new_n465_));
  INV_X1    g264(.A(G85gat), .ZN(new_n466_));
  INV_X1    g265(.A(G92gat), .ZN(new_n467_));
  OR3_X1    g266(.A1(new_n466_), .A2(new_n467_), .A3(KEYINPUT9), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n464_), .A2(new_n465_), .A3(new_n456_), .A4(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n461_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT8), .B1(new_n459_), .B2(new_n460_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n472_), .A2(KEYINPUT64), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(KEYINPUT64), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n454_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT66), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n473_), .A2(new_n454_), .A3(new_n474_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT65), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n446_), .B1(new_n476_), .B2(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n475_), .A2(KEYINPUT12), .ZN(new_n481_));
  INV_X1    g280(.A(new_n472_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n454_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(KEYINPUT12), .A3(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n477_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n446_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G120gat), .B(G148gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT5), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT67), .ZN(new_n491_));
  XOR2_X1   g290(.A(G176gat), .B(G204gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n480_), .A2(new_n488_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n480_), .B2(new_n488_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT13), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n496_), .A2(new_n497_), .A3(KEYINPUT13), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(G8gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT74), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n504_), .A2(new_n505_), .ZN(new_n507_));
  XOR2_X1   g306(.A(G15gat), .B(G22gat), .Z(new_n508_));
  NOR3_X1   g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G1gat), .B(G8gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G29gat), .B(G36gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G43gat), .B(G50gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n511_), .B(new_n514_), .Z(new_n515_));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n514_), .B(KEYINPUT15), .ZN(new_n518_));
  MUX2_X1   g317(.A(new_n514_), .B(new_n518_), .S(new_n511_), .Z(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G113gat), .B(G141gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT82), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G169gat), .B(G197gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT81), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n520_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n502_), .A2(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n445_), .A2(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G190gat), .B(G218gat), .Z(new_n530_));
  XNOR2_X1  g329(.A(G134gat), .B(G162gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT36), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n533_), .B(KEYINPUT70), .Z(new_n534_));
  AND2_X1   g333(.A1(new_n473_), .A2(new_n474_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n514_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n482_), .A2(new_n518_), .B1(new_n541_), .B2(new_n540_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n536_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n543_), .B1(new_n536_), .B2(new_n544_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n534_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT71), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT71), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n550_), .B(new_n534_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n547_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n532_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(KEYINPUT36), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n545_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G127gat), .B(G155gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT16), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT75), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G183gat), .B(G211gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT77), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n511_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(new_n483_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT78), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT79), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n572_), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n563_), .B(KEYINPUT17), .Z(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n558_), .A2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n529_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n202_), .B1(new_n579_), .B2(new_n404_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT104), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT73), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT37), .ZN(new_n583_));
  INV_X1    g382(.A(new_n555_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n546_), .A2(new_n547_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT69), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT69), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n556_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n583_), .B1(new_n589_), .B2(new_n548_), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT72), .B(KEYINPUT37), .Z(new_n591_));
  AOI211_X1 g390(.A(new_n585_), .B(new_n591_), .C1(new_n549_), .C2(new_n551_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n582_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n591_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n552_), .A2(new_n556_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n548_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n595_), .B(KEYINPUT73), .C1(new_n583_), .C2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n577_), .B1(new_n593_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n502_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT80), .Z(new_n602_));
  NAND2_X1  g401(.A1(new_n441_), .A2(new_n428_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n427_), .B1(new_n315_), .B2(new_n420_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n416_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT103), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n442_), .A2(KEYINPUT103), .A3(new_n416_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n417_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n602_), .A2(new_n609_), .A3(new_n527_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n404_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(G1gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(KEYINPUT38), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT38), .ZN(new_n614_));
  INV_X1    g413(.A(new_n610_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n612_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n614_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n617_), .A2(KEYINPUT105), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(KEYINPUT105), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n581_), .B(new_n613_), .C1(new_n618_), .C2(new_n619_), .ZN(G1324gat));
  NOR2_X1   g419(.A1(new_n315_), .A2(G8gat), .ZN(new_n621_));
  INV_X1    g420(.A(new_n315_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n579_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(G8gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n610_), .A2(new_n621_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n624_), .A2(new_n625_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(G1325gat));
  INV_X1    g429(.A(new_n416_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n579_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(G15gat), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n633_), .A2(KEYINPUT41), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(KEYINPUT41), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n416_), .A2(G15gat), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n634_), .B(new_n635_), .C1(new_n615_), .C2(new_n636_), .ZN(G1326gat));
  INV_X1    g436(.A(G22gat), .ZN(new_n638_));
  INV_X1    g437(.A(new_n375_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n579_), .B2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT42), .Z(new_n641_));
  NAND3_X1  g440(.A1(new_n610_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1327gat));
  NAND2_X1  g442(.A1(new_n558_), .A2(new_n577_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n529_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(G29gat), .B1(new_n646_), .B2(new_n404_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n500_), .A2(new_n577_), .A3(new_n526_), .A4(new_n501_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT107), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n593_), .A2(new_n598_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n609_), .A2(KEYINPUT43), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT43), .ZN(new_n652_));
  INV_X1    g451(.A(new_n650_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n445_), .B2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(KEYINPUT44), .B(new_n649_), .C1(new_n651_), .C2(new_n654_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n655_), .A2(G29gat), .A3(new_n404_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n651_), .A2(new_n654_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n649_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n657_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n647_), .B1(new_n656_), .B2(new_n660_), .ZN(G1328gat));
  INV_X1    g460(.A(KEYINPUT109), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(KEYINPUT46), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT110), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n655_), .A2(new_n622_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT43), .B1(new_n609_), .B2(new_n650_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n445_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT44), .B1(new_n669_), .B2(new_n649_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G36gat), .B1(new_n666_), .B2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n315_), .A2(G36gat), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n445_), .A2(new_n528_), .A3(new_n645_), .A4(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n662_), .A2(KEYINPUT46), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n665_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n678_), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT110), .B(new_n680_), .C1(new_n671_), .C2(new_n676_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n664_), .B1(new_n679_), .B2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n660_), .A2(new_n622_), .A3(new_n655_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n675_), .B1(new_n683_), .B2(G36gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT110), .B1(new_n684_), .B2(new_n680_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n677_), .A2(new_n665_), .A3(new_n678_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n663_), .A3(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n682_), .A2(new_n687_), .ZN(G1329gat));
  NAND2_X1  g487(.A1(new_n660_), .A2(new_n655_), .ZN(new_n689_));
  INV_X1    g488(.A(G43gat), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n416_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G43gat), .B1(new_n646_), .B2(new_n631_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(G1330gat));
  OAI21_X1  g494(.A(G50gat), .B1(new_n689_), .B2(new_n375_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n375_), .A2(G50gat), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT112), .Z(new_n698_));
  NAND2_X1  g497(.A1(new_n646_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(G1331gat));
  NOR2_X1   g499(.A1(new_n600_), .A2(new_n526_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n445_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n599_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n611_), .B1(new_n703_), .B2(KEYINPUT113), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n704_), .B1(KEYINPUT113), .B2(new_n703_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n702_), .A2(new_n578_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n611_), .A2(new_n391_), .ZN(new_n707_));
  AOI22_X1  g506(.A1(new_n705_), .A2(new_n391_), .B1(new_n706_), .B2(new_n707_), .ZN(G1332gat));
  INV_X1    g507(.A(G64gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n706_), .B2(new_n622_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT48), .Z(new_n711_));
  NAND2_X1  g510(.A1(new_n622_), .A2(new_n709_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n703_), .B2(new_n712_), .ZN(G1333gat));
  INV_X1    g512(.A(new_n706_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G71gat), .B1(new_n714_), .B2(new_n416_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT49), .ZN(new_n716_));
  OR3_X1    g515(.A1(new_n703_), .A2(G71gat), .A3(new_n416_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT114), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n716_), .A2(KEYINPUT114), .A3(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1334gat));
  OAI21_X1  g521(.A(G78gat), .B1(new_n714_), .B2(new_n375_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT50), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n375_), .A2(G78gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n703_), .B2(new_n725_), .ZN(G1335gat));
  AND2_X1   g525(.A1(new_n702_), .A2(new_n645_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(new_n466_), .A3(new_n404_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n669_), .A2(new_n577_), .A3(new_n701_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(new_n404_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n728_), .B1(new_n730_), .B2(new_n466_), .ZN(G1336gat));
  NAND3_X1  g530(.A1(new_n727_), .A2(new_n467_), .A3(new_n622_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n729_), .A2(new_n622_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n467_), .ZN(G1337gat));
  NAND3_X1  g533(.A1(new_n727_), .A2(new_n462_), .A3(new_n631_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(KEYINPUT115), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n729_), .A2(new_n631_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(G99gat), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(KEYINPUT115), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n739_), .B(new_n740_), .Z(G1338gat));
  AOI21_X1  g540(.A(new_n463_), .B1(new_n729_), .B2(new_n639_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n743_));
  OR2_X1    g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n743_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n727_), .A2(new_n463_), .A3(new_n639_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT116), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(new_n745_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT53), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n744_), .A2(new_n750_), .A3(new_n745_), .A4(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1339gat));
  INV_X1    g551(.A(KEYINPUT120), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n524_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n754_), .A2(KEYINPUT119), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n519_), .A2(new_n516_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n754_), .B2(KEYINPUT119), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n524_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n520_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n753_), .B1(new_n498_), .B2(new_n761_), .ZN(new_n762_));
  AOI211_X1 g561(.A(KEYINPUT120), .B(new_n760_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n481_), .A2(new_n485_), .A3(KEYINPUT55), .A4(new_n446_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n486_), .A2(new_n487_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT56), .B1(new_n769_), .B2(new_n494_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n494_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n769_), .A2(new_n771_), .A3(KEYINPUT56), .A4(new_n494_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n527_), .A2(new_n495_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n764_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n557_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT121), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n770_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n773_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n495_), .A2(new_n760_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT58), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT122), .B1(new_n650_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n785_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT58), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT122), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n593_), .A4(new_n598_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n784_), .A2(KEYINPUT58), .A3(new_n785_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n787_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n558_), .B1(new_n764_), .B2(new_n777_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT121), .B1(new_n795_), .B2(KEYINPUT57), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(KEYINPUT57), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n782_), .A2(new_n794_), .A3(new_n796_), .A4(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n577_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n599_), .A2(new_n527_), .A3(new_n600_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT54), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n376_), .A2(new_n611_), .A3(new_n416_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT59), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n779_), .A2(new_n781_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n794_), .A2(new_n806_), .A3(new_n797_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n577_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n801_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n803_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n805_), .A2(new_n526_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G113gat), .ZN(new_n813_));
  OR3_X1    g612(.A1(new_n804_), .A2(G113gat), .A3(new_n527_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1340gat));
  NAND3_X1  g614(.A1(new_n805_), .A2(new_n502_), .A3(new_n811_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(G120gat), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n600_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(KEYINPUT60), .B2(G120gat), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n804_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n817_), .A2(new_n820_), .ZN(G1341gat));
  NAND3_X1  g620(.A1(new_n805_), .A2(new_n808_), .A3(new_n811_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(G127gat), .ZN(new_n823_));
  OR3_X1    g622(.A1(new_n804_), .A2(G127gat), .A3(new_n577_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(G1342gat));
  AND2_X1   g624(.A1(new_n805_), .A2(new_n811_), .ZN(new_n826_));
  XOR2_X1   g625(.A(KEYINPUT123), .B(G134gat), .Z(new_n827_));
  NOR2_X1   g626(.A1(new_n650_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(G134gat), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n802_), .A2(new_n558_), .A3(new_n803_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n826_), .A2(new_n828_), .B1(new_n829_), .B2(new_n830_), .ZN(G1343gat));
  NOR4_X1   g630(.A1(new_n631_), .A2(new_n622_), .A3(new_n611_), .A4(new_n375_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n802_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n526_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n502_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g637(.A1(new_n833_), .A2(new_n577_), .ZN(new_n839_));
  XOR2_X1   g638(.A(KEYINPUT61), .B(G155gat), .Z(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1346gat));
  OR3_X1    g640(.A1(new_n833_), .A2(G162gat), .A3(new_n557_), .ZN(new_n842_));
  OAI21_X1  g641(.A(G162gat), .B1(new_n833_), .B2(new_n650_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1347gat));
  NOR3_X1   g643(.A1(new_n416_), .A2(new_n315_), .A3(new_n404_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(new_n639_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n809_), .A2(new_n526_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(G169gat), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT124), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(G169gat), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT62), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n848_), .A2(new_n854_), .A3(new_n849_), .A4(G169gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n851_), .A2(new_n853_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n809_), .A2(new_n847_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n526_), .A2(new_n231_), .A3(new_n235_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT125), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n856_), .A2(new_n861_), .ZN(G1348gat));
  AOI21_X1  g661(.A(G176gat), .B1(new_n858_), .B2(new_n502_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n800_), .B(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n798_), .B2(new_n577_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n639_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n600_), .A2(new_n205_), .A3(new_n846_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n863_), .B1(new_n867_), .B2(new_n868_), .ZN(G1349gat));
  NAND3_X1  g668(.A1(new_n867_), .A2(new_n808_), .A3(new_n845_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n577_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n870_), .A2(new_n220_), .B1(new_n858_), .B2(new_n871_), .ZN(G1350gat));
  OAI21_X1  g671(.A(G190gat), .B1(new_n857_), .B2(new_n650_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n558_), .A2(new_n219_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n857_), .B2(new_n874_), .ZN(G1351gat));
  NOR2_X1   g674(.A1(new_n631_), .A2(new_n375_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n611_), .A3(new_n622_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n802_), .A2(KEYINPUT126), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT126), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n866_), .B2(new_n877_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(G197gat), .B1(new_n882_), .B2(new_n526_), .ZN(new_n883_));
  AOI211_X1 g682(.A(new_n245_), .B(new_n527_), .C1(new_n879_), .C2(new_n881_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1352gat));
  AND2_X1   g684(.A1(new_n879_), .A2(new_n881_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G204gat), .B1(new_n886_), .B2(new_n600_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n882_), .A2(new_n246_), .A3(new_n502_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1353gat));
  NOR2_X1   g688(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(KEYINPUT127), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n577_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n882_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n892_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n891_), .ZN(new_n895_));
  AOI211_X1 g694(.A(new_n894_), .B(new_n895_), .C1(new_n879_), .C2(new_n881_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n893_), .A2(new_n896_), .ZN(G1354gat));
  OAI21_X1  g696(.A(G218gat), .B1(new_n886_), .B2(new_n650_), .ZN(new_n898_));
  INV_X1    g697(.A(G218gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n882_), .A2(new_n899_), .A3(new_n558_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1355gat));
endmodule


