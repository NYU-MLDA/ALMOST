//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G29gat), .B(G36gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT77), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT77), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n206_), .B(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(new_n208_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n205_), .B1(new_n210_), .B2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G1gat), .B(G8gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT80), .B(G8gat), .ZN(new_n216_));
  INV_X1    g015(.A(G1gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT14), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n215_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n218_), .A2(new_n219_), .A3(new_n215_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n212_), .A2(new_n208_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n207_), .A2(new_n209_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(KEYINPUT15), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n214_), .A2(new_n223_), .A3(new_n226_), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n224_), .A2(new_n225_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n230_), .B(KEYINPUT83), .Z(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n221_), .A2(new_n222_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n224_), .A2(new_n225_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(G229gat), .B(G233gat), .C1(new_n235_), .C2(new_n228_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n204_), .B1(new_n237_), .B2(KEYINPUT84), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT84), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n232_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(KEYINPUT85), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n204_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n237_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT85), .B1(new_n238_), .B2(new_n240_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(KEYINPUT86), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT86), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n241_), .A2(new_n244_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(new_n250_), .B2(new_n246_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G127gat), .B(G134gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G113gat), .B(G120gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT93), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G141gat), .A2(G148gat), .ZN(new_n258_));
  INV_X1    g057(.A(G141gat), .ZN(new_n259_));
  INV_X1    g058(.A(G148gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT94), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT1), .ZN(new_n264_));
  OR2_X1    g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n264_), .B(new_n265_), .C1(KEYINPUT1), .C2(new_n262_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n263_), .B1(new_n262_), .B2(KEYINPUT1), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n258_), .B(new_n261_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT95), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT3), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(new_n259_), .A4(new_n260_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n258_), .A2(new_n272_), .ZN(new_n273_));
  OAI22_X1  g072(.A1(KEYINPUT95), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n271_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  OAI22_X1  g074(.A1(new_n258_), .A2(new_n272_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n262_), .B(new_n265_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n268_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n257_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n279_), .B2(new_n256_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G225gat), .A2(G233gat), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT105), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(KEYINPUT104), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT93), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n256_), .B(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(new_n284_), .A3(new_n278_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT104), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n282_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n279_), .A2(new_n256_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n292_), .B(KEYINPUT4), .C1(new_n257_), .C2(new_n279_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n285_), .A2(new_n290_), .A3(new_n291_), .A4(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n283_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n288_), .B(KEYINPUT104), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n296_), .A2(KEYINPUT105), .A3(new_n291_), .A4(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G1gat), .B(G29gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(G85gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT0), .B(G57gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  NAND2_X1  g101(.A1(new_n298_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT106), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT33), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n302_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT106), .B1(new_n308_), .B2(KEYINPUT33), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT103), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G8gat), .B(G36gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT18), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G64gat), .B(G92gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n313_), .B(new_n314_), .Z(new_n315_));
  INV_X1    g114(.A(KEYINPUT20), .ZN(new_n316_));
  XOR2_X1   g115(.A(KEYINPUT90), .B(G176gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT22), .B(G169gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT91), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n320_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT91), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT89), .B(KEYINPUT23), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G183gat), .A2(G190gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n329_), .A2(KEYINPUT23), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n322_), .B(new_n325_), .C1(new_n326_), .C2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT88), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n336_), .A2(KEYINPUT24), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n328_), .A2(KEYINPUT23), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n338_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(KEYINPUT24), .A3(new_n320_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT25), .B(G183gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT26), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT87), .B1(new_n343_), .B2(G190gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT26), .B(G190gat), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n342_), .B(new_n344_), .C1(new_n345_), .C2(KEYINPUT87), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n340_), .A2(new_n341_), .A3(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n333_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G211gat), .B(G218gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT96), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G197gat), .B(G204gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT21), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n350_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n352_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n350_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n316_), .B1(new_n348_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n337_), .A2(new_n332_), .A3(KEYINPUT102), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT102), .B1(new_n337_), .B2(new_n332_), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n345_), .B(KEYINPUT101), .Z(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n342_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n363_), .A2(new_n364_), .A3(new_n341_), .A4(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n321_), .B1(new_n339_), .B2(new_n326_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n358_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n360_), .A2(new_n362_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n369_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n359_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n333_), .A2(new_n347_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n316_), .B1(new_n374_), .B2(new_n358_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n362_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n311_), .B(new_n315_), .C1(new_n371_), .C2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n373_), .A2(new_n375_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n362_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n360_), .A2(new_n362_), .A3(new_n370_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n315_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n377_), .A2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n315_), .B1(new_n371_), .B2(new_n376_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT103), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n308_), .A2(KEYINPUT33), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n296_), .A2(new_n282_), .A3(new_n293_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n302_), .B1(new_n281_), .B2(new_n291_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n384_), .A2(new_n386_), .A3(new_n387_), .A4(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n295_), .A2(new_n297_), .A3(new_n307_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(new_n308_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n380_), .A2(new_n381_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n315_), .A2(KEYINPUT32), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n360_), .A2(new_n379_), .A3(new_n370_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n358_), .B(KEYINPUT98), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n372_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n379_), .B1(new_n400_), .B2(new_n375_), .ZN(new_n401_));
  OAI211_X1 g200(.A(KEYINPUT32), .B(new_n315_), .C1(new_n398_), .C2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n397_), .A2(new_n402_), .ZN(new_n403_));
  OAI22_X1  g202(.A1(new_n310_), .A2(new_n391_), .B1(new_n394_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n278_), .A2(KEYINPUT29), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G228gat), .A2(G233gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n359_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n406_), .A2(KEYINPUT97), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n406_), .A2(KEYINPUT97), .ZN(new_n411_));
  OR3_X1    g210(.A1(new_n399_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n409_), .B1(new_n412_), .B2(new_n408_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n414_), .B(KEYINPUT99), .Z(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT100), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G22gat), .B(G50gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n278_), .A2(KEYINPUT29), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n419_), .A2(KEYINPUT28), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(KEYINPUT28), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n418_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n421_), .A3(new_n418_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n416_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n426_), .A2(new_n415_), .A3(new_n422_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n413_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  OAI22_X1  g227(.A1(new_n426_), .A2(new_n422_), .B1(KEYINPUT100), .B2(new_n415_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n415_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n423_), .A2(new_n430_), .A3(new_n424_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n399_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n432_), .A2(new_n407_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n429_), .B(new_n431_), .C1(new_n433_), .C2(new_n409_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n428_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G227gat), .A2(G233gat), .ZN(new_n437_));
  INV_X1    g236(.A(G71gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G15gat), .B(G43gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT92), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n441_), .B(KEYINPUT30), .Z(new_n442_));
  NAND2_X1  g241(.A1(new_n374_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n374_), .A2(new_n442_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n439_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n445_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n439_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n443_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n287_), .B(KEYINPUT31), .ZN(new_n451_));
  INV_X1    g250(.A(G99gat), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n452_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n446_), .A2(new_n449_), .A3(new_n453_), .A4(new_n454_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n436_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n404_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n386_), .A2(new_n377_), .A3(new_n383_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT27), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n382_), .B1(new_n398_), .B2(new_n401_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n463_), .B1(new_n395_), .B2(new_n315_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n462_), .A2(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n435_), .A2(new_n459_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n458_), .A2(new_n428_), .A3(new_n434_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT107), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(new_n393_), .B2(new_n308_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n303_), .A2(KEYINPUT107), .A3(new_n392_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n466_), .A2(new_n469_), .A3(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n253_), .B1(new_n461_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G230gat), .A2(G233gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(G85gat), .B2(G92gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT64), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT64), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n481_), .B1(new_n482_), .B2(new_n478_), .ZN(new_n483_));
  XOR2_X1   g282(.A(KEYINPUT10), .B(G99gat), .Z(new_n484_));
  INV_X1    g283(.A(G106gat), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n480_), .A2(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT65), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(KEYINPUT6), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(KEYINPUT65), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n488_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(KEYINPUT65), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n489_), .A2(KEYINPUT6), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n487_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n493_), .A2(KEYINPUT66), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT66), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n494_), .A2(new_n495_), .A3(new_n487_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n487_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n486_), .A2(new_n497_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT70), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n504_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n493_), .A2(KEYINPUT70), .A3(new_n496_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT67), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT7), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT7), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT67), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n508_), .A2(new_n510_), .B1(new_n452_), .B2(new_n485_), .ZN(new_n511_));
  AOI211_X1 g310(.A(G99gat), .B(G106gat), .C1(new_n507_), .C2(KEYINPUT7), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n505_), .A2(new_n506_), .A3(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G85gat), .B(G92gat), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n515_), .A2(KEYINPUT69), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(KEYINPUT69), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT8), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n501_), .A2(new_n497_), .A3(new_n513_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT68), .B(KEYINPUT8), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n503_), .B1(new_n520_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT72), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G57gat), .B(G64gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT11), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT71), .B(G71gat), .ZN(new_n529_));
  INV_X1    g328(.A(G78gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n529_), .B(G78gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n527_), .A2(KEYINPUT11), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n525_), .A2(new_n526_), .A3(new_n537_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n521_), .A2(new_n523_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT8), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n540_), .B1(new_n514_), .B2(new_n518_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n537_), .B(new_n502_), .C1(new_n539_), .C2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT72), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n525_), .A2(new_n537_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n477_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n477_), .B1(new_n525_), .B2(new_n537_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n502_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT12), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n536_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n549_), .B1(new_n548_), .B2(new_n536_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n547_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n546_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT73), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT73), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n546_), .A2(new_n555_), .A3(new_n552_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G120gat), .B(G148gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT5), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G176gat), .B(G204gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT74), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n554_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n546_), .A2(new_n552_), .A3(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT13), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT75), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n565_), .B(KEYINPUT13), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT75), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n548_), .A2(new_n226_), .A3(new_n214_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n525_), .A2(new_n234_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT76), .B(KEYINPUT34), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT35), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n572_), .A2(new_n573_), .A3(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n577_), .A2(new_n578_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n581_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n572_), .A2(new_n573_), .A3(new_n583_), .A4(new_n579_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G190gat), .B(G218gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT78), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n585_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT37), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n589_), .B(KEYINPUT36), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n585_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n595_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT79), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n585_), .B2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n582_), .A2(KEYINPUT79), .A3(new_n584_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n592_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n597_), .B1(new_n602_), .B2(KEYINPUT37), .ZN(new_n603_));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT16), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT81), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n536_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(new_n233_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n607_), .B1(new_n612_), .B2(KEYINPUT17), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(KEYINPUT82), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n607_), .A2(KEYINPUT17), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n614_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n603_), .A2(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n475_), .A2(new_n569_), .A3(new_n571_), .A4(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n621_), .A2(G1gat), .A3(new_n473_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT38), .Z(new_n623_));
  NAND2_X1  g422(.A1(new_n245_), .A2(new_n247_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n569_), .A2(new_n571_), .A3(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n394_), .A2(new_n403_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n386_), .A2(new_n377_), .A3(new_n383_), .A4(new_n390_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n387_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n306_), .A2(new_n309_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n460_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n474_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n602_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n618_), .A3(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n625_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n473_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n217_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT108), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n623_), .A2(new_n639_), .ZN(G1324gat));
  XNOR2_X1  g439(.A(KEYINPUT111), .B(KEYINPUT40), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT112), .ZN(new_n643_));
  INV_X1    g442(.A(G8gat), .ZN(new_n644_));
  INV_X1    g443(.A(new_n466_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n636_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT110), .B(KEYINPUT39), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n216_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT109), .B1(new_n621_), .B2(new_n649_), .ZN(new_n650_));
  AND4_X1   g449(.A1(new_n569_), .A2(new_n633_), .A3(new_n571_), .A4(new_n252_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT109), .ZN(new_n652_));
  INV_X1    g451(.A(new_n649_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n620_), .A4(new_n653_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n646_), .A2(new_n648_), .B1(new_n650_), .B2(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n625_), .A2(new_n635_), .A3(new_n466_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n647_), .B1(new_n656_), .B2(new_n644_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n643_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n650_), .A2(new_n654_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n625_), .A2(new_n635_), .ZN(new_n660_));
  OAI211_X1 g459(.A(G8gat), .B(new_n648_), .C1(new_n660_), .C2(new_n466_), .ZN(new_n661_));
  AND4_X1   g460(.A1(new_n643_), .A2(new_n659_), .A3(new_n661_), .A4(new_n657_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n642_), .B1(new_n658_), .B2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(new_n661_), .A3(new_n657_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT112), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n655_), .A2(new_n643_), .A3(new_n657_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n666_), .A3(new_n641_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n667_), .ZN(G1325gat));
  OAI21_X1  g467(.A(G15gat), .B1(new_n660_), .B2(new_n458_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT41), .Z(new_n670_));
  NOR3_X1   g469(.A1(new_n621_), .A2(G15gat), .A3(new_n458_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT113), .Z(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1326gat));
  OAI21_X1  g472(.A(G22gat), .B1(new_n660_), .B2(new_n435_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT42), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n435_), .A2(G22gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n621_), .B2(new_n676_), .ZN(G1327gat));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n603_), .A2(KEYINPUT114), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n603_), .A2(KEYINPUT114), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n633_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n603_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(KEYINPUT43), .ZN(new_n683_));
  AOI22_X1  g482(.A1(new_n681_), .A2(KEYINPUT43), .B1(new_n633_), .B2(new_n683_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n569_), .A2(new_n571_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n624_), .A3(new_n619_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n678_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n681_), .A2(KEYINPUT43), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n633_), .A2(new_n683_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n625_), .A2(new_n618_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(KEYINPUT44), .A3(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n687_), .A2(new_n692_), .A3(G29gat), .A4(new_n637_), .ZN(new_n693_));
  INV_X1    g492(.A(G29gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n634_), .A2(new_n618_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n651_), .A2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n696_), .B2(new_n473_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n693_), .A2(new_n697_), .ZN(G1328gat));
  NAND3_X1  g497(.A1(new_n687_), .A2(new_n692_), .A3(new_n645_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G36gat), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n466_), .A2(G36gat), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n696_), .A2(KEYINPUT45), .A3(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT45), .B1(new_n696_), .B2(new_n701_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n700_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n700_), .A2(KEYINPUT46), .A3(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1329gat));
  NAND4_X1  g508(.A1(new_n687_), .A2(new_n692_), .A3(G43gat), .A4(new_n459_), .ZN(new_n710_));
  INV_X1    g509(.A(G43gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n711_), .B1(new_n696_), .B2(new_n458_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g513(.A1(new_n696_), .A2(G50gat), .A3(new_n435_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n687_), .A2(new_n692_), .A3(new_n436_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT115), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(new_n717_), .A3(G50gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n716_), .B2(G50gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n715_), .B1(new_n718_), .B2(new_n719_), .ZN(G1331gat));
  INV_X1    g519(.A(G57gat), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n624_), .B(new_n685_), .C1(new_n474_), .C2(new_n461_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n620_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n721_), .B1(new_n723_), .B2(new_n473_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT116), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(KEYINPUT116), .B(new_n721_), .C1(new_n723_), .C2(new_n473_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n685_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n618_), .A2(new_n251_), .A3(new_n248_), .ZN(new_n729_));
  AND4_X1   g528(.A1(new_n728_), .A2(new_n634_), .A3(new_n633_), .A4(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n473_), .A2(new_n721_), .ZN(new_n731_));
  AOI22_X1  g530(.A1(new_n726_), .A2(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1332gat));
  INV_X1    g531(.A(G64gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n730_), .B2(new_n645_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT48), .Z(new_n735_));
  INV_X1    g534(.A(new_n723_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n733_), .A3(new_n645_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1333gat));
  AOI21_X1  g537(.A(new_n438_), .B1(new_n730_), .B2(new_n459_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT49), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n736_), .A2(new_n438_), .A3(new_n459_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1334gat));
  AOI21_X1  g541(.A(new_n530_), .B1(new_n730_), .B2(new_n436_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT50), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n736_), .A2(new_n530_), .A3(new_n436_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1335gat));
  AND2_X1   g545(.A1(new_n722_), .A2(new_n695_), .ZN(new_n747_));
  INV_X1    g546(.A(G85gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n637_), .ZN(new_n749_));
  AOI211_X1 g548(.A(new_n624_), .B(new_n618_), .C1(new_n569_), .C2(new_n571_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n690_), .A2(new_n750_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(new_n637_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n749_), .B1(new_n748_), .B2(new_n752_), .ZN(G1336gat));
  INV_X1    g552(.A(G92gat), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n722_), .A2(new_n695_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(new_n466_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT117), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT117), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n758_), .B(new_n754_), .C1(new_n755_), .C2(new_n466_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n466_), .A2(new_n754_), .ZN(new_n760_));
  AOI22_X1  g559(.A1(new_n757_), .A2(new_n759_), .B1(new_n751_), .B2(new_n760_), .ZN(G1337gat));
  NAND3_X1  g560(.A1(new_n747_), .A2(new_n484_), .A3(new_n459_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n751_), .A2(new_n459_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n762_), .B(new_n763_), .C1(new_n764_), .C2(new_n452_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n484_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n755_), .A2(new_n766_), .A3(new_n458_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n452_), .B1(new_n751_), .B2(new_n459_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT51), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n765_), .A2(new_n769_), .ZN(G1338gat));
  NAND3_X1  g569(.A1(new_n690_), .A2(new_n436_), .A3(new_n750_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(KEYINPUT118), .B(KEYINPUT52), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n771_), .A2(G106gat), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n771_), .B2(G106gat), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n436_), .A2(new_n485_), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n773_), .A2(new_n774_), .B1(new_n755_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT53), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778_));
  OAI221_X1 g577(.A(new_n778_), .B1(new_n755_), .B2(new_n775_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1339gat));
  OAI21_X1  g579(.A(new_n564_), .B1(new_n250_), .B2(new_n246_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n542_), .A2(new_n476_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT12), .B1(new_n525_), .B2(new_n537_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n548_), .A2(new_n549_), .A3(new_n536_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT55), .B1(new_n785_), .B2(KEYINPUT120), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT120), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n552_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n550_), .A2(new_n551_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n477_), .B1(new_n790_), .B2(new_n544_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n786_), .A2(new_n789_), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n562_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT56), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n792_), .A2(KEYINPUT56), .A3(new_n562_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n781_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n231_), .B1(new_n235_), .B2(new_n228_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n227_), .A2(new_n229_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n798_), .B(new_n242_), .C1(new_n799_), .C2(new_n231_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n244_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT57), .B(new_n634_), .C1(new_n797_), .C2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT121), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n634_), .B1(new_n797_), .B2(new_n802_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n553_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n245_), .A2(new_n247_), .B1(new_n809_), .B2(new_n560_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n792_), .A2(KEYINPUT56), .A3(new_n562_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT56), .B1(new_n792_), .B2(new_n562_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n801_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n565_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n816_), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n634_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n801_), .B1(new_n809_), .B2(new_n560_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT58), .B(new_n818_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n603_), .A3(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n805_), .A2(new_n808_), .A3(new_n817_), .A4(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n619_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n682_), .A2(new_n729_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n567_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n826_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n570_), .A2(new_n682_), .A3(new_n729_), .A4(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n825_), .A2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n645_), .A2(new_n467_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n637_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(G113gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n624_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n835_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n473_), .B1(new_n825_), .B2(new_n832_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(KEYINPUT59), .A3(new_n834_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n253_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n838_), .B1(new_n843_), .B2(new_n837_), .ZN(G1340gat));
  XOR2_X1   g643(.A(KEYINPUT122), .B(G120gat), .Z(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n685_), .B2(KEYINPUT60), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n836_), .B(new_n846_), .C1(KEYINPUT60), .C2(new_n845_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n685_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(new_n845_), .ZN(G1341gat));
  INV_X1    g648(.A(G127gat), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n619_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n853_));
  AOI21_X1  g652(.A(G127gat), .B1(new_n836_), .B2(new_n618_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT123), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT59), .B1(new_n841_), .B2(new_n834_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n831_), .B1(new_n824_), .B2(new_n619_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n834_), .ZN(new_n858_));
  NOR4_X1   g657(.A1(new_n857_), .A2(new_n839_), .A3(new_n473_), .A4(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n851_), .B1(new_n856_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n850_), .B1(new_n835_), .B2(new_n619_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n855_), .A2(new_n863_), .ZN(G1342gat));
  INV_X1    g663(.A(G134gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n836_), .A2(new_n865_), .A3(new_n602_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n682_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n865_), .ZN(G1343gat));
  NOR4_X1   g667(.A1(new_n857_), .A2(new_n473_), .A3(new_n645_), .A4(new_n468_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n624_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n728_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT124), .B(G148gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1345gat));
  NAND2_X1  g673(.A1(new_n869_), .A2(new_n618_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1346gat));
  AOI21_X1  g676(.A(G162gat), .B1(new_n869_), .B2(new_n602_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n680_), .A2(G162gat), .A3(new_n679_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT125), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n869_), .B2(new_n880_), .ZN(G1347gat));
  NOR3_X1   g680(.A1(new_n637_), .A2(new_n466_), .A3(new_n458_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n883_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n436_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n833_), .A2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n624_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G169gat), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n888_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n892_));
  INV_X1    g691(.A(new_n318_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n891_), .B(new_n892_), .C1(new_n893_), .C2(new_n888_), .ZN(G1348gat));
  AOI21_X1  g693(.A(new_n317_), .B1(new_n887_), .B2(new_n728_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n833_), .A2(new_n886_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n896_), .A2(G176gat), .A3(new_n685_), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT127), .B1(new_n895_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(G176gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n887_), .A2(new_n899_), .A3(new_n728_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT127), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n896_), .A2(new_n685_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n900_), .B(new_n901_), .C1(new_n317_), .C2(new_n902_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n898_), .A2(new_n903_), .ZN(G1349gat));
  NOR2_X1   g703(.A1(new_n896_), .A2(new_n619_), .ZN(new_n905_));
  MUX2_X1   g704(.A(G183gat), .B(new_n342_), .S(new_n905_), .Z(G1350gat));
  NAND3_X1  g705(.A1(new_n887_), .A2(new_n602_), .A3(new_n365_), .ZN(new_n907_));
  OAI21_X1  g706(.A(G190gat), .B1(new_n896_), .B2(new_n682_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1351gat));
  NOR4_X1   g708(.A1(new_n857_), .A2(new_n637_), .A3(new_n466_), .A4(new_n468_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n624_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n728_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n618_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT63), .B(G211gat), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n915_), .B2(new_n918_), .ZN(G1354gat));
  INV_X1    g718(.A(G218gat), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n910_), .A2(new_n920_), .A3(new_n602_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n910_), .A2(new_n603_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n920_), .ZN(G1355gat));
endmodule


