//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n969_, new_n970_, new_n971_, new_n973_,
    new_n974_, new_n975_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n982_, new_n983_, new_n984_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(G50gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205_));
  NOR3_X1   g004(.A1(new_n204_), .A2(new_n205_), .A3(G43gat), .ZN(new_n206_));
  INV_X1    g005(.A(G43gat), .ZN(new_n207_));
  OR2_X1    g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G29gat), .A2(G36gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n203_), .B1(new_n206_), .B2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n212_));
  OAI21_X1  g011(.A(G43gat), .B1(new_n204_), .B2(new_n205_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(new_n213_), .A3(G50gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G99gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT10), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT10), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G99gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT64), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G92gat), .ZN(new_n227_));
  NOR3_X1   g026(.A1(new_n227_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(G92gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(G85gat), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G85gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(G92gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n227_), .A2(G85gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT9), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G99gat), .A2(G106gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT6), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n226_), .A2(new_n231_), .A3(new_n235_), .A4(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT7), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(new_n216_), .A3(new_n221_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n243_), .A2(new_n238_), .A3(new_n239_), .A4(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(G85gat), .B(G92gat), .Z(new_n246_));
  NAND2_X1  g045(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n215_), .B(new_n241_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n249_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n226_), .A2(new_n235_), .A3(new_n240_), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n251_), .A2(new_n252_), .B1(new_n253_), .B2(new_n231_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT15), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n212_), .A2(new_n213_), .A3(G50gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(G50gat), .B1(new_n212_), .B2(new_n213_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n211_), .A2(KEYINPUT15), .A3(new_n214_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n250_), .B1(new_n254_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT70), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G232gat), .A2(G233gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT34), .Z(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n261_), .A2(KEYINPUT70), .A3(new_n264_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT35), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n261_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n264_), .B1(new_n261_), .B2(KEYINPUT70), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n241_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(new_n259_), .A3(new_n258_), .ZN(new_n274_));
  AOI211_X1 g073(.A(new_n272_), .B(new_n265_), .C1(new_n274_), .C2(new_n250_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n268_), .B1(new_n271_), .B2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n270_), .A2(new_n276_), .A3(KEYINPUT36), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G190gat), .B(G218gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G134gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(G162gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n270_), .A2(new_n276_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT36), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n281_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n283_), .B1(new_n281_), .B2(new_n285_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n202_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n281_), .A2(new_n285_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n283_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n281_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(KEYINPUT37), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G57gat), .ZN(new_n294_));
  INV_X1    g093(.A(G64gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G57gat), .A2(G64gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT11), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT67), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(G71gat), .ZN(new_n301_));
  INV_X1    g100(.A(G71gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n302_), .A2(KEYINPUT67), .ZN(new_n303_));
  OAI21_X1  g102(.A(G78gat), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT11), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n296_), .A2(new_n305_), .A3(new_n297_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(KEYINPUT67), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n300_), .A2(G71gat), .ZN(new_n308_));
  INV_X1    g107(.A(G78gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n299_), .A2(new_n304_), .A3(new_n306_), .A4(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n305_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n309_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G231gat), .A2(G233gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT14), .ZN(new_n320_));
  AND2_X1   g119(.A1(KEYINPUT72), .A2(G8gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(KEYINPUT72), .A2(G8gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n320_), .B1(new_n323_), .B2(G1gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(G15gat), .B(G22gat), .Z(new_n325_));
  NOR3_X1   g124(.A1(new_n324_), .A2(KEYINPUT73), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT72), .B(G8gat), .ZN(new_n328_));
  INV_X1    g127(.A(G1gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT14), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n325_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n327_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(G1gat), .B1(new_n326_), .B2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT73), .B1(new_n324_), .B2(new_n325_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n330_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n329_), .A3(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(G8gat), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(G8gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n336_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n329_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n319_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n337_), .ZN(new_n343_));
  AOI21_X1  g142(.A(G8gat), .B1(new_n333_), .B2(new_n336_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n318_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n346_), .A2(KEYINPUT74), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT16), .B(G183gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(G211gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G127gat), .B(G155gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n349_), .B(new_n350_), .Z(new_n351_));
  INV_X1    g150(.A(KEYINPUT17), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n347_), .B(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n346_), .A2(new_n352_), .A3(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n288_), .A2(new_n293_), .A3(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT75), .ZN(new_n358_));
  INV_X1    g157(.A(new_n316_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n273_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n316_), .B(new_n241_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(KEYINPUT12), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT12), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n359_), .A2(new_n273_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G230gat), .A2(G233gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT68), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n369_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n367_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G120gat), .B(G148gat), .ZN(new_n373_));
  INV_X1    g172(.A(G204gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT5), .ZN(new_n376_));
  INV_X1    g175(.A(G176gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n372_), .A2(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n367_), .A2(new_n370_), .A3(new_n371_), .A4(new_n378_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n382_), .A2(KEYINPUT13), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(KEYINPUT13), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT69), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G113gat), .B(G141gat), .ZN(new_n388_));
  INV_X1    g187(.A(G169gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(G197gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n215_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G229gat), .A2(G233gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n341_), .A2(new_n337_), .A3(new_n260_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n341_), .A2(new_n337_), .A3(new_n215_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n395_), .B1(new_n394_), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n392_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n395_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n343_), .A2(new_n344_), .A3(new_n393_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n215_), .B1(new_n341_), .B2(new_n337_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n392_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT95), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n410_), .A2(KEYINPUT33), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT85), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT2), .ZN(new_n415_));
  OR3_X1    g214(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT2), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n413_), .A2(KEYINPUT85), .A3(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .A4(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(G155gat), .A2(G162gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT1), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(G141gat), .ZN(new_n427_));
  INV_X1    g226(.A(G148gat), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n421_), .A2(KEYINPUT1), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n413_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n430_), .ZN(new_n431_));
  OR2_X1    g230(.A1(G113gat), .A2(G120gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G113gat), .A2(G120gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT83), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(new_n436_), .A3(new_n433_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G127gat), .B(G134gat), .Z(new_n438_));
  AND3_X1   g237(.A1(new_n435_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n439_), .A2(new_n440_), .A3(KEYINPUT84), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n435_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT84), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n431_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n431_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G225gat), .A2(G233gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT94), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n435_), .A2(new_n437_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n438_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(new_n443_), .A3(new_n442_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n439_), .A2(KEYINPUT84), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n456_), .A2(new_n457_), .B1(new_n424_), .B2(new_n430_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT4), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n452_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n445_), .A2(KEYINPUT4), .A3(new_n447_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n445_), .A2(new_n447_), .A3(new_n452_), .A4(KEYINPUT4), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n451_), .B1(new_n464_), .B2(new_n450_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT0), .B(G57gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(G85gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(G1gat), .B(G29gat), .Z(new_n468_));
  XOR2_X1   g267(.A(new_n467_), .B(new_n468_), .Z(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n412_), .B1(new_n465_), .B2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n449_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n472_));
  NOR4_X1   g271(.A1(new_n472_), .A2(new_n451_), .A3(new_n469_), .A4(new_n411_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  OR2_X1    g273(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G183gat), .A2(G190gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT77), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT77), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n475_), .A2(new_n480_), .A3(new_n476_), .A4(new_n477_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n479_), .B(new_n481_), .C1(KEYINPUT23), .C2(new_n476_), .ZN(new_n482_));
  OR2_X1    g281(.A1(G183gat), .A2(G190gat), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n482_), .A2(new_n483_), .B1(G169gat), .B2(G176gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT22), .B(G169gat), .Z(new_n485_));
  OR2_X1    g284(.A1(new_n485_), .A2(G176gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT24), .B1(new_n389_), .B2(new_n377_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G169gat), .A2(G176gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT25), .B(G183gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT26), .B(G190gat), .ZN(new_n493_));
  AOI211_X1 g292(.A(new_n488_), .B(new_n491_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n475_), .A2(new_n477_), .ZN(new_n495_));
  MUX2_X1   g294(.A(new_n495_), .B(KEYINPUT23), .S(new_n476_), .Z(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n487_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G197gat), .B(G204gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT87), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT87), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(new_n391_), .A3(G204gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(KEYINPUT21), .A3(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G211gat), .B(G218gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT21), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT88), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n505_), .A2(KEYINPUT88), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n499_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT89), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n503_), .A2(new_n511_), .A3(new_n504_), .A4(new_n508_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n504_), .A2(new_n499_), .A3(new_n505_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n498_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n484_), .A2(new_n486_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n514_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT91), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n496_), .A2(new_n483_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT22), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT78), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n525_), .A2(new_n490_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT79), .B1(new_n525_), .B2(new_n389_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT79), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n377_), .B1(new_n528_), .B2(KEYINPUT22), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n526_), .A2(new_n527_), .B1(G169gat), .B2(new_n529_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n494_), .A2(new_n482_), .B1(new_n523_), .B2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n522_), .B1(new_n520_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n518_), .A2(new_n521_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G226gat), .A2(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT19), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n535_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n522_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n531_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT92), .B1(new_n516_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT92), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n520_), .A2(new_n531_), .A3(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n537_), .B(new_n538_), .C1(new_n540_), .C2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n536_), .A2(KEYINPUT93), .A3(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n540_), .A2(new_n542_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT93), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(new_n537_), .A4(new_n538_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT18), .B(G64gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(G92gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G8gat), .B(G36gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  NAND2_X1  g351(.A1(new_n548_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n552_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n544_), .A2(new_n547_), .A3(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n469_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT96), .Z(new_n557_));
  INV_X1    g356(.A(new_n464_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n557_), .B1(new_n450_), .B2(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n474_), .A2(new_n553_), .A3(new_n555_), .A4(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n552_), .A2(KEYINPUT32), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n548_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n465_), .A2(new_n470_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n469_), .B1(new_n472_), .B2(new_n451_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(KEYINPUT97), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n465_), .A2(new_n566_), .A3(new_n470_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n540_), .A2(new_n542_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n538_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n535_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n535_), .B2(new_n533_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n561_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n562_), .A2(new_n565_), .A3(new_n567_), .A4(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n560_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT82), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT31), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n441_), .A2(new_n577_), .A3(new_n444_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT31), .B1(new_n456_), .B2(new_n457_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n576_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n531_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n577_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n456_), .A2(new_n457_), .A3(KEYINPUT31), .ZN(new_n583_));
  AOI21_X1  g382(.A(KEYINPUT82), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n539_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G15gat), .B(G43gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n581_), .A2(new_n585_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n581_), .B2(new_n585_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G227gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT30), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G71gat), .B(G99gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n593_), .B(new_n594_), .Z(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n590_), .A2(new_n591_), .A3(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n580_), .A2(new_n531_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n584_), .A2(new_n539_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n588_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n581_), .A2(new_n585_), .A3(new_n589_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n595_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n597_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT29), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n446_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n520_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT86), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(G233gat), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n607_), .A2(G233gat), .ZN(new_n610_));
  OAI21_X1  g409(.A(G228gat), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n606_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n611_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n520_), .A2(new_n605_), .A3(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G22gat), .B(G50gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT28), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n446_), .A2(new_n604_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n617_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n619_), .B1(new_n431_), .B2(KEYINPUT29), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(G78gat), .B(G106gat), .Z(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(KEYINPUT90), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n618_), .A2(new_n625_), .A3(new_n620_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n615_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n624_), .B(new_n626_), .C1(new_n612_), .C2(new_n614_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n603_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n575_), .A2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n630_), .B1(new_n597_), .B2(new_n602_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n630_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n596_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n600_), .A2(new_n595_), .A3(new_n601_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  AOI22_X1  g437(.A1(new_n634_), .A2(new_n638_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n543_), .A2(KEYINPUT93), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n546_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n543_), .B2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT98), .B1(new_n642_), .B2(new_n554_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT27), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n571_), .B2(new_n554_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n548_), .A2(new_n646_), .A3(new_n552_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n643_), .A2(new_n645_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n553_), .A2(new_n555_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(new_n644_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n639_), .A2(new_n648_), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n409_), .B1(new_n633_), .B2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(KEYINPUT99), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n654_));
  AOI211_X1 g453(.A(new_n654_), .B(new_n409_), .C1(new_n633_), .C2(new_n651_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n358_), .B(new_n387_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n565_), .A2(new_n567_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n657_), .A2(new_n329_), .A3(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  OR3_X1    g461(.A1(new_n660_), .A2(KEYINPUT101), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n356_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n286_), .A2(new_n287_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n652_), .A2(new_n385_), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT102), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n652_), .A2(new_n385_), .A3(new_n666_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n658_), .B1(new_n668_), .B2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n661_), .B1(new_n672_), .B2(new_n329_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n660_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT101), .B1(new_n660_), .B2(new_n662_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n663_), .A2(new_n674_), .A3(new_n675_), .ZN(G1324gat));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT39), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n648_), .A2(new_n650_), .ZN(new_n680_));
  AOI211_X1 g479(.A(new_n338_), .B(new_n679_), .C1(new_n667_), .C2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n677_), .A2(new_n678_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n657_), .A2(new_n328_), .A3(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n682_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n683_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1325gat));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n603_), .B1(new_n668_), .B2(new_n671_), .ZN(new_n690_));
  INV_X1    g489(.A(G15gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT104), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n690_), .A2(KEYINPUT104), .A3(new_n691_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n689_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n694_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(KEYINPUT41), .A3(new_n692_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n603_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n657_), .A2(new_n691_), .A3(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n695_), .A2(new_n697_), .A3(new_n699_), .ZN(G1326gat));
  INV_X1    g499(.A(G22gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n657_), .A2(new_n701_), .A3(new_n635_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n668_), .A2(new_n671_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n635_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n703_), .B1(new_n705_), .B2(G22gat), .ZN(new_n706_));
  AOI211_X1 g505(.A(KEYINPUT42), .B(new_n701_), .C1(new_n704_), .C2(new_n635_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n702_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n702_), .B(KEYINPUT105), .C1(new_n706_), .C2(new_n707_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1327gat));
  AND2_X1   g511(.A1(new_n288_), .A2(new_n293_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n633_), .B2(new_n651_), .ZN(new_n714_));
  AND2_X1   g513(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n715_));
  NOR2_X1   g514(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n664_), .B1(new_n714_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n633_), .A2(new_n651_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n288_), .A2(new_n293_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n720_), .A2(new_n721_), .A3(new_n715_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n719_), .A2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n723_), .A2(new_n385_), .A3(new_n408_), .A4(new_n725_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n639_), .A2(new_n648_), .A3(new_n650_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n631_), .B1(new_n560_), .B2(new_n574_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n721_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n356_), .B1(new_n729_), .B2(new_n717_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n714_), .A2(new_n715_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n730_), .A2(new_n385_), .A3(new_n408_), .A4(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n724_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n726_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G29gat), .B1(new_n734_), .B2(new_n658_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n291_), .A2(new_n292_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(new_n356_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n385_), .B(new_n737_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n658_), .A2(G29gat), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT108), .Z(new_n740_));
  OAI21_X1  g539(.A(new_n735_), .B1(new_n738_), .B2(new_n740_), .ZN(G1328gat));
  NAND3_X1  g540(.A1(new_n726_), .A2(new_n733_), .A3(new_n680_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G36gat), .ZN(new_n743_));
  INV_X1    g542(.A(new_n680_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(G36gat), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT109), .B1(new_n738_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n385_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n408_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n654_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n652_), .A2(KEYINPUT99), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n748_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n737_), .A4(new_n745_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n747_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n747_), .A2(KEYINPUT45), .A3(new_n754_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n743_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n743_), .A2(new_n757_), .A3(KEYINPUT46), .A4(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1329gat));
  OAI21_X1  g562(.A(G43gat), .B1(new_n734_), .B2(new_n603_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n738_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(new_n207_), .A3(new_n698_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n764_), .A2(new_n768_), .A3(new_n766_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1330gat));
  OAI21_X1  g571(.A(G50gat), .B1(new_n734_), .B2(new_n630_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n765_), .A2(new_n203_), .A3(new_n635_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1331gat));
  AND3_X1   g574(.A1(new_n720_), .A2(new_n386_), .A3(new_n409_), .ZN(new_n776_));
  AND4_X1   g575(.A1(G57gat), .A2(new_n776_), .A3(new_n659_), .A4(new_n666_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n358_), .A2(new_n720_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n385_), .A2(new_n408_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G57gat), .B1(new_n781_), .B2(new_n659_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n782_), .A2(KEYINPUT111), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(KEYINPUT111), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n777_), .B1(new_n783_), .B2(new_n784_), .ZN(G1332gat));
  NAND3_X1  g584(.A1(new_n776_), .A2(new_n680_), .A3(new_n666_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(G64gat), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT48), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n787_), .B1(new_n786_), .B2(G64gat), .ZN(new_n791_));
  OR3_X1    g590(.A1(new_n789_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n781_), .A2(new_n295_), .A3(new_n680_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n790_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(G1333gat));
  NAND3_X1  g594(.A1(new_n776_), .A2(new_n698_), .A3(new_n666_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(G71gat), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(KEYINPUT49), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(KEYINPUT49), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n698_), .A2(new_n302_), .ZN(new_n800_));
  OAI22_X1  g599(.A1(new_n798_), .A2(new_n799_), .B1(new_n780_), .B2(new_n800_), .ZN(new_n801_));
  XOR2_X1   g600(.A(new_n801_), .B(KEYINPUT113), .Z(G1334gat));
  NAND3_X1  g601(.A1(new_n781_), .A2(new_n309_), .A3(new_n635_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n776_), .A2(new_n635_), .A3(new_n666_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(G78gat), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(KEYINPUT50), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n805_), .A2(KEYINPUT50), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1335gat));
  NAND2_X1  g609(.A1(new_n776_), .A2(new_n737_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G85gat), .B1(new_n812_), .B2(new_n659_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n730_), .A2(new_n731_), .A3(new_n779_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(new_n232_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n813_), .B1(new_n816_), .B2(new_n659_), .ZN(G1336gat));
  AOI21_X1  g616(.A(G92gat), .B1(new_n812_), .B2(new_n680_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n230_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n229_), .A2(G92gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n744_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n818_), .B1(new_n814_), .B2(new_n821_), .ZN(G1337gat));
  OAI21_X1  g621(.A(G99gat), .B1(new_n815_), .B2(new_n603_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n812_), .A2(new_n220_), .A3(new_n698_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g625(.A1(new_n812_), .A2(new_n225_), .A3(new_n635_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n814_), .A2(new_n635_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(G106gat), .ZN(new_n830_));
  AOI211_X1 g629(.A(KEYINPUT52), .B(new_n221_), .C1(new_n814_), .C2(new_n635_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n827_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT53), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n827_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1339gat));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n385_), .A2(new_n409_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n357_), .A2(KEYINPUT115), .A3(new_n837_), .A4(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT54), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n288_), .A2(new_n293_), .A3(new_n356_), .A4(new_n842_), .ZN(new_n843_));
  OAI22_X1  g642(.A1(new_n843_), .A2(new_n838_), .B1(new_n841_), .B2(KEYINPUT54), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n840_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n395_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n394_), .A2(new_n401_), .A3(new_n396_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n392_), .A3(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n407_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT55), .B1(new_n365_), .B2(new_n366_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853_));
  INV_X1    g652(.A(new_n366_), .ZN(new_n854_));
  AOI211_X1 g653(.A(new_n853_), .B(new_n854_), .C1(new_n362_), .C2(new_n364_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n362_), .A2(new_n854_), .A3(new_n364_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n852_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n851_), .B1(new_n858_), .B2(new_n378_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n367_), .A2(new_n853_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n365_), .A2(KEYINPUT55), .A3(new_n366_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n856_), .A3(new_n861_), .ZN(new_n862_));
  OR2_X1    g661(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n862_), .A2(new_n379_), .A3(new_n850_), .A4(new_n863_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n849_), .A2(new_n859_), .A3(new_n864_), .A4(new_n381_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(KEYINPUT58), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n850_), .B1(new_n862_), .B2(new_n379_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n407_), .A2(new_n848_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n867_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n871_), .A2(new_n381_), .A3(new_n872_), .A4(new_n864_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n868_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n293_), .B2(new_n288_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n862_), .A2(new_n379_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n877_), .A2(new_n879_), .B1(new_n400_), .B2(new_n407_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n381_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n852_), .A2(new_n855_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n378_), .B1(new_n882_), .B2(new_n856_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n883_), .B2(new_n878_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n880_), .A2(new_n884_), .B1(new_n382_), .B2(new_n849_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n876_), .B1(new_n885_), .B2(new_n665_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n877_), .A2(new_n879_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n862_), .A2(new_n379_), .A3(new_n878_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n887_), .A2(new_n408_), .A3(new_n888_), .A4(new_n381_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n849_), .A2(new_n382_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n736_), .A3(KEYINPUT57), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n886_), .A2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n664_), .B1(new_n875_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n845_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(KEYINPUT119), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n680_), .A2(new_n658_), .A3(new_n634_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n845_), .A2(new_n894_), .A3(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n896_), .A2(new_n897_), .A3(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G113gat), .B1(new_n901_), .B2(new_n408_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n895_), .A2(new_n903_), .A3(new_n897_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n900_), .B2(KEYINPUT59), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n905_), .A2(new_n408_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n902_), .B1(new_n906_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g706(.A(G120gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n385_), .B2(KEYINPUT60), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n901_), .B(new_n909_), .C1(KEYINPUT60), .C2(new_n908_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n905_), .A2(new_n386_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n908_), .ZN(G1341gat));
  NAND2_X1  g711(.A1(new_n356_), .A2(G127gat), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT120), .Z(new_n914_));
  NAND2_X1  g713(.A1(new_n905_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(G127gat), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n900_), .B2(new_n664_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n915_), .A2(KEYINPUT121), .A3(new_n917_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1342gat));
  AOI21_X1  g721(.A(G134gat), .B1(new_n901_), .B2(new_n665_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n905_), .A2(new_n721_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n924_), .B2(G134gat), .ZN(G1343gat));
  AND3_X1   g724(.A1(new_n845_), .A2(new_n894_), .A3(new_n898_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n898_), .B1(new_n845_), .B2(new_n894_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n926_), .A2(new_n927_), .A3(new_n638_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n680_), .A2(new_n658_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(new_n409_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(new_n427_), .ZN(G1344gat));
  NOR2_X1   g731(.A1(new_n930_), .A2(new_n387_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n428_), .ZN(G1345gat));
  INV_X1    g733(.A(new_n930_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n356_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT61), .B(G155gat), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n936_), .B(new_n937_), .ZN(G1346gat));
  AND3_X1   g737(.A1(new_n935_), .A2(G162gat), .A3(new_n721_), .ZN(new_n939_));
  AOI21_X1  g738(.A(G162gat), .B1(new_n935_), .B2(new_n665_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1347gat));
  NOR3_X1   g740(.A1(new_n744_), .A2(new_n659_), .A3(new_n634_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n895_), .A2(new_n942_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n943_), .A2(new_n409_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n389_), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n945_), .B(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n944_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n485_), .B2(new_n948_), .ZN(G1348gat));
  OAI21_X1  g748(.A(new_n377_), .B1(new_n943_), .B2(new_n385_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n926_), .A2(new_n927_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n744_), .A2(new_n659_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n951_), .A2(new_n630_), .A3(new_n952_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n386_), .A2(G176gat), .A3(new_n698_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n950_), .B1(new_n953_), .B2(new_n954_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(KEYINPUT122), .ZN(G1349gat));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n957_));
  NAND4_X1  g756(.A1(new_n951_), .A2(new_n957_), .A3(new_n356_), .A4(new_n942_), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n896_), .A2(new_n356_), .A3(new_n899_), .A4(new_n942_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(KEYINPUT123), .ZN(new_n960_));
  INV_X1    g759(.A(G183gat), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n958_), .A2(new_n960_), .A3(new_n961_), .ZN(new_n962_));
  OR3_X1    g761(.A1(new_n943_), .A2(new_n664_), .A3(new_n492_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT124), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n962_), .A2(KEYINPUT124), .A3(new_n963_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(new_n967_), .ZN(G1350gat));
  OAI21_X1  g767(.A(G190gat), .B1(new_n943_), .B2(new_n713_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n665_), .A2(new_n493_), .ZN(new_n970_));
  XOR2_X1   g769(.A(new_n970_), .B(KEYINPUT125), .Z(new_n971_));
  OAI21_X1  g770(.A(new_n969_), .B1(new_n943_), .B2(new_n971_), .ZN(G1351gat));
  INV_X1    g771(.A(new_n638_), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n951_), .A2(new_n973_), .A3(new_n952_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n974_), .A2(new_n409_), .ZN(new_n975_));
  XNOR2_X1  g774(.A(new_n975_), .B(new_n391_), .ZN(G1352gat));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977_));
  OAI22_X1  g776(.A1(new_n974_), .A2(new_n387_), .B1(new_n977_), .B2(G204gat), .ZN(new_n978_));
  OAI21_X1  g777(.A(new_n978_), .B1(KEYINPUT126), .B2(new_n374_), .ZN(new_n979_));
  OAI211_X1 g778(.A(new_n977_), .B(G204gat), .C1(new_n974_), .C2(new_n387_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n979_), .A2(new_n980_), .ZN(G1353gat));
  OR2_X1    g780(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n982_));
  XNOR2_X1  g781(.A(KEYINPUT63), .B(G211gat), .ZN(new_n983_));
  NOR2_X1   g782(.A1(new_n974_), .A2(new_n664_), .ZN(new_n984_));
  MUX2_X1   g783(.A(new_n982_), .B(new_n983_), .S(new_n984_), .Z(G1354gat));
  INV_X1    g784(.A(G218gat), .ZN(new_n986_));
  OAI21_X1  g785(.A(new_n986_), .B1(new_n974_), .B2(new_n736_), .ZN(new_n987_));
  NAND4_X1  g786(.A1(new_n928_), .A2(G218gat), .A3(new_n721_), .A4(new_n952_), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n987_), .A2(new_n988_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n989_), .A2(KEYINPUT127), .ZN(new_n990_));
  INV_X1    g789(.A(KEYINPUT127), .ZN(new_n991_));
  NAND3_X1  g790(.A1(new_n987_), .A2(new_n991_), .A3(new_n988_), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n990_), .A2(new_n992_), .ZN(G1355gat));
endmodule


