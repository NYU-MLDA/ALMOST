//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206_));
  INV_X1    g005(.A(G85gat), .ZN(new_n207_));
  INV_X1    g006(.A(G92gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n206_), .B(new_n209_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n209_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n210_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT10), .B(G99gat), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n213_), .B(new_n214_), .C1(G106gat), .C2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n218_), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(KEYINPUT6), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n217_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(KEYINPUT6), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n218_), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(KEYINPUT65), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n216_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228_));
  AND2_X1   g027(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n229_));
  NOR2_X1   g028(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n228_), .A2(new_n230_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n222_), .A2(new_n231_), .A3(new_n232_), .A4(new_n225_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT67), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n228_), .A2(new_n230_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n235_), .B1(new_n228_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(new_n225_), .A4(new_n222_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n209_), .A2(new_n210_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT68), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT8), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n209_), .A2(new_n243_), .A3(new_n210_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n241_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n234_), .A2(new_n239_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n232_), .A2(new_n231_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n223_), .A2(new_n224_), .A3(KEYINPUT69), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT69), .B1(new_n223_), .B2(new_n224_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n241_), .A2(new_n244_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT8), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n227_), .B1(new_n247_), .B2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G57gat), .B(G64gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT11), .ZN(new_n256_));
  XOR2_X1   g055(.A(G71gat), .B(G78gat), .Z(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n256_), .A2(new_n257_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n255_), .A2(KEYINPUT11), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT12), .B1(new_n254_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT12), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n245_), .B1(new_n233_), .B2(KEYINPUT67), .ZN(new_n265_));
  INV_X1    g064(.A(new_n250_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n223_), .A2(new_n224_), .A3(KEYINPUT69), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n237_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n252_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n239_), .A2(new_n265_), .B1(new_n270_), .B2(KEYINPUT8), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n264_), .B(new_n261_), .C1(new_n271_), .C2(new_n227_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G230gat), .A2(G233gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n254_), .B2(new_n262_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n263_), .A2(new_n272_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AOI211_X1 g076(.A(new_n227_), .B(new_n261_), .C1(new_n247_), .C2(new_n253_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT71), .B1(new_n278_), .B2(new_n274_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n247_), .A2(new_n253_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n227_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n262_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT70), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n281_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n261_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n254_), .A2(new_n286_), .A3(new_n262_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n283_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n277_), .A2(new_n279_), .B1(new_n288_), .B2(new_n274_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n205_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n274_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n263_), .A2(new_n272_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n282_), .A2(new_n276_), .A3(new_n273_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n279_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(KEYINPUT72), .ZN(new_n297_));
  NOR3_X1   g096(.A1(new_n291_), .A2(new_n297_), .A3(KEYINPUT73), .ZN(new_n298_));
  INV_X1    g097(.A(new_n205_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(new_n296_), .B2(KEYINPUT72), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n289_), .A2(new_n290_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n292_), .A2(new_n295_), .A3(new_n299_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n300_), .A2(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT74), .B1(new_n298_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n303_), .ZN(new_n306_));
  OAI22_X1  g105(.A1(new_n291_), .A2(new_n297_), .B1(new_n306_), .B2(KEYINPUT73), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n300_), .A2(new_n302_), .A3(new_n301_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT13), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n305_), .A2(KEYINPUT13), .A3(new_n310_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G29gat), .B(G36gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G43gat), .B(G50gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT15), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n284_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G232gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT34), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n322_), .A2(KEYINPUT35), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n254_), .A2(new_n318_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(KEYINPUT35), .A3(new_n322_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(KEYINPUT35), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n320_), .A2(new_n327_), .A3(new_n323_), .A4(new_n324_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(KEYINPUT77), .A3(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G190gat), .B(G218gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(G134gat), .B(G162gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(KEYINPUT36), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(new_n336_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n326_), .A2(KEYINPUT77), .A3(new_n328_), .A4(new_n335_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n326_), .A2(new_n328_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(KEYINPUT36), .A3(new_n334_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT37), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT37), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n339_), .A2(new_n344_), .A3(new_n341_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G1gat), .B(G8gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT78), .B(G8gat), .ZN(new_n348_));
  INV_X1    g147(.A(G1gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT14), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G15gat), .B(G22gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n347_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n353_), .A3(new_n347_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G231gat), .A2(G233gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n261_), .B(new_n358_), .Z(new_n359_));
  XNOR2_X1  g158(.A(new_n357_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT17), .ZN(new_n362_));
  XOR2_X1   g161(.A(G127gat), .B(G155gat), .Z(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G183gat), .B(G211gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  OR3_X1    g166(.A1(new_n361_), .A2(new_n362_), .A3(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(KEYINPUT17), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n361_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n315_), .A2(new_n346_), .A3(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G113gat), .B(G141gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G169gat), .B(G197gat), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n373_), .B(new_n374_), .Z(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(KEYINPUT83), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G229gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n356_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n318_), .B1(new_n379_), .B2(new_n354_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n357_), .A2(KEYINPUT81), .A3(new_n318_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n357_), .A2(new_n318_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n378_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n357_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n319_), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n378_), .B(KEYINPUT82), .Z(new_n390_));
  NAND3_X1  g189(.A1(new_n384_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n377_), .B1(new_n387_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n391_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n393_), .A2(new_n386_), .A3(new_n376_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT24), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT85), .B1(G169gat), .B2(G176gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR3_X1   g197(.A1(KEYINPUT85), .A2(G169gat), .A3(G176gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n396_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT23), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT23), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(G183gat), .A3(G190gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT86), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n409_));
  INV_X1    g208(.A(G169gat), .ZN(new_n410_));
  INV_X1    g209(.A(G176gat), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n397_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n413_), .A2(new_n396_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT86), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n416_));
  INV_X1    g215(.A(G190gat), .ZN(new_n417_));
  OR3_X1    g216(.A1(new_n416_), .A2(new_n417_), .A3(KEYINPUT26), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT25), .B(G183gat), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT26), .B1(new_n416_), .B2(new_n417_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G169gat), .A2(G176gat), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n412_), .A2(KEYINPUT24), .A3(new_n397_), .A4(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n408_), .A2(new_n415_), .A3(new_n421_), .A4(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G183gat), .A2(G190gat), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n403_), .B2(new_n401_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(new_n403_), .B2(new_n401_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n427_), .A2(new_n422_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT22), .B(G169gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT87), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n410_), .A2(KEYINPUT22), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n411_), .B1(new_n432_), .B2(KEYINPUT87), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n428_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n424_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G71gat), .B(G99gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(G43gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n435_), .B(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G127gat), .B(G134gat), .Z(new_n439_));
  XOR2_X1   g238(.A(G113gat), .B(G120gat), .Z(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n438_), .B(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G227gat), .A2(G233gat), .ZN(new_n444_));
  INV_X1    g243(.A(G15gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT30), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT31), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n443_), .B(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G155gat), .A2(G162gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT88), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT88), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(G155gat), .A3(G162gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT1), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n456_), .A2(KEYINPUT90), .ZN(new_n457_));
  NOR2_X1   g256(.A1(G155gat), .A2(G162gat), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n458_), .B1(new_n456_), .B2(KEYINPUT90), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n452_), .A2(new_n454_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n460_), .A2(KEYINPUT89), .A3(new_n455_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n452_), .A2(new_n454_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(KEYINPUT1), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n457_), .B(new_n459_), .C1(new_n461_), .C2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G141gat), .B(G148gat), .Z(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n468_), .B(KEYINPUT92), .Z(new_n469_));
  INV_X1    g268(.A(G141gat), .ZN(new_n470_));
  INV_X1    g269(.A(G148gat), .ZN(new_n471_));
  OAI22_X1  g270(.A1(new_n470_), .A2(new_n471_), .B1(KEYINPUT91), .B2(KEYINPUT2), .ZN(new_n472_));
  AND2_X1   g271(.A1(KEYINPUT91), .A2(KEYINPUT2), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT3), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n469_), .A2(new_n474_), .A3(new_n475_), .A4(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n460_), .A2(new_n458_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n467_), .A2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT99), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n481_), .A2(KEYINPUT99), .A3(new_n482_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G211gat), .B(G218gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT96), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G197gat), .ZN(new_n490_));
  INV_X1    g289(.A(G204gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT94), .B(G197gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(new_n491_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT97), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT97), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n496_), .B(new_n492_), .C1(new_n493_), .C2(new_n491_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n489_), .A2(new_n495_), .A3(KEYINPUT21), .A4(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT21), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n494_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n493_), .A2(new_n491_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT95), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n499_), .B1(G197gat), .B2(G204gat), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n502_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n488_), .B(new_n500_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n498_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G228gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT93), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n485_), .A2(new_n486_), .A3(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n481_), .A2(KEYINPUT29), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n509_), .B1(new_n512_), .B2(new_n507_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G22gat), .B(G50gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n515_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n511_), .A2(new_n513_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G78gat), .B(G106gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n481_), .A2(KEYINPUT29), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT28), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n521_), .A2(new_n522_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n520_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n525_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n520_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n523_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n519_), .A2(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n516_), .A2(new_n529_), .A3(new_n526_), .A4(new_n518_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G8gat), .B(G36gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT18), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G64gat), .B(G92gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G226gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT19), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT20), .ZN(new_n542_));
  INV_X1    g341(.A(new_n423_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT26), .B(G190gat), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT101), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n419_), .B(KEYINPUT100), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n543_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n406_), .A2(KEYINPUT102), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n406_), .A2(KEYINPUT102), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n429_), .B(KEYINPUT103), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n428_), .B1(new_n552_), .B2(G176gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n498_), .A2(new_n506_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n542_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n498_), .A2(new_n424_), .A3(new_n434_), .A4(new_n506_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n541_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n551_), .A2(new_n506_), .A3(new_n498_), .A4(new_n553_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(new_n435_), .ZN(new_n560_));
  AND4_X1   g359(.A1(KEYINPUT20), .A2(new_n559_), .A3(new_n560_), .A4(new_n541_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n538_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n406_), .B(KEYINPUT102), .ZN(new_n563_));
  INV_X1    g362(.A(new_n552_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n411_), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n563_), .A2(new_n548_), .B1(new_n565_), .B2(new_n428_), .ZN(new_n566_));
  OAI211_X1 g365(.A(KEYINPUT20), .B(new_n557_), .C1(new_n566_), .C2(new_n507_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n540_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n542_), .B1(new_n566_), .B2(new_n507_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(new_n541_), .A3(new_n560_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n570_), .A3(new_n537_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n562_), .A2(new_n571_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n465_), .A2(new_n466_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n442_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT104), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n573_), .B2(new_n442_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n481_), .A2(new_n576_), .A3(new_n441_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT4), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G225gat), .A2(G233gat), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT4), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n481_), .A2(new_n582_), .A3(new_n441_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n581_), .A3(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G1gat), .B(G29gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(new_n207_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT0), .B(G57gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n579_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n481_), .A2(new_n441_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n576_), .A3(new_n574_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n581_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n588_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n572_), .B1(new_n584_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT105), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n581_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n582_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n583_), .A2(new_n593_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n597_), .B(new_n588_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n596_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n593_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n599_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n580_), .B2(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n605_), .A2(KEYINPUT105), .A3(KEYINPUT33), .A4(new_n588_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n600_), .A2(new_n601_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n595_), .A2(new_n602_), .A3(new_n606_), .A4(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n537_), .A2(KEYINPUT32), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n568_), .A2(new_n570_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n609_), .B1(new_n610_), .B2(KEYINPUT106), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n568_), .A2(new_n570_), .A3(KEYINPUT106), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n569_), .A2(new_n560_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n540_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n556_), .A2(new_n541_), .A3(new_n557_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n614_), .A2(KEYINPUT32), .A3(new_n537_), .A4(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n611_), .B1(new_n612_), .B2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n605_), .A2(new_n588_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n600_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n617_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n533_), .B1(new_n608_), .B2(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n605_), .A2(new_n588_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT27), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n572_), .A2(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n614_), .A2(new_n615_), .ZN(new_n625_));
  OAI211_X1 g424(.A(KEYINPUT27), .B(new_n571_), .C1(new_n625_), .C2(new_n537_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n622_), .A2(new_n600_), .A3(new_n624_), .A4(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n531_), .A2(new_n532_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n450_), .B1(new_n621_), .B2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n618_), .A2(new_n619_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n449_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n626_), .A2(new_n624_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n633_), .A2(new_n628_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n395_), .B1(new_n630_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n372_), .A2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(G1gat), .A3(new_n631_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(KEYINPUT38), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT107), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(KEYINPUT38), .ZN(new_n642_));
  AOI211_X1 g441(.A(new_n342_), .B(new_n371_), .C1(new_n630_), .C2(new_n636_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n315_), .A2(new_n395_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G1gat), .B1(new_n645_), .B2(new_n631_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n641_), .A2(new_n642_), .A3(new_n646_), .ZN(G1324gat));
  INV_X1    g446(.A(KEYINPUT108), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n643_), .A2(new_n644_), .A3(new_n634_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n649_), .B2(G8gat), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n649_), .A2(new_n648_), .A3(G8gat), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n348_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n638_), .A2(new_n655_), .A3(new_n635_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(G1325gat));
  OAI21_X1  g459(.A(G15gat), .B1(new_n645_), .B2(new_n450_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT41), .Z(new_n662_));
  NAND2_X1  g461(.A1(new_n449_), .A2(new_n445_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n662_), .B1(new_n638_), .B2(new_n663_), .ZN(G1326gat));
  OAI21_X1  g463(.A(G22gat), .B1(new_n645_), .B2(new_n628_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT42), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n628_), .A2(G22gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n638_), .B2(new_n667_), .ZN(G1327gat));
  INV_X1    g467(.A(new_n346_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n630_), .B2(new_n636_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n672_), .A2(KEYINPUT44), .A3(new_n371_), .A4(new_n644_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n630_), .A2(new_n636_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n671_), .B1(new_n674_), .B2(new_n346_), .ZN(new_n675_));
  AOI211_X1 g474(.A(KEYINPUT43), .B(new_n669_), .C1(new_n630_), .C2(new_n636_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n371_), .B(new_n644_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n673_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(G29gat), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n680_), .A2(new_n681_), .A3(new_n631_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n308_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n683_), .A2(new_n684_), .A3(new_n312_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT13), .B1(new_n305_), .B2(new_n310_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n342_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n371_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n637_), .A2(new_n687_), .A3(new_n690_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n691_), .A2(new_n631_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n682_), .B1(new_n681_), .B2(new_n692_), .ZN(G1328gat));
  OAI21_X1  g492(.A(G36gat), .B1(new_n680_), .B2(new_n635_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n635_), .A2(KEYINPUT110), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n635_), .A2(KEYINPUT110), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n691_), .A2(G36gat), .A3(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT45), .Z(new_n700_));
  NAND2_X1  g499(.A1(new_n694_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n694_), .A2(KEYINPUT46), .A3(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1329gat));
  INV_X1    g504(.A(G43gat), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n450_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n673_), .A2(new_n679_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT111), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n673_), .A2(new_n679_), .A3(new_n710_), .A4(new_n707_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n706_), .B1(new_n691_), .B2(new_n450_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n709_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT47), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n709_), .A2(new_n715_), .A3(new_n711_), .A4(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1330gat));
  INV_X1    g516(.A(G50gat), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n680_), .A2(new_n718_), .A3(new_n628_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n691_), .A2(new_n628_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(new_n720_), .ZN(G1331gat));
  INV_X1    g520(.A(new_n395_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n630_), .B2(new_n636_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n346_), .A2(new_n371_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(new_n315_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n631_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G57gat), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT112), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n687_), .A2(new_n722_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(new_n643_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(G57gat), .A3(new_n726_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n728_), .A2(new_n731_), .ZN(G1332gat));
  INV_X1    g531(.A(G64gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n730_), .B2(new_n697_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT48), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n725_), .A2(new_n733_), .A3(new_n697_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1333gat));
  INV_X1    g536(.A(G71gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n730_), .B2(new_n449_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n725_), .A2(new_n738_), .A3(new_n449_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1334gat));
  INV_X1    g542(.A(G78gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n730_), .B2(new_n533_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT50), .Z(new_n746_));
  NAND3_X1  g545(.A1(new_n725_), .A2(new_n744_), .A3(new_n533_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1335gat));
  OAI211_X1 g547(.A(new_n371_), .B(new_n729_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G85gat), .B1(new_n749_), .B2(new_n631_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n723_), .A2(new_n315_), .A3(new_n690_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n751_), .A2(KEYINPUT114), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(KEYINPUT114), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n726_), .A2(new_n207_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n750_), .B1(new_n755_), .B2(new_n756_), .ZN(G1336gat));
  OAI21_X1  g556(.A(G92gat), .B1(new_n749_), .B2(new_n698_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n634_), .A2(new_n208_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n755_), .B2(new_n759_), .ZN(G1337gat));
  OAI21_X1  g559(.A(G99gat), .B1(new_n749_), .B2(new_n450_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n450_), .A2(new_n215_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n754_), .A2(KEYINPUT115), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT115), .B1(new_n754_), .B2(new_n762_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT51), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n761_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1338gat));
  INV_X1    g568(.A(G106gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n754_), .A2(new_n770_), .A3(new_n533_), .ZN(new_n771_));
  OAI21_X1  g570(.A(G106gat), .B1(new_n749_), .B2(new_n628_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(KEYINPUT52), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(G106gat), .C1(new_n749_), .C2(new_n628_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n771_), .B1(new_n773_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT53), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n771_), .C1(new_n773_), .C2(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1339gat));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n687_), .A2(new_n782_), .A3(new_n395_), .A4(new_n724_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n313_), .A2(new_n395_), .A3(new_n724_), .A4(new_n314_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT54), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n375_), .B1(new_n393_), .B2(new_n386_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n375_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n390_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n384_), .A2(new_n389_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n789_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n788_), .A2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n303_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n277_), .A2(KEYINPUT55), .A3(new_n279_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n295_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n293_), .A2(new_n283_), .A3(new_n287_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n274_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n797_), .A2(new_n799_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n205_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n205_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n796_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n795_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n342_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n306_), .B1(new_n788_), .B2(new_n793_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n806_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n205_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT58), .B(new_n812_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n346_), .A2(new_n818_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n809_), .A2(new_n811_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n807_), .B1(new_n311_), .B2(new_n794_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n810_), .B1(new_n821_), .B2(new_n342_), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n787_), .B(new_n689_), .C1(new_n820_), .C2(new_n822_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n305_), .A2(new_n310_), .B1(new_n793_), .B2(new_n788_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n811_), .B1(new_n824_), .B2(new_n807_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n817_), .A2(new_n346_), .A3(new_n818_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n342_), .B1(new_n795_), .B2(new_n808_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n825_), .B(new_n826_), .C1(new_n827_), .C2(KEYINPUT57), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT117), .B1(new_n828_), .B2(new_n371_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n786_), .B1(new_n823_), .B2(new_n829_), .ZN(new_n830_));
  NOR4_X1   g629(.A1(new_n631_), .A2(new_n533_), .A3(new_n634_), .A4(new_n450_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(KEYINPUT59), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n784_), .B(new_n782_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n689_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n831_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT59), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n834_), .A2(G113gat), .A3(new_n722_), .A4(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT57), .B1(new_n809_), .B2(new_n688_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n811_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n826_), .B1(new_n821_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n371_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n832_), .B1(new_n844_), .B2(new_n786_), .ZN(new_n845_));
  AOI21_X1  g644(.A(G113gat), .B1(new_n845_), .B2(new_n722_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT116), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n840_), .A2(new_n847_), .ZN(G1340gat));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849_));
  INV_X1    g648(.A(new_n833_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n844_), .A2(new_n787_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n828_), .A2(KEYINPUT117), .A3(new_n371_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n850_), .B1(new_n853_), .B2(new_n786_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n315_), .B1(new_n845_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n849_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n687_), .B1(new_n837_), .B2(KEYINPUT59), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n834_), .A2(new_n858_), .A3(KEYINPUT118), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n857_), .A2(G120gat), .A3(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n687_), .A2(KEYINPUT60), .ZN(new_n861_));
  MUX2_X1   g660(.A(new_n861_), .B(KEYINPUT60), .S(G120gat), .Z(new_n862_));
  NAND2_X1  g661(.A1(new_n845_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n863_), .ZN(G1341gat));
  AND2_X1   g663(.A1(new_n834_), .A2(new_n838_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n689_), .A2(G127gat), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(KEYINPUT120), .Z(new_n867_));
  AOI21_X1  g666(.A(G127gat), .B1(new_n845_), .B2(new_n689_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n868_), .A2(KEYINPUT119), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(KEYINPUT119), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n865_), .A2(new_n867_), .B1(new_n869_), .B2(new_n870_), .ZN(G1342gat));
  AOI21_X1  g670(.A(G134gat), .B1(new_n845_), .B2(new_n342_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT121), .B(G134gat), .Z(new_n873_));
  NOR2_X1   g672(.A1(new_n669_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n865_), .B2(new_n874_), .ZN(G1343gat));
  NAND2_X1  g674(.A1(new_n844_), .A2(new_n786_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n628_), .A2(new_n449_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n697_), .A2(new_n631_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n877_), .A3(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n395_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(new_n470_), .ZN(G1344gat));
  NOR2_X1   g680(.A1(new_n879_), .A2(new_n687_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(new_n471_), .ZN(G1345gat));
  AND2_X1   g682(.A1(new_n876_), .A2(new_n877_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n884_), .A2(KEYINPUT122), .A3(new_n689_), .A4(new_n878_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n879_), .B2(new_n371_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G155gat), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n885_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1346gat));
  INV_X1    g690(.A(new_n879_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G162gat), .B1(new_n892_), .B2(new_n342_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n346_), .A2(G162gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT123), .Z(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n892_), .B2(new_n895_), .ZN(G1347gat));
  NAND2_X1  g695(.A1(new_n697_), .A2(new_n633_), .ZN(new_n897_));
  XOR2_X1   g696(.A(new_n897_), .B(KEYINPUT124), .Z(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n533_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n830_), .A2(new_n722_), .A3(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n410_), .B1(new_n901_), .B2(KEYINPUT62), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(KEYINPUT125), .A3(new_n904_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n900_), .B(new_n902_), .C1(new_n901_), .C2(KEYINPUT62), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n900_), .A2(new_n552_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(G1348gat));
  NOR3_X1   g707(.A1(new_n898_), .A2(new_n411_), .A3(new_n687_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n533_), .B1(new_n844_), .B2(new_n786_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n830_), .A2(new_n315_), .A3(new_n899_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n411_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n912_), .A2(KEYINPUT126), .A3(new_n411_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n911_), .B1(new_n915_), .B2(new_n916_), .ZN(G1349gat));
  NAND2_X1  g716(.A1(new_n830_), .A2(new_n899_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n918_), .A2(new_n547_), .A3(new_n371_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n898_), .A2(new_n371_), .ZN(new_n920_));
  AOI21_X1  g719(.A(G183gat), .B1(new_n910_), .B2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n919_), .A2(new_n921_), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n918_), .B2(new_n669_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n342_), .A2(new_n546_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n918_), .B2(new_n924_), .ZN(G1351gat));
  NOR2_X1   g724(.A1(new_n698_), .A2(new_n726_), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n884_), .A2(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927_), .B2(new_n722_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n884_), .A2(new_n926_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n929_), .A2(new_n490_), .A3(new_n395_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1352gat));
  NAND3_X1  g730(.A1(new_n927_), .A2(new_n491_), .A3(new_n315_), .ZN(new_n932_));
  OAI21_X1  g731(.A(G204gat), .B1(new_n929_), .B2(new_n687_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1353gat));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n935_));
  INV_X1    g734(.A(G211gat), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n689_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(KEYINPUT127), .ZN(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(new_n940_));
  AND3_X1   g739(.A1(new_n927_), .A2(new_n937_), .A3(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n937_), .B1(new_n927_), .B2(new_n940_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1354gat));
  OAI21_X1  g742(.A(G218gat), .B1(new_n929_), .B2(new_n669_), .ZN(new_n944_));
  OR2_X1    g743(.A1(new_n688_), .A2(G218gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n929_), .B2(new_n945_), .ZN(G1355gat));
endmodule


