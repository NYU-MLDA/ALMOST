//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n909_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT81), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT83), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT2), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT84), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT84), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n207_), .A2(new_n215_), .A3(new_n210_), .A4(new_n212_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n205_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(new_n204_), .B(KEYINPUT1), .Z(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n203_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n209_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(new_n211_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n217_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G127gat), .B(G134gat), .Z(new_n224_));
  XOR2_X1   g023(.A(G113gat), .B(G120gat), .Z(new_n225_));
  XOR2_X1   g024(.A(new_n224_), .B(new_n225_), .Z(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n226_), .B1(new_n217_), .B2(new_n222_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT91), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(KEYINPUT91), .B(new_n226_), .C1(new_n217_), .C2(new_n222_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G225gat), .A2(G233gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT93), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT93), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n233_), .A2(new_n237_), .A3(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G1gat), .B(G29gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G85gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G57gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  NAND2_X1  g042(.A1(new_n233_), .A2(KEYINPUT4), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT92), .ZN(new_n245_));
  INV_X1    g044(.A(new_n229_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n234_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n244_), .A2(new_n245_), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n247_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT92), .B1(new_n253_), .B2(new_n250_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n239_), .A2(new_n243_), .A3(new_n252_), .A4(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT33), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT23), .ZN(new_n259_));
  OR2_X1    g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT22), .B(G169gat), .ZN(new_n263_));
  INV_X1    g062(.A(G176gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n261_), .A2(new_n262_), .A3(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT26), .B(G190gat), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT25), .B(G183gat), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n271_), .A2(KEYINPUT24), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT24), .A3(new_n262_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n259_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n266_), .B1(new_n270_), .B2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G211gat), .B(G218gat), .Z(new_n276_));
  INV_X1    g075(.A(KEYINPUT21), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G197gat), .B(G204gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT21), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n276_), .A3(KEYINPUT21), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n275_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT90), .ZN(new_n286_));
  OR3_X1    g085(.A1(new_n275_), .A2(new_n284_), .A3(KEYINPUT90), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT20), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G226gat), .A2(G233gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT19), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT22), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT78), .B1(new_n291_), .B2(G169gat), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n264_), .B(new_n292_), .C1(new_n263_), .C2(KEYINPUT78), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n261_), .A2(new_n293_), .A3(new_n262_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT77), .ZN(new_n295_));
  INV_X1    g094(.A(G190gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT26), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n296_), .A2(KEYINPUT26), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n269_), .B(new_n297_), .C1(new_n298_), .C2(new_n295_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n299_), .A2(new_n259_), .A3(new_n273_), .A4(new_n272_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n294_), .A2(new_n300_), .ZN(new_n301_));
  AOI211_X1 g100(.A(new_n288_), .B(new_n290_), .C1(new_n301_), .C2(new_n284_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n286_), .A2(new_n287_), .A3(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT20), .B1(new_n301_), .B2(new_n284_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n275_), .A2(new_n284_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT88), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT88), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n275_), .A2(new_n307_), .A3(new_n284_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n304_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT89), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n290_), .B(KEYINPUT87), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NOR3_X1   g111(.A1(new_n309_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n301_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n284_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n288_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n275_), .A2(new_n307_), .A3(new_n284_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n307_), .B1(new_n275_), .B2(new_n284_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT89), .B1(new_n319_), .B2(new_n311_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n303_), .B1(new_n313_), .B2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G8gat), .B(G36gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT18), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G64gat), .B(G92gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n321_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n303_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n310_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n319_), .A2(KEYINPUT89), .A3(new_n311_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n325_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n243_), .B1(new_n233_), .B2(new_n249_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n248_), .A2(new_n234_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n334_), .B1(new_n253_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT94), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n334_), .B(KEYINPUT94), .C1(new_n253_), .C2(new_n335_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n333_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n252_), .A2(new_n254_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n341_), .A2(KEYINPUT33), .A3(new_n243_), .A4(new_n239_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n257_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n238_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n237_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n252_), .B(new_n254_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n243_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n255_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n285_), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(new_n315_), .B2(new_n314_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT96), .B1(new_n285_), .B2(KEYINPUT20), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n290_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(new_n311_), .B2(new_n319_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n325_), .A2(KEYINPUT32), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT95), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n321_), .A2(new_n359_), .A3(new_n357_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT95), .B1(new_n331_), .B2(new_n356_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n358_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n343_), .B1(new_n350_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n217_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n365_), .A3(new_n221_), .ZN(new_n366_));
  XOR2_X1   g165(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n223_), .A2(new_n365_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT29), .B1(new_n217_), .B2(new_n222_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G22gat), .B(G50gat), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n284_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n374_), .B1(new_n372_), .B2(new_n284_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n371_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n379_), .A2(new_n375_), .A3(new_n370_), .A4(new_n368_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381_));
  INV_X1    g180(.A(G78gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n378_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n384_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT86), .B(G106gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n386_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n378_), .A2(new_n380_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n383_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n388_), .B1(new_n392_), .B2(new_n385_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G71gat), .B(G99gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(G43gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT30), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(new_n301_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(G15gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n397_), .A2(new_n301_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n397_), .A2(new_n301_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n401_), .A3(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n403_), .A2(KEYINPUT80), .A3(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n408_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n403_), .A2(KEYINPUT80), .A3(new_n410_), .A4(new_n406_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n409_), .A2(new_n226_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n226_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n394_), .A2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n414_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n389_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n412_), .A2(new_n413_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n392_), .A2(new_n388_), .A3(new_n385_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n349_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(new_n355_), .B2(new_n326_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n423_), .A2(new_n332_), .ZN(new_n424_));
  AOI21_X1  g223(.A(KEYINPUT27), .B1(new_n327_), .B2(new_n332_), .ZN(new_n425_));
  OR2_X1    g224(.A1(new_n425_), .A2(KEYINPUT97), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(KEYINPUT97), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n424_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n363_), .A2(new_n415_), .B1(new_n421_), .B2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G113gat), .B(G141gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G169gat), .B(G197gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n430_), .B(new_n431_), .Z(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G229gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT75), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT73), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT14), .ZN(new_n437_));
  INV_X1    g236(.A(G1gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT72), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT72), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(G1gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n437_), .B1(new_n442_), .B2(G8gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G15gat), .B(G22gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n436_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(G8gat), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n448_));
  OAI211_X1 g247(.A(KEYINPUT73), .B(new_n444_), .C1(new_n448_), .C2(new_n437_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G1gat), .B(G8gat), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n446_), .B2(new_n449_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G29gat), .B(G36gat), .Z(new_n453_));
  XOR2_X1   g252(.A(G43gat), .B(G50gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n451_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n455_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n450_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n449_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT72), .B(G1gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT14), .B1(new_n460_), .B2(new_n447_), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT73), .B1(new_n461_), .B2(new_n444_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n458_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n457_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n435_), .B1(new_n456_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n455_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n457_), .A3(new_n464_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(KEYINPUT75), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n434_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n451_), .A2(new_n452_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n455_), .B(KEYINPUT15), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n467_), .A3(new_n434_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n433_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n434_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n456_), .A2(new_n465_), .A3(new_n435_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT75), .B1(new_n467_), .B2(new_n468_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(new_n474_), .A3(new_n432_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT76), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n429_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT10), .B(G99gat), .Z(new_n485_));
  INV_X1    g284(.A(G106gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G85gat), .B(G92gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT9), .ZN(new_n489_));
  INV_X1    g288(.A(G99gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT6), .B1(new_n490_), .B2(new_n486_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(G99gat), .A3(G106gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G85gat), .ZN(new_n495_));
  INV_X1    g294(.A(G92gat), .ZN(new_n496_));
  OR3_X1    g295(.A1(new_n495_), .A2(new_n496_), .A3(KEYINPUT9), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n487_), .A2(new_n489_), .A3(new_n494_), .A4(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT7), .ZN(new_n499_));
  NOR2_X1   g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n499_), .B1(new_n500_), .B2(KEYINPUT64), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT64), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n502_), .A2(G99gat), .A3(G106gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT65), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n500_), .A2(KEYINPUT64), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n502_), .B1(G99gat), .B2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT65), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .A4(new_n499_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n490_), .A2(new_n486_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n491_), .A2(new_n493_), .B1(new_n509_), .B2(KEYINPUT7), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n504_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT8), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT66), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n488_), .A2(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n511_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n512_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n498_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT67), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT67), .B(new_n498_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G57gat), .B(G64gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(KEYINPUT11), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(KEYINPUT11), .ZN(new_n524_));
  XOR2_X1   g323(.A(G71gat), .B(G78gat), .Z(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n524_), .A2(new_n525_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT12), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n519_), .A2(new_n520_), .A3(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n498_), .B(new_n528_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT12), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n517_), .A2(new_n529_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G230gat), .A2(G233gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n532_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n533_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G120gat), .B(G148gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT5), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G176gat), .B(G204gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n544_), .B(new_n545_), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n542_), .B(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n548_), .A2(KEYINPUT13), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(KEYINPUT13), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n517_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT35), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT34), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n553_), .A2(new_n455_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n519_), .A2(new_n472_), .A3(new_n520_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT68), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n554_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n561_), .B(new_n562_), .C1(new_n517_), .C2(new_n457_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n557_), .A2(new_n554_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n560_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n564_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n566_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G134gat), .B(G162gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT69), .B(KEYINPUT36), .Z(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n565_), .A2(new_n567_), .A3(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n570_), .B(KEYINPUT36), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT37), .B1(new_n573_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT70), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n567_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n566_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT71), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT71), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n565_), .A2(new_n583_), .A3(new_n567_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n584_), .A3(new_n574_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n565_), .A2(new_n567_), .A3(new_n572_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT70), .B(KEYINPUT37), .C1(new_n573_), .C2(new_n576_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n579_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G127gat), .B(G155gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT16), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G183gat), .B(G211gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT17), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT74), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(new_n529_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n471_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n596_), .A2(new_n597_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n602_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n552_), .A2(new_n591_), .A3(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n484_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n484_), .A2(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT98), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n349_), .B(KEYINPUT99), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n611_), .A2(new_n460_), .A3(new_n613_), .A4(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT38), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n617_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n551_), .A2(new_n482_), .A3(new_n606_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT100), .Z(new_n621_));
  NAND3_X1  g420(.A1(new_n585_), .A2(KEYINPUT101), .A3(new_n587_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT101), .B1(new_n585_), .B2(new_n587_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n429_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n621_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G1gat), .B1(new_n628_), .B2(new_n350_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n618_), .A2(new_n619_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n618_), .A2(new_n619_), .A3(KEYINPUT102), .A4(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1324gat));
  XNOR2_X1  g433(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT103), .B1(new_n628_), .B2(new_n428_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n637_));
  INV_X1    g436(.A(new_n428_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n621_), .A2(new_n637_), .A3(new_n638_), .A4(new_n627_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n636_), .A2(G8gat), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n641_), .A2(KEYINPUT39), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n611_), .A2(new_n613_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n428_), .A2(G8gat), .ZN(new_n644_));
  AOI22_X1  g443(.A1(new_n640_), .A2(new_n642_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n636_), .A2(G8gat), .A3(new_n639_), .A4(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n635_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n640_), .A2(new_n642_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n643_), .A2(new_n644_), .ZN(new_n650_));
  AND4_X1   g449(.A1(new_n647_), .A2(new_n649_), .A3(new_n650_), .A4(new_n635_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n648_), .A2(new_n651_), .ZN(G1325gat));
  OAI21_X1  g451(.A(G15gat), .B1(new_n628_), .B2(new_n418_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT41), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n609_), .A2(new_n400_), .A3(new_n414_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1326gat));
  INV_X1    g455(.A(new_n394_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G22gat), .B1(new_n628_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT42), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n657_), .A2(G22gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n659_), .B1(new_n612_), .B2(new_n660_), .ZN(G1327gat));
  NAND2_X1  g460(.A1(new_n626_), .A2(new_n607_), .ZN(new_n662_));
  NOR4_X1   g461(.A1(new_n429_), .A2(new_n662_), .A3(new_n483_), .A4(new_n552_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G29gat), .B1(new_n663_), .B2(new_n349_), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT43), .B1(new_n429_), .B2(new_n590_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n257_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n362_), .B1(new_n348_), .B2(new_n255_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n415_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n416_), .A2(new_n420_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n428_), .A2(new_n669_), .A3(new_n350_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n591_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n665_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n482_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n552_), .A2(new_n675_), .A3(new_n606_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT44), .B1(new_n674_), .B2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n674_), .A2(KEYINPUT44), .A3(new_n676_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n674_), .A2(KEYINPUT106), .A3(KEYINPUT44), .A4(new_n676_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n677_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n615_), .A2(G29gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n664_), .B1(new_n682_), .B2(new_n683_), .ZN(G1328gat));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685_));
  INV_X1    g484(.A(G36gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n682_), .B2(new_n638_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n663_), .A2(new_n686_), .A3(new_n638_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT45), .Z(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n689_), .ZN(new_n691_));
  AOI211_X1 g490(.A(new_n428_), .B(new_n677_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n691_), .B(KEYINPUT46), .C1(new_n692_), .C2(new_n686_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(G1329gat));
  AOI21_X1  g493(.A(G43gat), .B1(new_n663_), .B2(new_n414_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n414_), .A2(G43gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n682_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1330gat));
  INV_X1    g498(.A(G50gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n663_), .A2(new_n700_), .A3(new_n394_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n682_), .A2(new_n702_), .A3(new_n394_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G50gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n702_), .B1(new_n682_), .B2(new_n394_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(G1331gat));
  NAND4_X1  g505(.A1(new_n627_), .A2(new_n483_), .A3(new_n552_), .A4(new_n606_), .ZN(new_n707_));
  INV_X1    g506(.A(G57gat), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n350_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT110), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n552_), .A2(new_n606_), .A3(new_n590_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n429_), .A2(new_n482_), .A3(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT108), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n713_), .A2(KEYINPUT109), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(KEYINPUT109), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n615_), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n710_), .B1(new_n716_), .B2(new_n708_), .ZN(G1332gat));
  OAI21_X1  g516(.A(G64gat), .B1(new_n707_), .B2(new_n428_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT48), .ZN(new_n719_));
  INV_X1    g518(.A(new_n713_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n428_), .A2(G64gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n720_), .B2(new_n721_), .ZN(G1333gat));
  OAI21_X1  g521(.A(G71gat), .B1(new_n707_), .B2(new_n418_), .ZN(new_n723_));
  XOR2_X1   g522(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n418_), .A2(G71gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n720_), .B2(new_n726_), .ZN(G1334gat));
  OAI21_X1  g526(.A(G78gat), .B1(new_n707_), .B2(new_n657_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT50), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n713_), .A2(new_n382_), .A3(new_n394_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1335gat));
  NAND3_X1  g530(.A1(new_n552_), .A2(new_n675_), .A3(new_n607_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n665_), .B2(new_n673_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G85gat), .B1(new_n734_), .B2(new_n350_), .ZN(new_n735_));
  NOR4_X1   g534(.A1(new_n429_), .A2(new_n662_), .A3(new_n482_), .A4(new_n551_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n495_), .A3(new_n615_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1336gat));
  OAI21_X1  g537(.A(G92gat), .B1(new_n734_), .B2(new_n428_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(new_n496_), .A3(new_n638_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1337gat));
  OAI21_X1  g540(.A(G99gat), .B1(new_n734_), .B2(new_n418_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n736_), .A2(new_n414_), .A3(new_n485_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n745_), .A2(KEYINPUT112), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n744_), .B(new_n746_), .ZN(G1338gat));
  NAND3_X1  g546(.A1(new_n736_), .A2(new_n486_), .A3(new_n394_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749_));
  AOI211_X1 g548(.A(new_n657_), .B(new_n732_), .C1(new_n665_), .C2(new_n673_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n486_), .B1(new_n750_), .B2(KEYINPUT113), .ZN(new_n751_));
  INV_X1    g550(.A(new_n732_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n672_), .B1(new_n671_), .B2(new_n591_), .ZN(new_n753_));
  AOI211_X1 g552(.A(KEYINPUT43), .B(new_n590_), .C1(new_n668_), .C2(new_n670_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n394_), .B(new_n752_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n749_), .B1(new_n751_), .B2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G106gat), .B1(new_n755_), .B2(new_n756_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT113), .B1(new_n733_), .B2(new_n394_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n759_), .A2(new_n760_), .A3(KEYINPUT52), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n748_), .B1(new_n758_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT53), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n764_), .B(new_n748_), .C1(new_n758_), .C2(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1339gat));
  NOR3_X1   g565(.A1(new_n614_), .A2(new_n638_), .A3(new_n416_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n434_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n473_), .A2(new_n467_), .A3(new_n477_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n433_), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n481_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n548_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n538_), .A2(KEYINPUT115), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n532_), .A2(new_n536_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n540_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n532_), .A2(new_n536_), .A3(KEYINPUT55), .A4(new_n537_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT115), .B1(new_n538_), .B2(new_n774_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n776_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n773_), .B1(new_n782_), .B2(new_n547_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n537_), .B1(new_n532_), .B2(new_n536_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n532_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(KEYINPUT55), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n538_), .A2(new_n774_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n789_), .A3(new_n775_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n546_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n783_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n538_), .A2(new_n541_), .A3(new_n547_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n482_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n482_), .B2(new_n794_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n772_), .B1(new_n792_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n585_), .A2(new_n587_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT101), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(KEYINPUT57), .A3(new_n622_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n798_), .A2(KEYINPUT116), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n546_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n546_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n797_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n772_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n623_), .A2(new_n624_), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n804_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n803_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n809_), .A2(new_n625_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n794_), .A2(new_n481_), .A3(new_n770_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n590_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n792_), .A2(KEYINPUT58), .A3(new_n815_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n814_), .A2(new_n810_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n606_), .B1(new_n813_), .B2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n551_), .A2(new_n590_), .A3(new_n483_), .A4(new_n606_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n767_), .B1(new_n821_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(G113gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n482_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n821_), .B2(new_n824_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n825_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  OAI221_X1 g631(.A(new_n767_), .B1(new_n829_), .B2(KEYINPUT59), .C1(new_n821_), .C2(new_n824_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n483_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n828_), .B1(new_n834_), .B2(new_n827_), .ZN(G1340gat));
  INV_X1    g634(.A(KEYINPUT60), .ZN(new_n836_));
  AOI21_X1  g635(.A(G120gat), .B1(new_n552_), .B2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n836_), .B2(G120gat), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n826_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n551_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n840_));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT118), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n844_), .B(new_n839_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1341gat));
  INV_X1    g645(.A(G127gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n826_), .A2(new_n847_), .A3(new_n606_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n607_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(G1342gat));
  XOR2_X1   g649(.A(KEYINPUT119), .B(G134gat), .Z(new_n851_));
  NAND2_X1  g650(.A1(new_n591_), .A2(new_n851_), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(KEYINPUT120), .Z(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856_));
  AOI21_X1  g655(.A(G134gat), .B1(new_n826_), .B2(new_n626_), .ZN(new_n857_));
  OR3_X1    g656(.A1(new_n855_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1343gat));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n814_), .A2(new_n810_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n818_), .A2(new_n819_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT116), .B1(new_n798_), .B2(new_n802_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n809_), .A2(new_n811_), .A3(new_n804_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .A4(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n824_), .B1(new_n866_), .B2(new_n607_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n420_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n614_), .A2(new_n638_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n861_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n420_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n871_), .B(new_n869_), .C1(new_n821_), .C2(new_n824_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(KEYINPUT122), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n482_), .B1(new_n870_), .B2(new_n873_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g674(.A1(new_n868_), .A2(new_n861_), .A3(new_n869_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n872_), .A2(KEYINPUT122), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n551_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT123), .B(G148gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1345gat));
  AOI21_X1  g679(.A(new_n607_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n881_));
  XOR2_X1   g680(.A(KEYINPUT61), .B(G155gat), .Z(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1346gat));
  INV_X1    g682(.A(G162gat), .ZN(new_n884_));
  AOI211_X1 g683(.A(new_n884_), .B(new_n590_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n625_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(G162gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n626_), .B1(new_n870_), .B2(new_n873_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n889_), .A2(KEYINPUT124), .A3(new_n884_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n885_), .B1(new_n888_), .B2(new_n890_), .ZN(G1347gat));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n892_));
  INV_X1    g691(.A(new_n867_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n614_), .A2(new_n638_), .A3(new_n414_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n894_), .A2(KEYINPUT125), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(KEYINPUT125), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n895_), .A2(new_n896_), .A3(new_n394_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n893_), .A2(new_n482_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n892_), .B1(new_n898_), .B2(G169gat), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900_));
  INV_X1    g699(.A(new_n898_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n899_), .A2(new_n900_), .B1(new_n901_), .B2(new_n263_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n899_), .A2(new_n900_), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n898_), .A2(new_n892_), .A3(G169gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(G1348gat));
  NAND2_X1  g704(.A1(new_n893_), .A2(new_n897_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n551_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n264_), .ZN(G1349gat));
  NOR2_X1   g707(.A1(new_n906_), .A2(new_n607_), .ZN(new_n909_));
  MUX2_X1   g708(.A(G183gat), .B(new_n269_), .S(new_n909_), .Z(G1350gat));
  OAI21_X1  g709(.A(G190gat), .B1(new_n906_), .B2(new_n590_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n626_), .A2(new_n268_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n906_), .B2(new_n912_), .ZN(G1351gat));
  NOR2_X1   g712(.A1(new_n428_), .A2(new_n349_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n868_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n482_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n552_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g719(.A1(new_n915_), .A2(new_n607_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n922_));
  OR2_X1    g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  OR3_X1    g722(.A1(new_n921_), .A2(new_n922_), .A3(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n921_), .B2(new_n923_), .ZN(new_n925_));
  XOR2_X1   g724(.A(KEYINPUT63), .B(G211gat), .Z(new_n926_));
  AOI22_X1  g725(.A1(new_n924_), .A2(new_n925_), .B1(new_n921_), .B2(new_n926_), .ZN(G1354gat));
  OR3_X1    g726(.A1(new_n915_), .A2(G218gat), .A3(new_n625_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G218gat), .B1(new_n915_), .B2(new_n590_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1355gat));
endmodule


