//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_;
  INV_X1    g000(.A(KEYINPUT7), .ZN(new_n202_));
  INV_X1    g001(.A(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT8), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(new_n215_), .A3(new_n212_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G92gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT65), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G92gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n221_), .A3(G85gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT9), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n222_), .A2(KEYINPUT66), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT66), .B1(new_n222_), .B2(new_n223_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(KEYINPUT67), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(G85gat), .A2(G92gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n224_), .A2(new_n225_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n203_), .A2(KEYINPUT10), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT10), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G99gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n234_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n204_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n208_), .A2(new_n209_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n217_), .B1(new_n233_), .B2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(KEYINPUT74), .B(G29gat), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G36gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT74), .B(G29gat), .ZN(new_n246_));
  INV_X1    g045(.A(G36gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G43gat), .B(G50gat), .Z(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n245_), .A2(new_n250_), .A3(new_n248_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(KEYINPUT15), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT15), .ZN(new_n255_));
  INV_X1    g054(.A(new_n253_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n250_), .B1(new_n245_), .B2(new_n248_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n243_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(new_n253_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n260_), .B(new_n217_), .C1(new_n242_), .C2(new_n233_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G232gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT73), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT34), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n264_), .A2(KEYINPUT35), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(KEYINPUT35), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n259_), .A2(new_n261_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT77), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT77), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n259_), .A2(new_n270_), .A3(new_n261_), .A4(new_n267_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n259_), .A2(new_n261_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(KEYINPUT75), .A3(new_n265_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT75), .B1(new_n273_), .B2(new_n265_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n272_), .B(KEYINPUT76), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G190gat), .B(G218gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G134gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(G162gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n280_), .A2(KEYINPUT36), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n273_), .A2(new_n265_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n286_), .A2(new_n274_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(KEYINPUT76), .A3(new_n281_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n283_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n287_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(KEYINPUT36), .A3(new_n280_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT37), .ZN(new_n293_));
  XOR2_X1   g092(.A(G57gat), .B(G64gat), .Z(new_n294_));
  INV_X1    g093(.A(KEYINPUT11), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G57gat), .B(G64gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT11), .ZN(new_n298_));
  XOR2_X1   g097(.A(G71gat), .B(G78gat), .Z(new_n299_));
  NAND3_X1  g098(.A1(new_n296_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n298_), .A2(new_n299_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G231gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT78), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n302_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G15gat), .B(G22gat), .ZN(new_n306_));
  INV_X1    g105(.A(G1gat), .ZN(new_n307_));
  INV_X1    g106(.A(G8gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT14), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G1gat), .B(G8gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n305_), .B(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(KEYINPUT68), .B(KEYINPUT79), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT17), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT16), .B(G183gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G211gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(G127gat), .B(G155gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  OR3_X1    g119(.A1(new_n315_), .A2(new_n316_), .A3(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(KEYINPUT17), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n313_), .A2(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n323_), .A2(KEYINPUT80), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(KEYINPUT80), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n321_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT37), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n289_), .A2(new_n327_), .A3(new_n291_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n293_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G15gat), .B(G43gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT30), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G227gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G71gat), .B(G99gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G127gat), .B(G134gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G113gat), .B(G120gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT87), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n337_), .B(new_n338_), .Z(new_n341_));
  AOI21_X1  g140(.A(new_n340_), .B1(new_n341_), .B2(KEYINPUT87), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT86), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n343_), .B(KEYINPUT31), .Z(new_n344_));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT23), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(new_n347_), .B2(new_n345_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT83), .B(G183gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(G190gat), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G169gat), .ZN(new_n352_));
  INV_X1    g151(.A(G176gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT22), .B(G169gat), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n354_), .B1(new_n355_), .B2(new_n353_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT85), .B1(new_n345_), .B2(KEYINPUT23), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n347_), .A2(new_n345_), .ZN(new_n359_));
  MUX2_X1   g158(.A(KEYINPUT85), .B(new_n358_), .S(new_n359_), .Z(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT26), .B(G190gat), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n350_), .A2(KEYINPUT25), .ZN(new_n362_));
  NOR2_X1   g161(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT24), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n360_), .A2(new_n364_), .A3(new_n367_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n354_), .A2(new_n366_), .A3(new_n365_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n357_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n344_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n344_), .A2(new_n370_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n336_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n373_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n371_), .A3(new_n335_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT88), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n376_), .A3(KEYINPUT88), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G78gat), .B(G106gat), .Z(new_n382_));
  XOR2_X1   g181(.A(G211gat), .B(G218gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT94), .B(G197gat), .ZN(new_n384_));
  INV_X1    g183(.A(G204gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT95), .B(G204gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n386_), .B1(new_n388_), .B2(G197gat), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n383_), .B1(new_n389_), .B2(KEYINPUT21), .ZN(new_n390_));
  INV_X1    g189(.A(G197gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n387_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT96), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n384_), .A2(new_n385_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT97), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n390_), .B1(new_n398_), .B2(KEYINPUT21), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(KEYINPUT21), .A3(new_n383_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(G155gat), .ZN(new_n402_));
  INV_X1    g201(.A(G162gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT3), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT92), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G141gat), .A2(G148gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G141gat), .A2(G148gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT2), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n404_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n402_), .A2(new_n403_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT1), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n404_), .B2(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n415_), .A2(KEYINPUT90), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(KEYINPUT90), .ZN(new_n417_));
  INV_X1    g216(.A(new_n404_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n416_), .B(new_n417_), .C1(KEYINPUT1), .C2(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n407_), .B(KEYINPUT89), .Z(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n409_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT91), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT91), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n419_), .A2(new_n423_), .A3(new_n409_), .A4(new_n420_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n413_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n401_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G233gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT93), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n429_), .A2(G228gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(G228gat), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n428_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n427_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n433_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n382_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n434_), .A2(new_n435_), .A3(new_n382_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n425_), .A2(new_n426_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G22gat), .B(G50gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT28), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n440_), .B(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n443_), .B1(new_n436_), .B2(KEYINPUT98), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n437_), .A2(KEYINPUT98), .A3(new_n438_), .A4(new_n443_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n381_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n377_), .A3(new_n446_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n341_), .B(KEYINPUT102), .Z(new_n451_));
  AND2_X1   g250(.A1(new_n425_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n425_), .A2(new_n342_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT4), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n425_), .A2(new_n342_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT4), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G225gat), .A2(G233gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n425_), .A2(new_n451_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n455_), .A2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(new_n460_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT0), .B(G57gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(G85gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(G1gat), .B(G29gat), .Z(new_n468_));
  XOR2_X1   g267(.A(new_n467_), .B(new_n468_), .Z(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n461_), .A2(new_n465_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n459_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n469_), .B1(new_n472_), .B2(new_n464_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT27), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT18), .B(G64gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G92gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(G183gat), .A2(G190gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n360_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n356_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n348_), .A2(new_n367_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT100), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT25), .B(G183gat), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n369_), .B1(new_n361_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n486_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n487_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n484_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT105), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n484_), .A2(new_n491_), .A3(KEYINPUT105), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n494_), .A2(new_n399_), .A3(new_n400_), .A4(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n401_), .A2(new_n370_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT101), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n401_), .A2(KEYINPUT101), .A3(new_n370_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n496_), .A2(new_n499_), .A3(KEYINPUT20), .A4(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT106), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G226gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT19), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n501_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n502_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT20), .B1(new_n401_), .B2(new_n370_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT99), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n504_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n401_), .A2(new_n492_), .ZN(new_n512_));
  OAI211_X1 g311(.A(KEYINPUT99), .B(KEYINPUT20), .C1(new_n401_), .C2(new_n370_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT107), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n481_), .B1(new_n507_), .B2(new_n515_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n499_), .A2(KEYINPUT20), .A3(new_n500_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n401_), .A2(new_n492_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n518_), .A2(new_n504_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n510_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n517_), .A2(new_n519_), .B1(new_n520_), .B2(new_n504_), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n516_), .A2(KEYINPUT108), .B1(new_n480_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT108), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n523_), .B(new_n481_), .C1(new_n507_), .C2(new_n515_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n476_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n521_), .B(new_n481_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n526_), .A2(new_n476_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n450_), .B(new_n475_), .C1(new_n525_), .C2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n480_), .A2(KEYINPUT32), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n521_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n507_), .A2(new_n515_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n474_), .B(new_n530_), .C1(new_n531_), .C2(new_n529_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n461_), .A2(new_n465_), .A3(KEYINPUT33), .A4(new_n470_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT103), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n472_), .A2(new_n464_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT103), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n535_), .A2(new_n536_), .A3(KEYINPUT33), .A4(new_n470_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n470_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n539_), .B1(new_n459_), .B2(new_n463_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n526_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT33), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n471_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT104), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT104), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n471_), .A2(new_n545_), .A3(new_n542_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n532_), .B1(new_n541_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n447_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n381_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n329_), .B1(new_n528_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT13), .ZN(new_n552_));
  XOR2_X1   g351(.A(G120gat), .B(G148gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(G176gat), .B(G204gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n555_), .B(new_n556_), .Z(new_n557_));
  INV_X1    g356(.A(new_n302_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n243_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT68), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n243_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n561_), .A3(KEYINPUT12), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT12), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n243_), .B(new_n558_), .C1(new_n560_), .C2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n217_), .B(new_n302_), .C1(new_n233_), .C2(new_n242_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT69), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT69), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n570_), .A3(new_n567_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT70), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n565_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n565_), .B2(new_n572_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n567_), .B1(new_n559_), .B2(new_n566_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n557_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n574_), .A2(new_n575_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n557_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n580_), .A2(new_n577_), .A3(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n552_), .B1(new_n579_), .B2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n576_), .A2(new_n578_), .A3(new_n557_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n581_), .B1(new_n580_), .B2(new_n577_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(KEYINPUT13), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n588_), .A2(KEYINPUT72), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(KEYINPUT72), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n312_), .B1(new_n253_), .B2(new_n252_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G229gat), .A2(G233gat), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n258_), .A2(new_n254_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n312_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n594_), .B(new_n595_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n260_), .A2(new_n597_), .ZN(new_n599_));
  OAI211_X1 g398(.A(G229gat), .B(G233gat), .C1(new_n599_), .C2(new_n593_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT81), .Z(new_n602_));
  XNOR2_X1  g401(.A(G113gat), .B(G141gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n352_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(new_n391_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n605_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n598_), .A2(new_n600_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT82), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n592_), .A2(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n551_), .A2(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n614_), .A2(new_n307_), .A3(new_n474_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT109), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n616_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT38), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n292_), .B1(new_n528_), .B2(new_n550_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n622_), .A2(new_n326_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n613_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G1gat), .B1(new_n624_), .B2(new_n475_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n617_), .A2(new_n618_), .A3(KEYINPUT38), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n621_), .A2(new_n625_), .A3(new_n626_), .ZN(G1324gat));
  NOR2_X1   g426(.A1(new_n525_), .A2(new_n527_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n623_), .A2(new_n613_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(KEYINPUT110), .A2(KEYINPUT39), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(G8gat), .A3(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(KEYINPUT110), .A2(KEYINPUT39), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n614_), .A2(new_n308_), .A3(new_n628_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n632_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n629_), .A2(G8gat), .A3(new_n635_), .A4(new_n630_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n633_), .A2(new_n634_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(G1325gat));
  INV_X1    g438(.A(G15gat), .ZN(new_n640_));
  INV_X1    g439(.A(new_n381_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n614_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n623_), .A2(new_n613_), .A3(new_n641_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n643_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT41), .B1(new_n643_), .B2(G15gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n642_), .B1(new_n644_), .B2(new_n645_), .ZN(G1326gat));
  INV_X1    g445(.A(G22gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n614_), .A2(new_n647_), .A3(new_n447_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G22gat), .B1(new_n624_), .B2(new_n549_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(KEYINPUT42), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(KEYINPUT42), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n648_), .B1(new_n650_), .B2(new_n651_), .ZN(G1327gat));
  NOR3_X1   g451(.A1(new_n592_), .A2(new_n612_), .A3(new_n326_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n292_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n528_), .B2(new_n550_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n474_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n528_), .A2(new_n550_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n328_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n327_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n658_), .B1(new_n659_), .B2(new_n663_), .ZN(new_n664_));
  AOI211_X1 g463(.A(KEYINPUT43), .B(new_n662_), .C1(new_n528_), .C2(new_n550_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n653_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT44), .B(new_n653_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(new_n475_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n657_), .B1(new_n671_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g471(.A1(new_n668_), .A2(new_n628_), .A3(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G36gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n656_), .A2(new_n247_), .A3(new_n628_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT45), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n674_), .A2(KEYINPUT46), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1329gat));
  NAND2_X1  g480(.A1(new_n377_), .A2(G43gat), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n656_), .A2(new_n641_), .ZN(new_n683_));
  OAI22_X1  g482(.A1(new_n670_), .A2(new_n682_), .B1(G43gat), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g484(.A(G50gat), .B1(new_n656_), .B2(new_n447_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n670_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n447_), .A2(G50gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n686_), .B1(new_n687_), .B2(new_n688_), .ZN(G1331gat));
  NOR2_X1   g488(.A1(new_n591_), .A2(new_n611_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n623_), .A2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G57gat), .B1(new_n691_), .B2(new_n475_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n551_), .A2(new_n690_), .ZN(new_n693_));
  INV_X1    g492(.A(G57gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n474_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT111), .Z(G1332gat));
  INV_X1    g496(.A(new_n691_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n628_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G64gat), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT112), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT112), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n699_), .A2(new_n702_), .A3(G64gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n701_), .A2(KEYINPUT48), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n702_), .B1(new_n699_), .B2(G64gat), .ZN(new_n706_));
  INV_X1    g505(.A(G64gat), .ZN(new_n707_));
  AOI211_X1 g506(.A(KEYINPUT112), .B(new_n707_), .C1(new_n698_), .C2(new_n628_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n693_), .A2(new_n707_), .A3(new_n628_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n704_), .A2(new_n709_), .A3(new_n710_), .ZN(G1333gat));
  INV_X1    g510(.A(G71gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n693_), .A2(new_n712_), .A3(new_n641_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G71gat), .B1(new_n691_), .B2(new_n381_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n714_), .A2(KEYINPUT49), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(KEYINPUT49), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n713_), .B1(new_n715_), .B2(new_n716_), .ZN(G1334gat));
  INV_X1    g516(.A(G78gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n693_), .A2(new_n718_), .A3(new_n447_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G78gat), .B1(new_n691_), .B2(new_n549_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(KEYINPUT50), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(KEYINPUT50), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n719_), .B1(new_n721_), .B2(new_n722_), .ZN(G1335gat));
  NOR3_X1   g522(.A1(new_n591_), .A2(new_n611_), .A3(new_n326_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n655_), .A2(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G85gat), .B1(new_n725_), .B2(new_n474_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n664_), .A2(new_n665_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(new_n724_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(new_n474_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n726_), .B1(new_n729_), .B2(G85gat), .ZN(G1336gat));
  NAND3_X1  g529(.A1(new_n628_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT113), .Z(new_n732_));
  NAND2_X1  g531(.A1(new_n728_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n725_), .A2(new_n628_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n218_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT114), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n733_), .A2(KEYINPUT114), .A3(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1337gat));
  OAI211_X1 g539(.A(new_n725_), .B(new_n377_), .C1(new_n239_), .C2(new_n238_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n641_), .B(new_n724_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n742_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT115), .B1(new_n742_), .B2(G99gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n741_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g545(.A1(new_n725_), .A2(new_n204_), .A3(new_n447_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n447_), .B(new_n724_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(new_n749_), .A3(G106gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n748_), .B2(G106gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g552(.A1(new_n628_), .A2(new_n475_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n611_), .A2(new_n584_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n567_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT117), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n566_), .ZN(new_n762_));
  AOI211_X1 g561(.A(KEYINPUT117), .B(new_n762_), .C1(new_n562_), .C2(new_n564_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n565_), .A2(new_n572_), .A3(KEYINPUT55), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n758_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n581_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(KEYINPUT56), .A3(new_n581_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n756_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n595_), .B1(new_n599_), .B2(new_n593_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n594_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n605_), .B(new_n772_), .C1(new_n773_), .C2(new_n595_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n610_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT118), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n610_), .A2(new_n777_), .A3(new_n774_), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n585_), .A2(new_n584_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n654_), .B1(new_n771_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI211_X1 g581(.A(KEYINPUT57), .B(new_n654_), .C1(new_n771_), .C2(new_n779_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n582_), .B1(new_n778_), .B2(new_n776_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n766_), .A2(KEYINPUT56), .A3(new_n581_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT56), .B1(new_n766_), .B2(new_n581_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n784_), .B(KEYINPUT58), .C1(new_n785_), .C2(new_n786_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n663_), .A3(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n782_), .A2(new_n783_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n326_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n782_), .A2(new_n791_), .A3(KEYINPUT119), .A4(new_n783_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n794_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n329_), .A2(new_n587_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n612_), .ZN(new_n800_));
  NOR4_X1   g599(.A1(new_n329_), .A2(new_n587_), .A3(KEYINPUT116), .A4(new_n611_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n588_), .A2(new_n662_), .A3(new_n612_), .A4(new_n326_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT116), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n799_), .A2(new_n798_), .A3(new_n612_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT54), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n803_), .A2(new_n807_), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n449_), .B(new_n755_), .C1(new_n797_), .C2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(G113gat), .B1(new_n809_), .B2(new_n611_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n802_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n805_), .A2(new_n806_), .A3(KEYINPUT54), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n782_), .A2(new_n791_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT120), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT120), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n782_), .A2(new_n818_), .A3(new_n791_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n783_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n815_), .B1(new_n820_), .B2(new_n795_), .ZN(new_n821_));
  NOR4_X1   g620(.A1(new_n821_), .A2(KEYINPUT59), .A3(new_n449_), .A4(new_n755_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n812_), .A2(new_n822_), .A3(new_n612_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n810_), .B1(new_n823_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g623(.A(G120gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n591_), .B2(KEYINPUT60), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(KEYINPUT121), .Z(new_n827_));
  OAI211_X1 g626(.A(new_n809_), .B(new_n827_), .C1(KEYINPUT60), .C2(new_n825_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n812_), .A2(new_n822_), .A3(new_n591_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n825_), .ZN(G1341gat));
  AOI21_X1  g629(.A(G127gat), .B1(new_n809_), .B2(new_n326_), .ZN(new_n831_));
  INV_X1    g630(.A(G127gat), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n812_), .A2(new_n822_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n831_), .B1(new_n833_), .B2(new_n326_), .ZN(G1342gat));
  AOI21_X1  g633(.A(G134gat), .B1(new_n809_), .B2(new_n292_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n812_), .A2(new_n822_), .A3(new_n662_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(G134gat), .ZN(G1343gat));
  AOI21_X1  g636(.A(new_n448_), .B1(new_n797_), .B2(new_n808_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n754_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n612_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT122), .B(G141gat), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(G1344gat));
  INV_X1    g641(.A(new_n839_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n592_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g644(.A1(new_n839_), .A2(new_n795_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT61), .B(G155gat), .Z(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1346gat));
  NOR3_X1   g647(.A1(new_n839_), .A2(new_n403_), .A3(new_n662_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n843_), .A2(new_n292_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n403_), .B2(new_n850_), .ZN(G1347gat));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n525_), .A2(new_n474_), .A3(new_n527_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n641_), .ZN(new_n854_));
  NOR4_X1   g653(.A1(new_n821_), .A2(new_n612_), .A3(new_n447_), .A4(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n852_), .B1(new_n855_), .B2(new_n352_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n854_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n820_), .A2(new_n795_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n549_), .B(new_n857_), .C1(new_n858_), .C2(new_n815_), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT62), .B(G169gat), .C1(new_n859_), .C2(new_n612_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n855_), .A2(new_n355_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n856_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT123), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n856_), .A2(new_n860_), .A3(new_n864_), .A4(new_n861_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1348gat));
  NOR3_X1   g665(.A1(new_n821_), .A2(new_n447_), .A3(new_n854_), .ZN(new_n867_));
  AOI21_X1  g666(.A(G176gat), .B1(new_n867_), .B2(new_n592_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT124), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n447_), .B1(new_n797_), .B2(new_n808_), .ZN(new_n870_));
  AND4_X1   g669(.A1(G176gat), .A2(new_n870_), .A3(new_n592_), .A4(new_n857_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1349gat));
  NOR3_X1   g671(.A1(new_n859_), .A2(new_n488_), .A3(new_n795_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n326_), .A3(new_n857_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n349_), .B2(new_n874_), .ZN(G1350gat));
  OAI21_X1  g674(.A(G190gat), .B1(new_n859_), .B2(new_n662_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n867_), .A2(new_n292_), .A3(new_n361_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1351gat));
  NAND2_X1  g677(.A1(new_n797_), .A2(new_n808_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n448_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(new_n880_), .A3(new_n853_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n838_), .A2(KEYINPUT125), .A3(new_n853_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n611_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G197gat), .ZN(G1352gat));
  AND4_X1   g686(.A1(KEYINPUT125), .A2(new_n879_), .A3(new_n880_), .A4(new_n853_), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT125), .B1(new_n838_), .B2(new_n853_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n592_), .B(new_n388_), .C1(new_n888_), .C2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n591_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n385_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT126), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n890_), .B(new_n894_), .C1(new_n891_), .C2(new_n385_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(G1353gat));
  INV_X1    g695(.A(KEYINPUT63), .ZN(new_n897_));
  INV_X1    g696(.A(G211gat), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT127), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n795_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n885_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n901_), .ZN(new_n903_));
  AOI211_X1 g702(.A(KEYINPUT127), .B(new_n903_), .C1(new_n883_), .C2(new_n884_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n899_), .B1(new_n902_), .B2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n901_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT127), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n885_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n907_), .A2(new_n908_), .A3(new_n897_), .A4(new_n898_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n909_), .ZN(G1354gat));
  AOI21_X1  g709(.A(G218gat), .B1(new_n885_), .B2(new_n292_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n662_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(G218gat), .B2(new_n912_), .ZN(G1355gat));
endmodule


