//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  XOR2_X1   g003(.A(G211gat), .B(G218gat), .Z(new_n205_));
  INV_X1    g004(.A(KEYINPUT92), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT21), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n210_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n209_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(KEYINPUT24), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(KEYINPUT24), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G183gat), .A3(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n220_), .B1(G183gat), .B2(G190gat), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G183gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT82), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n225_), .B2(G183gat), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n219_), .B(new_n224_), .C1(new_n227_), .C2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT83), .B(G176gat), .Z(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G169gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n221_), .A2(KEYINPUT84), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n221_), .A2(KEYINPUT84), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n223_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G183gat), .A2(G190gat), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n233_), .B(new_n216_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n230_), .A2(new_n238_), .ZN(new_n239_));
  AOI211_X1 g038(.A(new_n202_), .B(new_n204_), .C1(new_n213_), .C2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n216_), .B(KEYINPUT96), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n233_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n224_), .B1(G183gat), .B2(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n236_), .A2(new_n218_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n228_), .B(KEYINPUT94), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT25), .B(G183gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n245_), .A2(new_n248_), .A3(KEYINPUT95), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT95), .B1(new_n245_), .B2(new_n248_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n212_), .B(new_n244_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n240_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT20), .B1(new_n213_), .B2(new_n239_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n244_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n254_), .B1(new_n255_), .B2(new_n213_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n204_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n253_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G64gat), .B(G92gat), .Z(new_n259_));
  XNOR2_X1  g058(.A(G8gat), .B(G36gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n258_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n263_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n253_), .B(new_n265_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT27), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n230_), .A2(new_n238_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n202_), .B1(new_n271_), .B2(new_n212_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n244_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n245_), .A2(new_n248_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT95), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n273_), .B1(new_n276_), .B2(new_n249_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n272_), .B1(new_n277_), .B2(new_n212_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n278_), .A2(new_n204_), .B1(new_n252_), .B2(new_n240_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n270_), .B1(new_n279_), .B2(new_n265_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n278_), .A2(new_n204_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n274_), .A2(new_n244_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT101), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n274_), .A2(KEYINPUT101), .A3(new_n244_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n212_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n202_), .B1(new_n213_), .B2(new_n239_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n257_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n263_), .B1(new_n281_), .B2(new_n288_), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n267_), .A2(new_n269_), .B1(new_n280_), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G71gat), .B(G99gat), .ZN(new_n291_));
  INV_X1    g090(.A(G15gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT30), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n239_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G127gat), .B(G134gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G113gat), .B(G120gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT86), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT31), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n295_), .B(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(KEYINPUT85), .B(G43gat), .Z(new_n302_));
  NAND2_X1  g101(.A1(G227gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n301_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT89), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n309_), .A2(KEYINPUT3), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(KEYINPUT3), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT2), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n311_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT88), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT88), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(G155gat), .A3(G162gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT87), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n314_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n312_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(new_n307_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n319_), .A2(KEYINPUT1), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n321_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n319_), .A2(KEYINPUT1), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n324_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n306_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n329_));
  OAI211_X1 g128(.A(G228gat), .B(G233gat), .C1(new_n329_), .C2(new_n212_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n322_), .A2(new_n328_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT90), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n322_), .A2(new_n328_), .A3(KEYINPUT90), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n306_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G228gat), .A2(G233gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n213_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n330_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G78gat), .B(G106gat), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT93), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n339_), .B(new_n330_), .C1(new_n335_), .C2(new_n337_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n343_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(new_n341_), .A3(KEYINPUT93), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n333_), .A2(new_n334_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT28), .B1(new_n347_), .B2(KEYINPUT29), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n333_), .A2(new_n349_), .A3(new_n306_), .A4(new_n334_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G22gat), .B(G50gat), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n351_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT91), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n348_), .A2(new_n350_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n351_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT91), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n344_), .A2(new_n346_), .B1(new_n354_), .B2(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n357_), .A2(new_n341_), .A3(new_n343_), .A4(new_n359_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n290_), .B(new_n305_), .C1(new_n361_), .C2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n288_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n256_), .A2(new_n257_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n265_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n266_), .A2(KEYINPUT27), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n268_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT103), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n279_), .A2(new_n265_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n266_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n269_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n280_), .A2(new_n289_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT103), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n371_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n344_), .A2(new_n346_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n354_), .A2(new_n360_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n301_), .B(new_n304_), .Z(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n362_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n364_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n299_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n347_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n299_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n322_), .A2(new_n328_), .A3(new_n298_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT4), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n385_), .B1(new_n389_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n387_), .A2(new_n391_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n385_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(G57gat), .B(G85gat), .Z(new_n399_));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n401_), .B(new_n402_), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n398_), .A2(new_n404_), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n394_), .A2(new_n397_), .A3(new_n403_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n384_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n381_), .A2(new_n362_), .A3(new_n305_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n389_), .A2(new_n393_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT100), .B1(new_n410_), .B2(new_n385_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n403_), .B1(new_n395_), .B2(new_n385_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(KEYINPUT100), .A3(new_n385_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n267_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n398_), .A2(new_n404_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(KEYINPUT99), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT99), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT33), .B1(new_n406_), .B2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n415_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n265_), .A2(KEYINPUT32), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n279_), .A2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n281_), .A2(new_n288_), .ZN(new_n424_));
  OAI221_X1 g223(.A(new_n423_), .B1(new_n424_), .B2(new_n422_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n409_), .B1(new_n421_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n408_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G134gat), .B(G162gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT77), .ZN(new_n430_));
  XOR2_X1   g229(.A(G190gat), .B(G218gat), .Z(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n432_), .A2(KEYINPUT36), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT8), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT69), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n436_), .B1(G99gat), .B2(G106gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G99gat), .A2(G106gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(KEYINPUT6), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n435_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(KEYINPUT6), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n436_), .A2(G99gat), .A3(G106gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(KEYINPUT69), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n444_));
  INV_X1    g243(.A(G99gat), .ZN(new_n445_));
  INV_X1    g244(.A(G106gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n440_), .A2(new_n443_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(G85gat), .ZN(new_n451_));
  INV_X1    g250(.A(G92gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G85gat), .A2(G92gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n434_), .B1(new_n450_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n441_), .A2(new_n442_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n447_), .A2(new_n448_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n434_), .B(new_n456_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT70), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT70), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT69), .B1(new_n441_), .B2(new_n442_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n465_), .A2(new_n460_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n455_), .B1(new_n466_), .B2(new_n443_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n464_), .B(new_n461_), .C1(new_n467_), .C2(new_n434_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n463_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT71), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT68), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT10), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n472_), .A2(G99gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n445_), .A2(KEYINPUT10), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT64), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n445_), .A2(KEYINPUT10), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(G99gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT64), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT65), .B(G106gat), .Z(new_n481_));
  AOI21_X1  g280(.A(new_n459_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT66), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n454_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT67), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n485_), .A3(KEYINPUT9), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT67), .B1(new_n454_), .B2(new_n483_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT9), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n488_), .B1(new_n454_), .B2(KEYINPUT67), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n486_), .B(new_n453_), .C1(new_n487_), .C2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n471_), .B1(new_n482_), .B2(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n478_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n481_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  AND4_X1   g293(.A1(new_n471_), .A2(new_n494_), .A3(new_n490_), .A4(new_n458_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n470_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n482_), .A2(new_n471_), .A3(new_n490_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n490_), .A3(new_n458_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT68), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(new_n499_), .A3(KEYINPUT71), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n469_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT15), .ZN(new_n502_));
  INV_X1    g301(.A(G29gat), .ZN(new_n503_));
  INV_X1    g302(.A(G36gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G29gat), .A2(G36gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(G43gat), .A2(G50gat), .ZN(new_n508_));
  NOR2_X1   g307(.A1(G43gat), .A2(G50gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n505_), .B(new_n506_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n512_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n502_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n513_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n512_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(KEYINPUT15), .A3(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n501_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n497_), .A2(new_n499_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n457_), .A2(new_n462_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n519_), .A2(new_n520_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G232gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n523_), .A2(KEYINPUT76), .A3(new_n528_), .A4(new_n531_), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n501_), .A2(new_n522_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n532_), .B1(KEYINPUT35), .B2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n531_), .B1(new_n533_), .B2(KEYINPUT76), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n433_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n531_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n523_), .A2(new_n528_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT76), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n432_), .B(KEYINPUT36), .Z(new_n543_));
  NAND4_X1  g342(.A1(new_n540_), .A2(new_n542_), .A3(new_n532_), .A4(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n536_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G15gat), .B(G22gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G1gat), .A2(G8gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT14), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(G1gat), .A2(G8gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n547_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n546_), .A2(new_n547_), .A3(new_n550_), .A4(new_n548_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n557_), .A2(KEYINPUT11), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(KEYINPUT11), .ZN(new_n559_));
  XOR2_X1   g358(.A(G71gat), .B(G78gat), .Z(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n559_), .A2(new_n560_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n556_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(G211gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT16), .B(G183gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(KEYINPUT80), .A3(KEYINPUT17), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n564_), .B(new_n569_), .C1(KEYINPUT17), .C2(new_n568_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n563_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n461_), .B1(new_n467_), .B2(new_n434_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n576_), .A2(new_n497_), .A3(new_n499_), .A4(new_n563_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT12), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n563_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n501_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n575_), .A2(new_n582_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT72), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n577_), .A2(new_n587_), .A3(new_n579_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n587_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n581_), .B1(new_n586_), .B2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G120gat), .B(G148gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(G204gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT5), .B(G176gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n593_), .B(new_n594_), .Z(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n581_), .B(new_n595_), .C1(new_n586_), .C2(new_n590_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT13), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n597_), .A2(KEYINPUT13), .A3(new_n598_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT81), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n516_), .A2(new_n521_), .A3(new_n554_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n554_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n604_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n605_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n554_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n527_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n609_), .B1(new_n611_), .B2(new_n606_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G169gat), .B(G197gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n608_), .A2(new_n612_), .A3(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n616_), .B1(new_n608_), .B2(new_n612_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n603_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n608_), .A2(new_n612_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(new_n615_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n608_), .A2(new_n612_), .A3(new_n616_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(KEYINPUT81), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n619_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n602_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n428_), .A2(new_n545_), .A3(new_n573_), .A4(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G1gat), .B1(new_n627_), .B2(new_n407_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n426_), .B1(new_n384_), .B2(new_n407_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT37), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n536_), .A2(new_n631_), .A3(new_n544_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT78), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n536_), .A2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(KEYINPUT78), .B(new_n433_), .C1(new_n534_), .C2(new_n535_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n544_), .A2(KEYINPUT79), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n523_), .A2(KEYINPUT76), .A3(new_n528_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n637_), .A2(new_n531_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT79), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n540_), .A4(new_n543_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .A4(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n632_), .B1(new_n641_), .B2(KEYINPUT37), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n630_), .A2(new_n642_), .A3(new_n572_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n600_), .A2(new_n601_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT73), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT73), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n602_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n625_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n643_), .A2(new_n644_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n642_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n428_), .A2(new_n651_), .A3(new_n573_), .A4(new_n649_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT104), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(G1gat), .ZN(new_n655_));
  INV_X1    g454(.A(new_n407_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n654_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(KEYINPUT105), .A3(new_n629_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT105), .B1(new_n657_), .B2(new_n629_), .ZN(new_n659_));
  OAI221_X1 g458(.A(new_n628_), .B1(new_n629_), .B2(new_n657_), .C1(new_n658_), .C2(new_n659_), .ZN(G1324gat));
  INV_X1    g459(.A(new_n378_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G8gat), .B1(new_n627_), .B2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT39), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n661_), .A2(G8gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n654_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n665_), .ZN(new_n667_));
  AOI211_X1 g466(.A(KEYINPUT106), .B(new_n667_), .C1(new_n650_), .C2(new_n653_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n663_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n663_), .B(KEYINPUT40), .C1(new_n666_), .C2(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1325gat));
  OAI21_X1  g472(.A(G15gat), .B1(new_n627_), .B2(new_n305_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(KEYINPUT41), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(KEYINPUT41), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n382_), .A2(new_n292_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n675_), .B(new_n676_), .C1(new_n652_), .C2(new_n677_), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n361_), .A2(new_n363_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G22gat), .B1(new_n627_), .B2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT42), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n679_), .A2(G22gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n652_), .B2(new_n682_), .ZN(G1327gat));
  NOR3_X1   g482(.A1(new_n630_), .A2(new_n545_), .A3(new_n573_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n626_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(new_n503_), .A3(new_n656_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n688_), .A2(KEYINPUT43), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(KEYINPUT43), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n689_), .B(new_n690_), .C1(new_n630_), .C2(new_n651_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n428_), .A2(new_n688_), .A3(KEYINPUT43), .A4(new_n642_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n572_), .B1(KEYINPUT108), .B2(KEYINPUT44), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n602_), .A2(new_n625_), .A3(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n691_), .A2(new_n692_), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n691_), .A2(new_n692_), .A3(new_n696_), .A4(new_n694_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n656_), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT109), .B1(new_n701_), .B2(G29gat), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703_));
  AOI211_X1 g502(.A(new_n703_), .B(new_n503_), .C1(new_n700_), .C2(new_n656_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n687_), .B1(new_n702_), .B2(new_n704_), .ZN(G1328gat));
  NOR2_X1   g504(.A1(new_n661_), .A2(G36gat), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OR3_X1    g506(.A1(new_n685_), .A2(KEYINPUT45), .A3(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT45), .B1(new_n685_), .B2(new_n707_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n661_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(new_n504_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n710_), .B(KEYINPUT46), .C1(new_n711_), .C2(new_n504_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1329gat));
  AOI21_X1  g515(.A(G43gat), .B1(new_n686_), .B2(new_n382_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n382_), .A2(G43gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n700_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(G1330gat));
  OR3_X1    g520(.A1(new_n685_), .A2(G50gat), .A3(new_n679_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n679_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G50gat), .B1(new_n723_), .B2(new_n724_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(G1331gat));
  NAND3_X1  g526(.A1(new_n646_), .A2(new_n648_), .A3(new_n625_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n545_), .ZN(new_n729_));
  NOR4_X1   g528(.A1(new_n630_), .A2(new_n728_), .A3(new_n729_), .A4(new_n572_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(G57gat), .A3(new_n656_), .ZN(new_n731_));
  INV_X1    g530(.A(G57gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n643_), .A2(new_n602_), .A3(new_n625_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n407_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n731_), .B1(new_n734_), .B2(KEYINPUT111), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(KEYINPUT111), .B2(new_n734_), .ZN(G1332gat));
  OR3_X1    g535(.A1(new_n733_), .A2(G64gat), .A3(new_n661_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n730_), .A2(new_n378_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G64gat), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(KEYINPUT48), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(KEYINPUT48), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(G1333gat));
  OR3_X1    g541(.A1(new_n733_), .A2(G71gat), .A3(new_n305_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n730_), .A2(new_n382_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n744_), .A2(G71gat), .A3(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n744_), .B2(G71gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT113), .ZN(G1334gat));
  OR3_X1    g548(.A1(new_n733_), .A2(G78gat), .A3(new_n679_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n679_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n730_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G78gat), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(KEYINPUT50), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(KEYINPUT50), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n750_), .B1(new_n754_), .B2(new_n755_), .ZN(G1335gat));
  INV_X1    g555(.A(new_n728_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n684_), .A2(new_n757_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n758_), .A2(G85gat), .A3(new_n407_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n645_), .A2(new_n573_), .A3(new_n624_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n691_), .A2(new_n692_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n656_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n759_), .B1(new_n762_), .B2(G85gat), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT114), .ZN(G1336gat));
  INV_X1    g563(.A(new_n758_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G92gat), .B1(new_n765_), .B2(new_n378_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n661_), .A2(new_n452_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n761_), .B2(new_n767_), .ZN(G1337gat));
  NAND3_X1  g567(.A1(new_n765_), .A2(new_n480_), .A3(new_n382_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n761_), .A2(new_n382_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(new_n445_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n765_), .A2(new_n481_), .A3(new_n751_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n691_), .A2(new_n692_), .A3(new_n751_), .A4(new_n760_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(G106gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G106gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g578(.A(G113gat), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n598_), .A2(new_n624_), .A3(KEYINPUT117), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT117), .B1(new_n598_), .B2(new_n624_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n586_), .B2(new_n590_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n501_), .A2(new_n583_), .B1(new_n575_), .B2(new_n582_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n787_), .B(KEYINPUT55), .C1(new_n589_), .C2(new_n588_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n584_), .A2(new_n577_), .A3(new_n585_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n580_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n786_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n791_), .A2(KEYINPUT56), .A3(new_n596_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT56), .B1(new_n791_), .B2(new_n596_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n784_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n604_), .A2(new_n609_), .A3(new_n607_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n605_), .B1(new_n611_), .B2(new_n606_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n615_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n622_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n729_), .B1(new_n794_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n781_), .B1(new_n801_), .B2(KEYINPUT57), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n791_), .A2(new_n596_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n791_), .A2(KEYINPUT56), .A3(new_n596_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n799_), .B1(new_n808_), .B2(new_n784_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT118), .B(new_n803_), .C1(new_n809_), .C2(new_n729_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n794_), .A2(new_n800_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT57), .A3(new_n545_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n598_), .A2(new_n622_), .A3(new_n797_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n815_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n808_), .A2(new_n817_), .A3(new_n813_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n642_), .A2(new_n816_), .A3(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n802_), .A2(new_n810_), .A3(new_n812_), .A4(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n819_), .A2(new_n812_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n823_), .A2(KEYINPUT120), .A3(new_n810_), .A4(new_n802_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(new_n824_), .A3(new_n572_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n625_), .A2(new_n573_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT115), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n828_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n651_), .A2(new_n826_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT116), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n651_), .A2(new_n829_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT54), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n651_), .A2(new_n829_), .A3(new_n834_), .A4(new_n826_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n831_), .A2(new_n833_), .A3(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n825_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n378_), .A2(new_n383_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n656_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n780_), .B1(new_n841_), .B2(new_n625_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n819_), .A2(new_n812_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n801_), .A2(KEYINPUT57), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n572_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n836_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n840_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n625_), .A2(new_n780_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n839_), .B1(new_n825_), .B2(new_n836_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n848_), .B(new_n849_), .C1(new_n850_), .C2(new_n847_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n842_), .A2(new_n851_), .ZN(G1340gat));
  NAND2_X1  g651(.A1(new_n646_), .A2(new_n648_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n854_), .B(new_n848_), .C1(new_n850_), .C2(new_n847_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G120gat), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n645_), .A2(KEYINPUT60), .ZN(new_n857_));
  MUX2_X1   g656(.A(new_n857_), .B(KEYINPUT60), .S(G120gat), .Z(new_n858_));
  NAND2_X1  g657(.A1(new_n850_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n856_), .A2(new_n859_), .ZN(G1341gat));
  INV_X1    g659(.A(G127gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n841_), .B2(new_n572_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n572_), .A2(new_n861_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n848_), .B(new_n863_), .C1(new_n850_), .C2(new_n847_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1342gat));
  INV_X1    g664(.A(G134gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n841_), .B2(new_n545_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n651_), .A2(new_n866_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n848_), .B(new_n868_), .C1(new_n850_), .C2(new_n847_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n867_), .A2(new_n869_), .ZN(G1343gat));
  NOR2_X1   g669(.A1(new_n679_), .A2(new_n382_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n661_), .A3(new_n656_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT121), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n837_), .A2(new_n624_), .A3(new_n873_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g674(.A1(new_n837_), .A2(new_n854_), .A3(new_n873_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g676(.A1(new_n836_), .A2(new_n572_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n873_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1346gat));
  AND2_X1   g680(.A1(new_n837_), .A2(new_n873_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n729_), .ZN(new_n883_));
  INV_X1    g682(.A(G162gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n651_), .A2(new_n884_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n883_), .A2(new_n884_), .B1(new_n882_), .B2(new_n885_), .ZN(G1347gat));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n661_), .A2(new_n656_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n383_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  AOI211_X1 g689(.A(new_n625_), .B(new_n890_), .C1(new_n836_), .C2(new_n845_), .ZN(new_n891_));
  OAI21_X1  g690(.A(G169gat), .B1(new_n891_), .B2(KEYINPUT122), .ZN(new_n892_));
  INV_X1    g691(.A(new_n890_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n846_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n894_), .A2(new_n895_), .A3(new_n625_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n887_), .B1(new_n892_), .B2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n895_), .B1(new_n894_), .B2(new_n625_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n891_), .A2(KEYINPUT122), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n898_), .A2(new_n899_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n891_), .A2(new_n232_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n897_), .A2(new_n900_), .A3(new_n901_), .ZN(G1348gat));
  INV_X1    g701(.A(new_n894_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n602_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n893_), .A2(G176gat), .A3(new_n854_), .ZN(new_n905_));
  AOI22_X1  g704(.A1(new_n904_), .A2(new_n231_), .B1(new_n837_), .B2(new_n905_), .ZN(G1349gat));
  AOI21_X1  g705(.A(G183gat), .B1(new_n878_), .B2(new_n893_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n572_), .A2(new_n247_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n903_), .B2(new_n908_), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n894_), .B2(new_n651_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n729_), .A2(new_n246_), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n911_), .B(KEYINPUT123), .Z(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n894_), .B2(new_n912_), .ZN(G1351gat));
  NAND2_X1  g712(.A1(new_n888_), .A2(new_n871_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n837_), .A2(G197gat), .A3(new_n624_), .A4(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n837_), .A2(new_n624_), .A3(new_n915_), .ZN(new_n919_));
  INV_X1    g718(.A(G197gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n914_), .B1(new_n825_), .B2(new_n836_), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n922_), .A2(KEYINPUT124), .A3(G197gat), .A4(new_n624_), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n918_), .A2(new_n921_), .A3(new_n923_), .ZN(G1352gat));
  NOR2_X1   g723(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n925_));
  AND2_X1   g724(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n922_), .B(new_n854_), .C1(new_n925_), .C2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n837_), .A2(new_n915_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n853_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n927_), .B1(new_n929_), .B2(new_n925_), .ZN(G1353gat));
  AOI211_X1 g729(.A(KEYINPUT63), .B(G211gat), .C1(new_n922_), .C2(new_n573_), .ZN(new_n931_));
  OR2_X1    g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n572_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n933_));
  AND3_X1   g732(.A1(new_n922_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n931_), .A2(new_n934_), .ZN(G1354gat));
  AND3_X1   g734(.A1(new_n922_), .A2(G218gat), .A3(new_n642_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n837_), .A2(new_n729_), .A3(new_n915_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n938_));
  AOI21_X1  g737(.A(G218gat), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n922_), .A2(KEYINPUT126), .A3(new_n729_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n936_), .B1(new_n939_), .B2(new_n940_), .ZN(G1355gat));
endmodule


