//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n613_, new_n614_, new_n615_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NOR2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n205_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT8), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT10), .B(G99gat), .Z(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  AOI22_X1  g011(.A1(KEYINPUT9), .A2(new_n202_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  NOR3_X1   g014(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT9), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n208_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n210_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G57gat), .B(G64gat), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n220_), .A2(KEYINPUT11), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(KEYINPUT11), .ZN(new_n222_));
  XOR2_X1   g021(.A(G71gat), .B(G78gat), .Z(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n222_), .A2(new_n223_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n219_), .B(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT12), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT12), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n219_), .A2(new_n229_), .A3(new_n225_), .A4(new_n224_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G230gat), .A2(G233gat), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n227_), .A2(new_n232_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G120gat), .B(G148gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(G176gat), .B(G204gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT64), .B(KEYINPUT5), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT65), .B1(new_n235_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n240_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n241_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT13), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G29gat), .B(G36gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT66), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G43gat), .B(G50gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n249_), .A2(KEYINPUT66), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n249_), .A2(KEYINPUT66), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(new_n251_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G232gat), .A2(G233gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT34), .ZN(new_n259_));
  OAI22_X1  g058(.A1(new_n219_), .A2(new_n257_), .B1(KEYINPUT35), .B2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n257_), .B(KEYINPUT15), .Z(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(new_n219_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n263_));
  OAI211_X1 g062(.A(KEYINPUT35), .B(new_n259_), .C1(new_n260_), .C2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n262_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G190gat), .B(G218gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT68), .ZN(new_n267_));
  XOR2_X1   g066(.A(G134gat), .B(G162gat), .Z(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(KEYINPUT36), .Z(new_n270_));
  AND2_X1   g069(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n269_), .A2(KEYINPUT36), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n265_), .A2(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT37), .ZN(new_n275_));
  OR3_X1    g074(.A1(new_n271_), .A2(new_n273_), .A3(KEYINPUT37), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G15gat), .B(G22gat), .ZN(new_n278_));
  INV_X1    g077(.A(G1gat), .ZN(new_n279_));
  INV_X1    g078(.A(G8gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT14), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G1gat), .B(G8gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n226_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G231gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT17), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G127gat), .B(G155gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT16), .ZN(new_n291_));
  XOR2_X1   g090(.A(G183gat), .B(G211gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n288_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(KEYINPUT17), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n294_), .B1(new_n288_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT69), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT70), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n277_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n248_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G78gat), .B(G106gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT88), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304_));
  NOR2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT78), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n307_), .A2(KEYINPUT79), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT79), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n309_), .A2(KEYINPUT78), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n306_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(KEYINPUT78), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n307_), .A2(KEYINPUT79), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n305_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(KEYINPUT1), .Z(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  AND3_X1   g117(.A1(KEYINPUT77), .A2(G141gat), .A3(G148gat), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT77), .B1(G141gat), .B2(G148gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  NOR3_X1   g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT83), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n312_), .A2(new_n313_), .A3(new_n305_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n305_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n316_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT82), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  OAI211_X1 g128(.A(KEYINPUT82), .B(new_n316_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(G141gat), .ZN(new_n332_));
  INV_X1    g131(.A(G148gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT2), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT2), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT81), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(KEYINPUT80), .B2(KEYINPUT3), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n332_), .A2(new_n333_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT81), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n338_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n321_), .B(new_n337_), .C1(KEYINPUT80), .C2(KEYINPUT3), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n334_), .A2(new_n336_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n324_), .B1(new_n331_), .B2(new_n345_), .ZN(new_n346_));
  AOI211_X1 g145(.A(KEYINPUT83), .B(new_n344_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n304_), .B(new_n323_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT28), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT82), .B1(new_n315_), .B2(new_n316_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n316_), .ZN(new_n351_));
  AOI211_X1 g150(.A(new_n328_), .B(new_n351_), .C1(new_n311_), .C2(new_n314_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n345_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT83), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n331_), .A2(new_n324_), .A3(new_n345_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT28), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n356_), .A2(new_n357_), .A3(new_n304_), .A4(new_n323_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n349_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n349_), .B2(new_n358_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n303_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n323_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n357_), .B1(new_n365_), .B2(new_n304_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n348_), .A2(KEYINPUT28), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n359_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n301_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n349_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G211gat), .B(G218gat), .Z(new_n372_));
  INV_X1    g171(.A(G204gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G197gat), .ZN(new_n374_));
  INV_X1    g173(.A(G197gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(G204gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n372_), .A2(KEYINPUT21), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT85), .B1(new_n377_), .B2(KEYINPUT21), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT85), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT21), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n374_), .A2(new_n376_), .A3(new_n381_), .A4(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT84), .B1(new_n375_), .B2(G204gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT84), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n373_), .A3(G197gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n387_), .A3(new_n376_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n372_), .B1(new_n388_), .B2(KEYINPUT21), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n384_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n384_), .A2(new_n389_), .A3(KEYINPUT86), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n379_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n323_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n394_), .B1(new_n395_), .B2(KEYINPUT29), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT87), .ZN(new_n397_));
  OAI211_X1 g196(.A(G228gat), .B(G233gat), .C1(new_n394_), .C2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n396_), .B(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n363_), .A2(new_n371_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(new_n363_), .B2(new_n371_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT27), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n406_), .B(KEYINPUT90), .Z(new_n407_));
  AND3_X1   g206(.A1(new_n384_), .A2(new_n389_), .A3(KEYINPUT86), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT86), .B1(new_n384_), .B2(new_n389_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n378_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G183gat), .A2(G190gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT23), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT23), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(G183gat), .A3(G190gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(G183gat), .A2(G190gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(G169gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT25), .B(G183gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT26), .B(G190gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT24), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(G169gat), .B2(G176gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(G169gat), .B2(G176gat), .ZN(new_n427_));
  INV_X1    g226(.A(G169gat), .ZN(new_n428_));
  INV_X1    g227(.A(G176gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n425_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n424_), .A2(new_n427_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n414_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT73), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n412_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n411_), .A2(KEYINPUT73), .A3(KEYINPUT23), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n432_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n421_), .B1(new_n431_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT20), .B1(new_n410_), .B2(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n436_), .A2(new_n416_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n431_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n439_), .A2(new_n420_), .B1(new_n440_), .B2(new_n415_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n394_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n407_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G8gat), .B(G36gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G64gat), .B(G92gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n394_), .A2(new_n441_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n410_), .A2(new_n437_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n406_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(KEYINPUT20), .A4(new_n451_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n443_), .A2(new_n448_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n448_), .B1(new_n443_), .B2(new_n452_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n403_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n443_), .A2(new_n448_), .A3(new_n452_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n438_), .A2(new_n442_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n407_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n449_), .A2(new_n450_), .A3(KEYINPUT20), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n457_), .A2(new_n458_), .B1(new_n459_), .B2(new_n406_), .ZN(new_n460_));
  OAI211_X1 g259(.A(KEYINPUT27), .B(new_n456_), .C1(new_n460_), .C2(new_n448_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n455_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n402_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G127gat), .B(G134gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G113gat), .B(G120gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n464_), .B(new_n465_), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n365_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n395_), .A2(new_n466_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT4), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n471_), .B(KEYINPUT92), .Z(new_n472_));
  INV_X1    g271(.A(KEYINPUT94), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n467_), .B1(new_n356_), .B2(new_n323_), .ZN(new_n474_));
  XOR2_X1   g273(.A(KEYINPUT93), .B(KEYINPUT4), .Z(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n473_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  NOR4_X1   g276(.A1(new_n365_), .A2(KEYINPUT94), .A3(new_n467_), .A4(new_n475_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n470_), .B(new_n472_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n468_), .A2(new_n469_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n471_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G1gat), .B(G29gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(G85gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT0), .B(G57gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n483_), .B(new_n484_), .Z(new_n485_));
  AND3_X1   g284(.A1(new_n479_), .A2(new_n481_), .A3(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT75), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT74), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G227gat), .A2(G233gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(G15gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(G43gat), .ZN(new_n494_));
  INV_X1    g293(.A(G15gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n492_), .B(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(G43gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G71gat), .B(G99gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n494_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n500_), .B1(new_n494_), .B2(new_n498_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n491_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT30), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n437_), .A2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n421_), .B(KEYINPUT30), .C1(new_n431_), .C2(new_n436_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n504_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n503_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(KEYINPUT74), .A3(new_n501_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n490_), .B1(new_n508_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT31), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n510_), .A2(new_n504_), .A3(new_n506_), .A4(new_n507_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n513_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n467_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n508_), .A2(new_n511_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(new_n514_), .A3(KEYINPUT75), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT31), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(new_n515_), .A3(new_n466_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n463_), .A2(new_n489_), .A3(new_n523_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n518_), .A2(KEYINPUT76), .A3(new_n522_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT76), .B1(new_n518_), .B2(new_n522_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n479_), .A2(new_n481_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n485_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n479_), .A2(new_n481_), .A3(new_n485_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n462_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n399_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n361_), .A2(new_n362_), .A3(new_n301_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n302_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n363_), .A2(new_n371_), .A3(new_n399_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n527_), .B1(new_n532_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT33), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n531_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n443_), .A2(new_n452_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n448_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n456_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n471_), .B(new_n470_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n485_), .B1(new_n480_), .B2(new_n472_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n479_), .A2(KEYINPUT33), .A3(new_n481_), .A4(new_n485_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n541_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n448_), .A2(KEYINPUT32), .ZN(new_n551_));
  MUX2_X1   g350(.A(new_n460_), .B(new_n542_), .S(new_n551_), .Z(new_n552_));
  OAI21_X1  g351(.A(new_n552_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n550_), .A2(new_n402_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n539_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT95), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT95), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n539_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n524_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT71), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n257_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(new_n284_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G229gat), .A2(G233gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n561_), .A2(new_n284_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n261_), .A2(new_n284_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n563_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G113gat), .B(G141gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(G169gat), .B(G197gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n569_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n559_), .A2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n300_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(new_n279_), .A3(new_n489_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT38), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT96), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n248_), .A2(new_n576_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n297_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n274_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n559_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(G1gat), .B1(new_n588_), .B2(new_n488_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n582_), .B(new_n589_), .C1(new_n580_), .C2(new_n579_), .ZN(G1324gat));
  INV_X1    g389(.A(new_n578_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n591_), .A2(G8gat), .A3(new_n462_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n462_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n585_), .A2(new_n593_), .A3(new_n587_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT97), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n585_), .A2(new_n596_), .A3(new_n593_), .A4(new_n587_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n597_), .A3(G8gat), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT39), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n595_), .A2(new_n597_), .A3(new_n600_), .A4(G8gat), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n592_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n602_), .B(new_n604_), .ZN(G1325gat));
  INV_X1    g404(.A(new_n527_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G15gat), .B1(new_n588_), .B2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT99), .Z(new_n608_));
  OR2_X1    g407(.A1(new_n608_), .A2(KEYINPUT41), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(KEYINPUT41), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n578_), .A2(new_n495_), .A3(new_n527_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .ZN(G1326gat));
  OAI21_X1  g411(.A(G22gat), .B1(new_n588_), .B2(new_n402_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT42), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n402_), .A2(G22gat), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n614_), .B1(new_n591_), .B2(new_n615_), .ZN(G1327gat));
  INV_X1    g415(.A(new_n298_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n586_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n248_), .A2(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n619_), .A2(new_n577_), .ZN(new_n620_));
  AOI21_X1  g419(.A(G29gat), .B1(new_n620_), .B2(new_n489_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT44), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n559_), .A2(KEYINPUT43), .A3(new_n277_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n275_), .A2(KEYINPUT100), .A3(new_n276_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT100), .B1(new_n275_), .B2(new_n276_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT43), .B1(new_n559_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT101), .ZN(new_n628_));
  INV_X1    g427(.A(new_n524_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n539_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n557_), .B1(new_n539_), .B2(new_n554_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n629_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n277_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n275_), .A2(KEYINPUT100), .A3(new_n276_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n632_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(KEYINPUT43), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n623_), .B1(new_n628_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n583_), .A2(new_n617_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n622_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n623_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n638_), .B1(new_n637_), .B2(KEYINPUT43), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT43), .ZN(new_n645_));
  AOI211_X1 g444(.A(KEYINPUT101), .B(new_n645_), .C1(new_n632_), .C2(new_n636_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n643_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n641_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(KEYINPUT44), .A3(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n642_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n489_), .A2(G29gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n621_), .B1(new_n650_), .B2(new_n651_), .ZN(G1328gat));
  INV_X1    g451(.A(new_n620_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n653_), .A2(G36gat), .A3(new_n462_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT45), .Z(new_n655_));
  NAND3_X1  g454(.A1(new_n642_), .A2(new_n593_), .A3(new_n649_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n656_), .A2(new_n657_), .A3(G36gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n656_), .B2(G36gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI221_X1 g461(.A(new_n655_), .B1(KEYINPUT103), .B2(KEYINPUT46), .C1(new_n658_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1329gat));
  INV_X1    g463(.A(new_n523_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n650_), .A2(G43gat), .A3(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n497_), .B1(new_n653_), .B2(new_n606_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(G1330gat));
  AOI21_X1  g469(.A(G50gat), .B1(new_n620_), .B2(new_n538_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n538_), .A2(G50gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n650_), .B2(new_n672_), .ZN(G1331gat));
  INV_X1    g472(.A(new_n248_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(new_n299_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT105), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n559_), .A2(new_n575_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G57gat), .B1(new_n678_), .B2(new_n489_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n674_), .A2(new_n575_), .A3(new_n617_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n587_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(G57gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n489_), .B2(KEYINPUT106), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(KEYINPUT106), .B2(new_n683_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n679_), .B1(new_n682_), .B2(new_n685_), .ZN(G1332gat));
  OAI21_X1  g485(.A(G64gat), .B1(new_n681_), .B2(new_n462_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT48), .ZN(new_n688_));
  INV_X1    g487(.A(G64gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n678_), .A2(new_n689_), .A3(new_n593_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1333gat));
  OAI21_X1  g490(.A(G71gat), .B1(new_n681_), .B2(new_n606_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT49), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n606_), .A2(G71gat), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT107), .Z(new_n695_));
  NAND2_X1  g494(.A1(new_n678_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT108), .ZN(G1334gat));
  OAI21_X1  g497(.A(G78gat), .B1(new_n681_), .B2(new_n402_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT50), .ZN(new_n700_));
  INV_X1    g499(.A(G78gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n678_), .A2(new_n701_), .A3(new_n538_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1335gat));
  NOR4_X1   g502(.A1(new_n674_), .A2(new_n575_), .A3(new_n559_), .A4(new_n618_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G85gat), .B1(new_n704_), .B2(new_n489_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT109), .Z(new_n706_));
  NOR3_X1   g505(.A1(new_n674_), .A2(new_n575_), .A3(new_n298_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n647_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n488_), .A2(new_n214_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n706_), .B1(new_n710_), .B2(new_n711_), .ZN(G1336gat));
  XNOR2_X1  g511(.A(new_n708_), .B(KEYINPUT110), .ZN(new_n713_));
  OAI21_X1  g512(.A(G92gat), .B1(new_n713_), .B2(new_n462_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n704_), .A2(new_n215_), .A3(new_n593_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1337gat));
  INV_X1    g515(.A(G99gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n710_), .B2(new_n527_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n704_), .A2(new_n665_), .A3(new_n211_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT51), .B1(new_n718_), .B2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G99gat), .B1(new_n713_), .B2(new_n606_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT51), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n723_), .A3(new_n719_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(G1338gat));
  NAND3_X1  g524(.A1(new_n704_), .A2(new_n212_), .A3(new_n538_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n647_), .A2(KEYINPUT111), .A3(new_n538_), .A4(new_n707_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(G106gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n647_), .A2(new_n538_), .A3(new_n707_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n727_), .B1(new_n729_), .B2(new_n732_), .ZN(new_n733_));
  AND4_X1   g532(.A1(new_n727_), .A2(new_n732_), .A3(G106gat), .A4(new_n728_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n726_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT53), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n737_), .B(new_n726_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1339gat));
  NAND2_X1  g538(.A1(new_n235_), .A2(new_n240_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n562_), .A2(new_n563_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n566_), .A2(new_n567_), .A3(new_n564_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n572_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n572_), .B2(new_n569_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT115), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n232_), .B1(new_n231_), .B2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n228_), .A2(KEYINPUT113), .A3(new_n230_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n231_), .A2(new_n232_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n747_), .A2(new_n748_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n233_), .A2(KEYINPUT114), .A3(KEYINPUT55), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT114), .B1(new_n233_), .B2(KEYINPUT55), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n751_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(KEYINPUT56), .A3(new_n242_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT56), .B1(new_n754_), .B2(new_n242_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n740_), .B(new_n745_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT58), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT118), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n277_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n745_), .A2(new_n740_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n754_), .A2(new_n242_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n762_), .B1(new_n765_), .B2(new_n755_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(KEYINPUT58), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n760_), .A2(new_n761_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n758_), .A2(KEYINPUT117), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n766_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(new_n772_), .A3(new_n759_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n740_), .A2(new_n575_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n765_), .B2(new_n755_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n745_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n244_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n274_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n769_), .A2(new_n773_), .B1(KEYINPUT57), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n778_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n617_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n300_), .A2(new_n576_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT112), .B1(new_n785_), .B2(KEYINPUT54), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(KEYINPUT54), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n300_), .A2(new_n788_), .A3(new_n789_), .A4(new_n576_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n786_), .A2(new_n787_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n784_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n489_), .A2(new_n665_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n793_), .A2(new_n463_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(KEYINPUT59), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n792_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n782_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n778_), .A2(KEYINPUT116), .A3(new_n781_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n780_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n779_), .A2(KEYINPUT57), .ZN(new_n804_));
  INV_X1    g603(.A(new_n773_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n760_), .A2(new_n768_), .A3(new_n761_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n799_), .A2(new_n800_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT119), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n297_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n803_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n795_), .B1(new_n811_), .B2(new_n791_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n575_), .B(new_n797_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(G113gat), .ZN(new_n815_));
  INV_X1    g614(.A(G113gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n816_), .A3(new_n575_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1340gat));
  OAI211_X1 g617(.A(new_n248_), .B(new_n797_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G120gat), .ZN(new_n820_));
  INV_X1    g619(.A(G120gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n674_), .B2(KEYINPUT60), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n812_), .B(new_n822_), .C1(KEYINPUT60), .C2(new_n821_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(G1341gat));
  AOI21_X1  g623(.A(G127gat), .B1(new_n812_), .B2(new_n298_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n811_), .A2(new_n791_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n794_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n827_), .A2(KEYINPUT59), .B1(new_n792_), .B2(new_n796_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT120), .B(G127gat), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n810_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n825_), .B1(new_n828_), .B2(new_n830_), .ZN(G1342gat));
  OAI211_X1 g630(.A(new_n761_), .B(new_n797_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(G134gat), .ZN(new_n833_));
  INV_X1    g632(.A(G134gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n812_), .A2(new_n834_), .A3(new_n586_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1343gat));
  XNOR2_X1  g635(.A(KEYINPUT121), .B(G141gat), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n606_), .A2(new_n538_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n838_), .A2(new_n488_), .A3(new_n593_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n826_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n837_), .B1(new_n840_), .B2(new_n575_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n826_), .A2(new_n839_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n837_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n842_), .A2(new_n576_), .A3(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n841_), .A2(new_n844_), .ZN(G1344gat));
  NAND3_X1  g644(.A1(new_n840_), .A2(new_n333_), .A3(new_n248_), .ZN(new_n846_));
  OAI21_X1  g645(.A(G148gat), .B1(new_n842_), .B2(new_n674_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1345gat));
  XNOR2_X1  g647(.A(KEYINPUT61), .B(G155gat), .ZN(new_n849_));
  OR3_X1    g648(.A1(new_n842_), .A2(new_n617_), .A3(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n842_), .B2(new_n617_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1346gat));
  AOI21_X1  g651(.A(G162gat), .B1(new_n840_), .B2(new_n586_), .ZN(new_n853_));
  INV_X1    g652(.A(G162gat), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n842_), .A2(new_n854_), .A3(new_n626_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1347gat));
  NAND2_X1  g655(.A1(new_n488_), .A2(new_n593_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n606_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT122), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n538_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n784_), .B2(new_n791_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT22), .B(G169gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n575_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n575_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(KEYINPUT62), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n428_), .B1(new_n866_), .B2(KEYINPUT62), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n864_), .B1(new_n869_), .B2(new_n870_), .ZN(G1348gat));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n773_), .A2(new_n761_), .A3(new_n768_), .A4(new_n760_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n873_), .A2(new_n804_), .A3(new_n799_), .A4(new_n800_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n297_), .B1(new_n874_), .B2(KEYINPUT119), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n787_), .A2(new_n790_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n875_), .A2(new_n803_), .B1(new_n786_), .B2(new_n876_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n674_), .A2(new_n859_), .A3(new_n429_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n877_), .A2(new_n538_), .A3(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(G176gat), .B1(new_n862_), .B2(new_n248_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n872_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n792_), .A2(new_n248_), .A3(new_n860_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n429_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n826_), .A2(new_n402_), .A3(new_n878_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(KEYINPUT124), .A3(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n886_), .ZN(G1349gat));
  INV_X1    g686(.A(new_n862_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n888_), .A2(new_n422_), .A3(new_n810_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n859_), .A2(new_n617_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n826_), .A2(new_n402_), .A3(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(G183gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n889_), .B1(new_n891_), .B2(new_n892_), .ZN(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n888_), .B2(new_n277_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n862_), .A2(new_n423_), .A3(new_n586_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1351gat));
  NOR2_X1   g695(.A1(new_n838_), .A2(new_n857_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n826_), .A2(new_n897_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n898_), .A2(new_n375_), .A3(new_n576_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n897_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n877_), .A2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G197gat), .B1(new_n901_), .B2(new_n575_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n899_), .A2(new_n902_), .ZN(G1352gat));
  OAI211_X1 g702(.A(KEYINPUT125), .B(G204gat), .C1(new_n898_), .C2(new_n674_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n901_), .A2(new_n248_), .A3(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1353gat));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n908_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n909_));
  AOI211_X1 g708(.A(new_n909_), .B(new_n810_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n901_), .A2(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n908_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n913_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n901_), .A2(new_n912_), .A3(new_n910_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1354gat));
  NAND2_X1  g715(.A1(new_n901_), .A2(new_n586_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT127), .B(G218gat), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n277_), .A2(new_n918_), .ZN(new_n919_));
  AOI22_X1  g718(.A1(new_n917_), .A2(new_n918_), .B1(new_n901_), .B2(new_n919_), .ZN(G1355gat));
endmodule


