//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G43gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G183gat), .ZN(new_n206_));
  OR2_X1    g005(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n207_));
  NAND2_X1  g006(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT84), .ZN(new_n210_));
  INV_X1    g009(.A(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT26), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n212_), .B(KEYINPUT85), .Z(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(KEYINPUT84), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215_));
  AOI22_X1  g014(.A1(KEYINPUT25), .A2(new_n206_), .B1(new_n215_), .B2(G190gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n210_), .A2(new_n213_), .A3(new_n214_), .A4(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT86), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT86), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT24), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n224_), .B1(G169gat), .B2(G176gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT87), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT87), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n223_), .A2(new_n228_), .A3(new_n225_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT23), .B1(new_n206_), .B2(new_n211_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(G183gat), .A3(G190gat), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(new_n224_), .B2(new_n222_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n217_), .A2(new_n227_), .A3(new_n229_), .A4(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(G169gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n232_), .A2(new_n238_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n237_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n235_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT89), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT89), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n235_), .A2(new_n246_), .A3(new_n243_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G227gat), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(G15gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n245_), .A2(new_n247_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n251_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT90), .B(KEYINPUT30), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n253_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n256_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n205_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n253_), .A2(new_n255_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n256_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n205_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(new_n257_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n260_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT91), .ZN(new_n267_));
  XOR2_X1   g066(.A(G127gat), .B(G134gat), .Z(new_n268_));
  XOR2_X1   g067(.A(G113gat), .B(G120gat), .Z(new_n269_));
  AOI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n268_), .B(new_n269_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n271_), .B2(new_n267_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT31), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT92), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n266_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT92), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n260_), .A2(new_n276_), .A3(new_n273_), .A4(new_n265_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  NOR3_X1   g080(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT93), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT2), .ZN(new_n285_));
  INV_X1    g084(.A(G141gat), .ZN(new_n286_));
  INV_X1    g085(.A(G148gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n288_), .B(new_n289_), .C1(new_n290_), .C2(new_n291_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n280_), .B(new_n281_), .C1(new_n284_), .C2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT94), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT29), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n279_), .B1(KEYINPUT1), .B2(new_n281_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n281_), .A2(KEYINPUT1), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n286_), .A2(new_n287_), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n299_), .A2(new_n291_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n295_), .A2(new_n296_), .A3(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G22gat), .B(G50gat), .Z(new_n306_));
  OR2_X1    g105(.A1(new_n293_), .A2(new_n294_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n293_), .A2(new_n294_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n301_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n304_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n296_), .A3(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n305_), .A2(new_n306_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n306_), .B1(new_n305_), .B2(new_n311_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G211gat), .B(G218gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(KEYINPUT98), .B(G204gat), .Z(new_n318_));
  INV_X1    g117(.A(G197gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(KEYINPUT97), .B(G197gat), .Z(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(G204gat), .B2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n317_), .B1(new_n322_), .B2(KEYINPUT21), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(G204gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(new_n319_), .B2(new_n318_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n323_), .B1(KEYINPUT21), .B2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(KEYINPUT21), .A3(new_n317_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n309_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(G233gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT96), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n333_), .A2(G228gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(G228gat), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n332_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n331_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n337_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n339_), .B(new_n328_), .C1(new_n309_), .C2(new_n296_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G78gat), .B(G106gat), .Z(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT100), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT101), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n315_), .A2(KEYINPUT102), .A3(new_n342_), .A4(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n338_), .A2(new_n340_), .A3(new_n345_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n306_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n303_), .A2(new_n304_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n310_), .B1(new_n309_), .B2(new_n296_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(KEYINPUT102), .A3(new_n312_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n345_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n347_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n346_), .A2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n344_), .B(new_n341_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n295_), .A2(new_n302_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n272_), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n271_), .B(KEYINPUT103), .Z(new_n360_));
  NAND2_X1  g159(.A1(new_n309_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(KEYINPUT4), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT104), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n359_), .A2(KEYINPUT104), .A3(new_n361_), .A4(KEYINPUT4), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n358_), .A2(new_n367_), .A3(new_n272_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n366_), .A2(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n359_), .A2(new_n361_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n369_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G85gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT0), .B(G57gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  NAND3_X1  g178(.A1(new_n373_), .A2(new_n375_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n371_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n375_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n381_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G8gat), .B(G36gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT18), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G64gat), .B(G92gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n326_), .A2(new_n327_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT19), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n237_), .B1(new_n233_), .B2(new_n242_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n222_), .A2(new_n224_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT25), .B(G183gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n215_), .A2(G190gat), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n212_), .A3(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n226_), .A2(new_n396_), .A3(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n395_), .B1(new_n241_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT20), .B1(new_n328_), .B2(new_n401_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n392_), .A2(new_n394_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n394_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n245_), .A2(new_n391_), .A3(new_n247_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n406_), .B1(new_n328_), .B2(new_n401_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n390_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n407_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n394_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n254_), .A2(new_n328_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n402_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n404_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(new_n414_), .A3(new_n389_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n409_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT27), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n394_), .B1(new_n392_), .B2(new_n402_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n419_), .B1(new_n394_), .B2(new_n410_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n390_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(KEYINPUT27), .A3(new_n415_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  NOR4_X1   g222(.A1(new_n278_), .A2(new_n357_), .A3(new_n385_), .A4(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n385_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n357_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n368_), .A2(new_n369_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n428_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n359_), .A2(new_n370_), .A3(new_n361_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n381_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT105), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n428_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n366_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT105), .ZN(new_n435_));
  INV_X1    g234(.A(new_n431_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n382_), .A2(new_n383_), .A3(new_n381_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n432_), .A2(new_n437_), .B1(new_n438_), .B2(KEYINPUT33), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n416_), .B1(new_n380_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n389_), .A2(KEYINPUT32), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n411_), .A2(new_n414_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT106), .ZN(new_n444_));
  INV_X1    g243(.A(new_n442_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n420_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT106), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n411_), .A2(new_n414_), .A3(new_n447_), .A4(new_n442_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n444_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n439_), .A2(new_n441_), .B1(new_n385_), .B2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n427_), .B1(new_n450_), .B2(new_n357_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n424_), .B1(new_n451_), .B2(new_n278_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G190gat), .B(G218gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G134gat), .B(G162gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n455_), .B(KEYINPUT36), .Z(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(G85gat), .ZN(new_n458_));
  INV_X1    g257(.A(G92gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT8), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT6), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G99gat), .A3(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT64), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n466_), .A2(new_n468_), .A3(KEYINPUT64), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G99gat), .A2(G106gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT7), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT66), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n476_), .A2(KEYINPUT66), .A3(new_n477_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n475_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n464_), .B1(new_n473_), .B2(new_n482_), .ZN(new_n483_));
  NOR4_X1   g282(.A1(new_n479_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT66), .B1(new_n476_), .B2(new_n477_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n469_), .B(new_n474_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n463_), .B1(new_n486_), .B2(new_n462_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n466_), .A2(new_n468_), .A3(KEYINPUT64), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT64), .B1(new_n466_), .B2(new_n468_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n492_));
  INV_X1    g291(.A(G106gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n460_), .A2(KEYINPUT9), .A3(new_n461_), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n461_), .A2(KEYINPUT9), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT65), .B1(new_n491_), .B2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT65), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n473_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n488_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G29gat), .B(G36gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT35), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G232gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n504_), .A2(new_n507_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n499_), .B(new_n502_), .C1(new_n483_), .C2(new_n487_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n507_), .B(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT74), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n514_), .A2(KEYINPUT74), .A3(new_n516_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n513_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n512_), .A2(new_n508_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n522_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n513_), .A2(new_n524_), .A3(new_n519_), .A4(new_n520_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n457_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n455_), .A2(KEYINPUT36), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n523_), .A2(new_n527_), .A3(new_n525_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT75), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n523_), .A2(KEYINPUT75), .A3(new_n527_), .A4(new_n525_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n526_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT108), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AOI211_X1 g333(.A(KEYINPUT108), .B(new_n526_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n452_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G1gat), .B(G8gat), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n539_), .A2(KEYINPUT77), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(KEYINPUT77), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G15gat), .B(G22gat), .ZN(new_n543_));
  INV_X1    g342(.A(G8gat), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n540_), .A2(new_n545_), .A3(new_n543_), .A4(new_n541_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n550_), .B(KEYINPUT78), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n549_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT67), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT11), .ZN(new_n556_));
  INV_X1    g355(.A(G57gat), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n557_), .A2(G64gat), .ZN(new_n558_));
  INV_X1    g357(.A(G64gat), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(G57gat), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n556_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(G71gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(G78gat), .ZN(new_n563_));
  INV_X1    g362(.A(G78gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(G71gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n555_), .B1(new_n561_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n559_), .A2(G57gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n557_), .A2(G64gat), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT11), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G71gat), .B(G78gat), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n570_), .A2(KEYINPUT67), .A3(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n554_), .B1(new_n567_), .B2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT67), .B1(new_n570_), .B2(new_n571_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n566_), .B(new_n555_), .C1(new_n553_), .C2(KEYINPUT11), .ZN(new_n575_));
  INV_X1    g374(.A(new_n554_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT69), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n573_), .A2(KEYINPUT69), .A3(new_n577_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n552_), .B(new_n582_), .Z(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n584_));
  XOR2_X1   g383(.A(G127gat), .B(G155gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n583_), .A2(new_n584_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n578_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n552_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n552_), .A2(new_n591_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n589_), .B(KEYINPUT17), .Z(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n590_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n504_), .A2(KEYINPUT68), .A3(new_n591_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n514_), .A2(new_n578_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT68), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(new_n514_), .B2(new_n578_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n504_), .B2(new_n591_), .ZN(new_n605_));
  XOR2_X1   g404(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n606_));
  NAND2_X1  g405(.A1(new_n599_), .A2(new_n606_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n576_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n608_), .A2(new_n609_), .A3(new_n579_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT69), .B1(new_n573_), .B2(new_n577_), .ZN(new_n611_));
  OAI211_X1 g410(.A(KEYINPUT12), .B(new_n514_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n605_), .A2(new_n607_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n604_), .A2(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(G120gat), .B(G148gat), .Z(new_n615_));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n604_), .A2(new_n613_), .A3(new_n619_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT13), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n621_), .A2(KEYINPUT13), .A3(new_n622_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n516_), .A2(new_n549_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n547_), .A2(new_n548_), .A3(new_n507_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(G229gat), .A2(G233gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n629_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n507_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n630_), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G113gat), .B(G141gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G169gat), .B(G197gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n637_), .B(new_n638_), .Z(new_n639_));
  NAND3_X1  g438(.A1(new_n633_), .A2(new_n636_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT81), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT82), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n642_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n633_), .A2(new_n636_), .ZN(new_n646_));
  OAI22_X1  g445(.A1(new_n644_), .A2(new_n645_), .B1(new_n646_), .B2(new_n639_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n645_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n646_), .A2(new_n639_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n643_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n628_), .A2(new_n651_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n538_), .A2(new_n597_), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n202_), .B1(new_n653_), .B2(new_n385_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT37), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n530_), .A2(new_n531_), .ZN(new_n656_));
  OAI211_X1 g455(.A(KEYINPUT76), .B(new_n655_), .C1(new_n656_), .C2(new_n526_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT76), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT37), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(KEYINPUT37), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n532_), .A2(new_n659_), .A3(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n657_), .A2(new_n627_), .A3(new_n597_), .A4(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n452_), .A2(new_n651_), .A3(new_n663_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n385_), .A2(KEYINPUT107), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n385_), .A2(KEYINPUT107), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(new_n202_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT38), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n654_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n672_), .B1(new_n670_), .B2(new_n669_), .ZN(G1324gat));
  NAND3_X1  g472(.A1(new_n664_), .A2(new_n544_), .A3(new_n423_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT39), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n653_), .A2(new_n423_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(G8gat), .ZN(new_n677_));
  AOI211_X1 g476(.A(KEYINPUT39), .B(new_n544_), .C1(new_n653_), .C2(new_n423_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT40), .B(new_n674_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1325gat));
  INV_X1    g482(.A(new_n278_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n250_), .B1(new_n653_), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT41), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n664_), .A2(new_n250_), .A3(new_n684_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1326gat));
  INV_X1    g487(.A(G22gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n653_), .B2(new_n357_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n664_), .A2(new_n689_), .A3(new_n357_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1327gat));
  NOR2_X1   g493(.A1(new_n357_), .A2(new_n423_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n684_), .A2(new_n695_), .A3(new_n426_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n355_), .A2(new_n356_), .A3(new_n380_), .A4(new_n384_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n423_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n449_), .A2(new_n385_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n437_), .A2(new_n432_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n438_), .A2(KEYINPUT33), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n415_), .B(new_n409_), .C1(new_n438_), .C2(KEYINPUT33), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n355_), .A2(new_n356_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n698_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n696_), .B1(new_n706_), .B2(new_n684_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n651_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n536_), .A2(new_n597_), .ZN(new_n709_));
  AND4_X1   g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n627_), .A4(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G29gat), .B1(new_n710_), .B2(new_n385_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n657_), .A2(new_n662_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(KEYINPUT43), .B1(new_n452_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n707_), .A2(new_n715_), .A3(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n652_), .A2(new_n596_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT44), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n452_), .A2(KEYINPUT43), .A3(new_n713_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n715_), .B1(new_n707_), .B2(new_n712_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT44), .B(new_n719_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT110), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n718_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(new_n726_), .A3(KEYINPUT44), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n720_), .B1(new_n724_), .B2(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n668_), .A2(G29gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n711_), .B1(new_n728_), .B2(new_n729_), .ZN(G1328gat));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731_));
  INV_X1    g530(.A(G36gat), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n724_), .A2(new_n727_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n423_), .B1(new_n725_), .B2(KEYINPUT44), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n732_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n710_), .A2(new_n732_), .A3(new_n423_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT45), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n731_), .B1(new_n736_), .B2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n734_), .B1(new_n724_), .B2(new_n727_), .ZN(new_n741_));
  OAI211_X1 g540(.A(KEYINPUT46), .B(new_n738_), .C1(new_n741_), .C2(new_n732_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1329gat));
  NOR2_X1   g542(.A1(new_n278_), .A2(new_n204_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n745_), .B(new_n720_), .C1(new_n724_), .C2(new_n727_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G43gat), .B1(new_n710_), .B2(new_n684_), .ZN(new_n747_));
  OAI21_X1  g546(.A(KEYINPUT47), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n728_), .A2(new_n744_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750_));
  INV_X1    g549(.A(new_n747_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n748_), .A2(new_n752_), .ZN(G1330gat));
  AOI21_X1  g552(.A(G50gat), .B1(new_n710_), .B2(new_n357_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n357_), .A2(G50gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n728_), .B2(new_n755_), .ZN(G1331gat));
  NOR3_X1   g555(.A1(new_n627_), .A2(new_n708_), .A3(new_n596_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n538_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G57gat), .B1(new_n759_), .B2(new_n426_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n452_), .A2(new_n708_), .A3(new_n627_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n761_), .A2(new_n597_), .A3(new_n713_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n557_), .A3(new_n668_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n760_), .A2(new_n763_), .ZN(G1332gat));
  AOI21_X1  g563(.A(new_n559_), .B1(new_n758_), .B2(new_n423_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT48), .Z(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(new_n559_), .A3(new_n423_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1333gat));
  AOI21_X1  g567(.A(new_n562_), .B1(new_n758_), .B2(new_n684_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT49), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n762_), .A2(new_n562_), .A3(new_n684_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1334gat));
  AOI21_X1  g571(.A(new_n564_), .B1(new_n758_), .B2(new_n357_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT50), .Z(new_n774_));
  NAND3_X1  g573(.A1(new_n762_), .A2(new_n564_), .A3(new_n357_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1335gat));
  NOR3_X1   g575(.A1(new_n627_), .A2(new_n708_), .A3(new_n597_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n717_), .A2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT111), .ZN(new_n779_));
  OAI21_X1  g578(.A(G85gat), .B1(new_n779_), .B2(new_n426_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n761_), .A2(new_n709_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n458_), .A3(new_n668_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1336gat));
  OAI21_X1  g582(.A(G92gat), .B1(new_n779_), .B2(new_n425_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(new_n459_), .A3(new_n423_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(G1337gat));
  OAI21_X1  g585(.A(G99gat), .B1(new_n778_), .B2(new_n278_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n781_), .A2(new_n684_), .A3(new_n492_), .A4(new_n494_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n787_), .A2(new_n788_), .B1(KEYINPUT112), .B2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(KEYINPUT112), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n790_), .B(new_n791_), .ZN(G1338gat));
  NAND3_X1  g591(.A1(new_n781_), .A2(new_n493_), .A3(new_n357_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n717_), .A2(new_n357_), .A3(new_n777_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n794_), .A2(new_n795_), .A3(G106gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n794_), .B2(G106gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n793_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT53), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n800_), .B(new_n793_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1339gat));
  OR3_X1    g601(.A1(new_n663_), .A2(KEYINPUT54), .A3(new_n708_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT54), .B1(new_n663_), .B2(new_n708_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n647_), .A2(new_n650_), .A3(new_n622_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n605_), .A2(new_n607_), .A3(new_n612_), .A4(KEYINPUT55), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT12), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n491_), .A2(KEYINPUT65), .A3(new_n498_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n501_), .B1(new_n473_), .B2(new_n500_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n464_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n474_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n491_), .B2(new_n815_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n486_), .A2(new_n462_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n463_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n810_), .B1(new_n813_), .B2(new_n818_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n582_), .A2(new_n819_), .B1(new_n599_), .B2(new_n606_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n820_), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(new_n605_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n809_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n613_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT113), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n613_), .A2(new_n826_), .A3(new_n823_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n820_), .A2(new_n601_), .A3(new_n598_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n603_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n822_), .A2(new_n825_), .A3(new_n827_), .A4(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n620_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n620_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n806_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n630_), .A2(new_n635_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n639_), .B1(new_n836_), .B2(new_n632_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n629_), .A2(new_n631_), .A3(new_n634_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n646_), .A2(new_n639_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n623_), .A2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n536_), .B1(new_n835_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(KEYINPUT115), .A3(new_n842_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n536_), .B(KEYINPUT57), .C1(new_n835_), .C2(new_n840_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n622_), .A2(new_n839_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT116), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n620_), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT56), .B1(new_n830_), .B2(new_n620_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n849_), .B(KEYINPUT58), .C1(new_n850_), .C2(new_n851_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n712_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .A4(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n805_), .B1(new_n857_), .B2(new_n596_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n684_), .A2(new_n695_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n667_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n858_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(G113gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n708_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT59), .B1(new_n858_), .B2(new_n861_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT117), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n867_), .B(KEYINPUT59), .C1(new_n858_), .C2(new_n861_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n843_), .A2(new_n847_), .A3(new_n856_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT118), .B1(new_n870_), .B2(new_n596_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n805_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n870_), .A2(KEYINPUT118), .A3(new_n596_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(new_n876_), .A3(new_n860_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n869_), .A2(new_n708_), .A3(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n864_), .B1(new_n878_), .B2(new_n863_), .ZN(G1340gat));
  INV_X1    g678(.A(G120gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n627_), .B2(KEYINPUT60), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n862_), .B(new_n881_), .C1(KEYINPUT60), .C2(new_n880_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n873_), .A2(new_n871_), .A3(new_n805_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n860_), .A2(new_n876_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n628_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G120gat), .B1(new_n886_), .B2(KEYINPUT119), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888_));
  AOI211_X1 g687(.A(new_n888_), .B(new_n885_), .C1(new_n866_), .C2(new_n868_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n882_), .B1(new_n887_), .B2(new_n889_), .ZN(G1341gat));
  NOR3_X1   g689(.A1(new_n858_), .A2(new_n596_), .A3(new_n861_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892_));
  OR3_X1    g691(.A1(new_n891_), .A2(new_n892_), .A3(G127gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n891_), .B2(G127gat), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n869_), .A2(new_n877_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n597_), .A2(G127gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(G1342gat));
  INV_X1    g697(.A(G134gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n862_), .A2(new_n899_), .A3(new_n537_), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n869_), .A2(new_n712_), .A3(new_n877_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(G1343gat));
  NOR2_X1   g701(.A1(new_n858_), .A2(new_n684_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n667_), .A2(new_n705_), .A3(new_n423_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n651_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT121), .B(G141gat), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1344gat));
  NOR2_X1   g707(.A1(new_n905_), .A2(new_n627_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(new_n287_), .ZN(G1345gat));
  OAI21_X1  g709(.A(KEYINPUT122), .B1(new_n905_), .B2(new_n596_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n903_), .A2(new_n912_), .A3(new_n597_), .A4(new_n904_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT61), .B(G155gat), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n911_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n911_), .B2(new_n913_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1346gat));
  OAI21_X1  g716(.A(G162gat), .B1(new_n905_), .B2(new_n713_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n536_), .A2(G162gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n905_), .B2(new_n919_), .ZN(G1347gat));
  NAND3_X1  g719(.A1(new_n667_), .A2(new_n684_), .A3(new_n423_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n357_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n875_), .A2(new_n708_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(KEYINPUT124), .B1(new_n923_), .B2(G169gat), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n925_));
  INV_X1    g724(.A(new_n923_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(KEYINPUT22), .B(G169gat), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n924_), .A2(new_n925_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  OR2_X1    g727(.A1(new_n924_), .A2(new_n925_), .ZN(new_n929_));
  AND3_X1   g728(.A1(new_n923_), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n928_), .B1(new_n929_), .B2(new_n930_), .ZN(G1348gat));
  INV_X1    g730(.A(G176gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n875_), .A2(new_n922_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(new_n627_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n858_), .A2(new_n357_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n921_), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n935_), .A2(G176gat), .A3(new_n628_), .A4(new_n936_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n934_), .A2(new_n937_), .ZN(G1349gat));
  NOR3_X1   g737(.A1(new_n933_), .A2(new_n397_), .A3(new_n596_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n935_), .A2(new_n597_), .A3(new_n936_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n939_), .B1(new_n206_), .B2(new_n940_), .ZN(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n933_), .B2(new_n713_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n537_), .A2(new_n212_), .A3(new_n398_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n933_), .B2(new_n943_), .ZN(G1351gat));
  NOR2_X1   g743(.A1(new_n425_), .A2(new_n697_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n903_), .A2(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n946_), .A2(new_n651_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(new_n319_), .ZN(G1352gat));
  INV_X1    g747(.A(G204gat), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(KEYINPUT125), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n318_), .B1(new_n951_), .B2(new_n949_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n946_), .A2(new_n627_), .ZN(new_n953_));
  MUX2_X1   g752(.A(new_n950_), .B(new_n952_), .S(new_n953_), .Z(G1353gat));
  NAND2_X1  g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n597_), .A2(new_n955_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(KEYINPUT126), .ZN(new_n957_));
  OAI21_X1  g756(.A(KEYINPUT127), .B1(new_n946_), .B2(new_n957_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960_));
  INV_X1    g759(.A(new_n957_), .ZN(new_n961_));
  NAND4_X1  g760(.A1(new_n903_), .A2(new_n960_), .A3(new_n945_), .A4(new_n961_), .ZN(new_n962_));
  AND3_X1   g761(.A1(new_n958_), .A2(new_n959_), .A3(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n959_), .B1(new_n958_), .B2(new_n962_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n963_), .A2(new_n964_), .ZN(G1354gat));
  OAI21_X1  g764(.A(G218gat), .B1(new_n946_), .B2(new_n713_), .ZN(new_n966_));
  OR2_X1    g765(.A1(new_n536_), .A2(G218gat), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n966_), .B1(new_n946_), .B2(new_n967_), .ZN(G1355gat));
endmodule


