//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n927_, new_n928_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n952_, new_n953_,
    new_n954_, new_n956_, new_n957_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n967_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G1gat), .A2(G8gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT14), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G29gat), .B(G36gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n212_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT73), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT73), .B1(new_n213_), .B2(new_n214_), .ZN(new_n218_));
  NOR3_X1   g017(.A1(new_n210_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n213_), .A2(new_n214_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT73), .ZN(new_n221_));
  INV_X1    g020(.A(new_n218_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n209_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n203_), .B1(new_n219_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(KEYINPUT15), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n215_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n227_), .A3(new_n209_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n210_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT74), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .A4(new_n202_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n224_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n229_), .A3(new_n202_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT74), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G113gat), .B(G141gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT75), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G169gat), .B(G197gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n232_), .A2(KEYINPUT76), .A3(new_n234_), .A4(new_n238_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n234_), .A2(new_n224_), .A3(new_n231_), .A4(new_n238_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT76), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n232_), .A2(new_n234_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n238_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n239_), .A2(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT24), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n246_), .B1(G169gat), .B2(G176gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT78), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(G169gat), .B2(G176gat), .ZN(new_n249_));
  INV_X1    g048(.A(G169gat), .ZN(new_n250_));
  INV_X1    g049(.A(G176gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(KEYINPUT78), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n247_), .A2(new_n249_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT24), .B1(new_n252_), .B2(new_n249_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n256_));
  INV_X1    g055(.A(G183gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT77), .B(G183gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(new_n256_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G190gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT23), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(G183gat), .A3(G190gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT79), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT79), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n266_), .A2(new_n263_), .A3(G183gat), .A4(G190gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(G190gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT23), .B1(new_n257_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n255_), .A2(new_n262_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n264_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n259_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n273_), .B1(new_n274_), .B2(G190gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(G169gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n272_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G227gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G15gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n279_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT31), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G71gat), .B(G99gat), .ZN(new_n285_));
  INV_X1    g084(.A(G43gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G127gat), .B(G134gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G113gat), .B(G120gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n289_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n284_), .B(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT81), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT2), .ZN(new_n301_));
  NAND3_X1  g100(.A1(KEYINPUT81), .A2(G141gat), .A3(G148gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n307_));
  INV_X1    g106(.A(G141gat), .ZN(new_n308_));
  INV_X1    g107(.A(G148gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT84), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT84), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n312_), .A2(new_n307_), .A3(new_n308_), .A4(new_n309_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n303_), .A2(new_n306_), .A3(new_n311_), .A4(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT82), .ZN(new_n315_));
  INV_X1    g114(.A(G155gat), .ZN(new_n316_));
  INV_X1    g115(.A(G162gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n314_), .A2(new_n321_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n300_), .A2(new_n302_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n308_), .A2(new_n309_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT83), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(new_n320_), .B2(KEYINPUT1), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n327_), .A2(KEYINPUT83), .A3(G155gat), .A4(G162gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n320_), .A2(KEYINPUT1), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n318_), .A2(new_n330_), .A3(new_n319_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n323_), .B(new_n324_), .C1(new_n329_), .C2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n322_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n293_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n322_), .A2(new_n292_), .A3(new_n332_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(KEYINPUT4), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n292_), .B1(new_n322_), .B2(new_n332_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n337_), .A2(KEYINPUT98), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT98), .B1(new_n337_), .B2(new_n338_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n297_), .B(new_n336_), .C1(new_n339_), .C2(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n334_), .A2(new_n335_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n296_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(G85gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT0), .B(G57gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n346_), .B(new_n347_), .Z(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n344_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n341_), .A2(new_n343_), .A3(new_n348_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT29), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n322_), .A2(new_n353_), .A3(new_n332_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT85), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n322_), .A2(KEYINPUT85), .A3(new_n332_), .A4(new_n353_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n358_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G22gat), .B(G50gat), .Z(new_n361_));
  NOR3_X1   g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n361_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n358_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n329_), .A2(new_n331_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n323_), .A2(new_n324_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n365_), .A2(new_n366_), .B1(new_n314_), .B2(new_n321_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT85), .B1(new_n367_), .B2(new_n353_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n357_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n364_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n363_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G78gat), .B(G106gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G218gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(G211gat), .ZN(new_n376_));
  INV_X1    g175(.A(G211gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G218gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n379_), .A2(KEYINPUT21), .ZN(new_n380_));
  INV_X1    g179(.A(G197gat), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT87), .B1(new_n381_), .B2(G204gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT87), .ZN(new_n383_));
  INV_X1    g182(.A(G204gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n384_), .A3(G197gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n381_), .A2(G204gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n382_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n380_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n384_), .A2(G197gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n386_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n379_), .B1(KEYINPUT21), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT89), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n393_), .A2(new_n382_), .A3(new_n386_), .A4(new_n385_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n391_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n392_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n388_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G228gat), .A2(G233gat), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n398_), .B(new_n399_), .C1(new_n353_), .C2(new_n367_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n381_), .A2(G204gat), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n384_), .A2(G197gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT21), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n379_), .ZN(new_n404_));
  XOR2_X1   g203(.A(KEYINPUT88), .B(KEYINPUT21), .Z(new_n405_));
  OAI211_X1 g204(.A(new_n403_), .B(new_n404_), .C1(new_n387_), .C2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT89), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n407_), .A2(new_n395_), .B1(new_n387_), .B2(new_n380_), .ZN(new_n408_));
  XOR2_X1   g207(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n409_));
  AOI21_X1  g208(.A(new_n409_), .B1(new_n322_), .B2(new_n332_), .ZN(new_n410_));
  OAI211_X1 g209(.A(G228gat), .B(G233gat), .C1(new_n408_), .C2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n374_), .B1(new_n400_), .B2(new_n411_), .ZN(new_n412_));
  OAI22_X1  g211(.A1(new_n362_), .A2(new_n372_), .B1(new_n412_), .B2(KEYINPUT91), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n400_), .A2(new_n411_), .A3(new_n374_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n361_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n370_), .A2(new_n363_), .A3(new_n371_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n420_), .A2(KEYINPUT91), .A3(new_n415_), .A4(new_n414_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n352_), .B1(new_n417_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT27), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(KEYINPUT93), .B(KEYINPUT20), .C1(new_n398_), .C2(new_n279_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n250_), .A2(KEYINPUT22), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT22), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G169gat), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n429_), .A2(new_n431_), .A3(KEYINPUT96), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT96), .B1(new_n429_), .B2(new_n431_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n251_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n263_), .B1(G183gat), .B2(G190gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(G183gat), .A2(G190gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT97), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT97), .ZN(new_n441_));
  INV_X1    g240(.A(new_n439_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n271_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n436_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n445_), .B1(new_n270_), .B2(new_n264_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT95), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n435_), .A2(KEYINPUT24), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n449_), .A2(KEYINPUT94), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(KEYINPUT94), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n450_), .A2(new_n249_), .A3(new_n252_), .A4(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT25), .B(G183gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n261_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n448_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n398_), .B1(new_n444_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n428_), .A2(new_n457_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n438_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n459_), .A2(new_n262_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n408_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT93), .B1(new_n461_), .B2(KEYINPUT20), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n427_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G8gat), .B(G36gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT18), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G64gat), .B(G92gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n398_), .B2(new_n279_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n443_), .A2(new_n440_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n436_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n446_), .B(KEYINPUT95), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n454_), .A3(new_n452_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n408_), .A3(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n469_), .A2(new_n475_), .A3(new_n426_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n463_), .A2(new_n467_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n467_), .B1(new_n463_), .B2(new_n476_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n423_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n463_), .A2(new_n467_), .A3(new_n476_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n426_), .B1(new_n469_), .B2(new_n475_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n458_), .A2(new_n462_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n481_), .B1(new_n482_), .B2(new_n426_), .ZN(new_n483_));
  OAI211_X1 g282(.A(KEYINPUT27), .B(new_n480_), .C1(new_n483_), .C2(new_n467_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n422_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n417_), .A2(new_n421_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n351_), .A2(KEYINPUT33), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT33), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n341_), .A2(new_n488_), .A3(new_n343_), .A4(new_n348_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n467_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n468_), .B1(new_n408_), .B2(new_n460_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n472_), .A2(new_n474_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n492_), .A2(KEYINPUT93), .B1(new_n493_), .B2(new_n398_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n461_), .A2(KEYINPUT20), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT93), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n426_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n476_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n491_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n348_), .B1(new_n342_), .B2(new_n297_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n336_), .A2(new_n296_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n339_), .A2(new_n340_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n490_), .A2(new_n500_), .A3(new_n480_), .A4(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n467_), .A2(KEYINPUT32), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT99), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n463_), .A2(new_n476_), .A3(new_n507_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n352_), .B(new_n508_), .C1(new_n483_), .C2(new_n506_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n486_), .B1(new_n505_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n295_), .B1(new_n485_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n479_), .A2(new_n484_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n512_), .A2(new_n486_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n295_), .A2(new_n352_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n245_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n517_));
  INV_X1    g316(.A(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT64), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT64), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(G106gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n517_), .A2(new_n519_), .A3(new_n521_), .A4(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT6), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(G99gat), .A3(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n529_), .A2(KEYINPUT9), .ZN(new_n530_));
  INV_X1    g329(.A(G85gat), .ZN(new_n531_));
  INV_X1    g330(.A(G92gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(KEYINPUT9), .A3(new_n529_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n523_), .A2(new_n528_), .A3(new_n530_), .A4(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n533_), .A2(KEYINPUT65), .A3(new_n529_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n525_), .A2(new_n527_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT7), .ZN(new_n539_));
  INV_X1    g338(.A(G99gat), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n518_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n537_), .B1(new_n538_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT8), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n528_), .A2(new_n542_), .A3(new_n541_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT8), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n537_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n536_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n215_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT70), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G232gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT34), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(KEYINPUT35), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n225_), .A2(new_n227_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n533_), .A2(KEYINPUT65), .A3(new_n529_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n541_), .A2(new_n542_), .ZN(new_n557_));
  AOI211_X1 g356(.A(KEYINPUT8), .B(new_n556_), .C1(new_n557_), .C2(new_n528_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n547_), .B1(new_n546_), .B2(new_n537_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n535_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n554_), .B1(new_n555_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n551_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n553_), .A2(KEYINPUT35), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n563_), .B(KEYINPUT69), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n551_), .A2(new_n566_), .A3(new_n561_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G190gat), .B(G218gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G134gat), .B(G162gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT36), .Z(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n571_), .A2(KEYINPUT36), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n565_), .A2(new_n574_), .A3(new_n567_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(KEYINPUT71), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT37), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n573_), .A2(KEYINPUT71), .A3(KEYINPUT37), .A4(new_n575_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT12), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n560_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(G71gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(G78gat), .ZN(new_n584_));
  INV_X1    g383(.A(G78gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(G71gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G57gat), .B(G64gat), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n587_), .B1(new_n588_), .B2(KEYINPUT11), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT66), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n588_), .B2(KEYINPUT11), .ZN(new_n591_));
  INV_X1    g390(.A(G64gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(G57gat), .ZN(new_n593_));
  INV_X1    g392(.A(G57gat), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(G64gat), .ZN(new_n595_));
  AND4_X1   g394(.A1(new_n590_), .A2(new_n593_), .A3(new_n595_), .A4(KEYINPUT11), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n589_), .B1(new_n591_), .B2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n593_), .A2(new_n595_), .A3(KEYINPUT11), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT66), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n593_), .A2(new_n595_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT11), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n593_), .A2(new_n595_), .A3(new_n590_), .A4(KEYINPUT11), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n599_), .A2(new_n602_), .A3(new_n587_), .A4(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n597_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n560_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n597_), .A2(new_n604_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n545_), .A2(new_n548_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n608_), .B2(new_n535_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n582_), .B1(new_n606_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n581_), .B1(new_n549_), .B2(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT67), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n560_), .A2(new_n605_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT67), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(new_n581_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n610_), .A2(new_n612_), .A3(new_n613_), .A4(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n608_), .A2(new_n535_), .A3(new_n607_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n613_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(G120gat), .B(G148gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G176gat), .B(G204gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n622_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n627_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n617_), .A2(new_n621_), .A3(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n631_), .A2(KEYINPUT13), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(KEYINPUT13), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n210_), .B(new_n607_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT72), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G127gat), .B(G155gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT16), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G183gat), .B(G211gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT17), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n638_), .B(new_n643_), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n637_), .A2(KEYINPUT17), .A3(new_n642_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n580_), .A2(new_n634_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n516_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n352_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n649_), .A2(G1gat), .A3(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT38), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n511_), .A2(new_n515_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n573_), .A2(new_n575_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n655_), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT100), .B(new_n657_), .C1(new_n511_), .C2(new_n515_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n634_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n239_), .A2(new_n242_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n243_), .A2(new_n244_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(new_n647_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n659_), .A2(new_n352_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n652_), .B1(G1gat), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT101), .ZN(G1324gat));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n659_), .A2(new_n665_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n512_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G8gat), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT39), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n649_), .A2(G8gat), .A3(new_n671_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT102), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n677_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n669_), .B1(new_n675_), .B2(new_n678_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n672_), .A2(new_n673_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n680_), .A2(KEYINPUT40), .A3(new_n674_), .A4(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1325gat));
  OAI21_X1  g481(.A(G15gat), .B1(new_n670_), .B2(new_n295_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT41), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n649_), .A2(G15gat), .A3(new_n295_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1326gat));
  INV_X1    g485(.A(new_n486_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G22gat), .B1(new_n670_), .B2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n687_), .A2(G22gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n649_), .B2(new_n691_), .ZN(G1327gat));
  NOR2_X1   g491(.A1(new_n646_), .A2(new_n655_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n516_), .A2(new_n660_), .A3(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n352_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n664_), .A2(new_n646_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n654_), .A2(new_n580_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(KEYINPUT43), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n578_), .A2(new_n579_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n704_), .B2(KEYINPUT104), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n698_), .B1(new_n701_), .B2(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(KEYINPUT44), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT43), .B1(new_n699_), .B2(new_n700_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n704_), .A2(KEYINPUT104), .A3(new_n702_), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT44), .B(new_n697_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n706_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n707_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n352_), .A2(G29gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n696_), .B1(new_n714_), .B2(new_n715_), .ZN(G1328gat));
  NOR3_X1   g515(.A1(new_n694_), .A2(G36gat), .A3(new_n671_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT45), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n512_), .B1(new_n706_), .B2(KEYINPUT44), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n721_));
  INV_X1    g520(.A(G36gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n719_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OAI211_X1 g524(.A(KEYINPUT46), .B(new_n719_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1329gat));
  NAND2_X1  g526(.A1(new_n712_), .A2(new_n713_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n707_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n295_), .A2(new_n286_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n728_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n295_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G43gat), .B1(new_n695_), .B2(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT47), .B1(new_n731_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n714_), .A2(new_n730_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736_));
  INV_X1    g535(.A(new_n733_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n735_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n734_), .A2(new_n738_), .ZN(G1330gat));
  AND2_X1   g538(.A1(new_n486_), .A2(G50gat), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n728_), .A2(new_n729_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G50gat), .B1(new_n695_), .B2(new_n486_), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT106), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n714_), .A2(new_n740_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n745_));
  INV_X1    g544(.A(new_n742_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n744_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n743_), .A2(new_n747_), .ZN(G1331gat));
  NOR2_X1   g547(.A1(new_n660_), .A2(new_n663_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n654_), .A2(new_n749_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n750_), .A2(new_n646_), .A3(new_n703_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(new_n594_), .A3(new_n352_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n660_), .A2(new_n647_), .A3(new_n663_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n753_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT107), .B(new_n753_), .C1(new_n656_), .C2(new_n658_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n352_), .A3(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n752_), .B1(new_n758_), .B2(new_n594_), .ZN(G1332gat));
  NAND2_X1  g558(.A1(new_n512_), .A2(new_n592_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT109), .Z(new_n761_));
  NAND2_X1  g560(.A1(new_n751_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n756_), .A2(new_n512_), .A3(new_n757_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(G64gat), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G64gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(G1333gat));
  NAND3_X1  g566(.A1(new_n751_), .A2(new_n583_), .A3(new_n732_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n756_), .A2(new_n732_), .A3(new_n757_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G71gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G71gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(G1334gat));
  NAND3_X1  g572(.A1(new_n751_), .A2(new_n585_), .A3(new_n486_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n756_), .A2(new_n486_), .A3(new_n757_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(G78gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n775_), .B2(G78gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(KEYINPUT110), .B(new_n774_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1335gat));
  NAND2_X1  g582(.A1(new_n750_), .A2(new_n693_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n531_), .B1(new_n784_), .B2(new_n650_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n749_), .A2(new_n647_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n701_), .B2(new_n705_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n352_), .A2(G85gat), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT111), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n785_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT112), .ZN(G1336gat));
  OAI21_X1  g591(.A(G92gat), .B1(new_n788_), .B2(new_n671_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n512_), .A2(new_n532_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n784_), .B2(new_n794_), .ZN(G1337gat));
  AOI21_X1  g594(.A(new_n540_), .B1(new_n787_), .B2(new_n732_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n517_), .A2(new_n522_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n784_), .A2(new_n295_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799_));
  OAI22_X1  g598(.A1(new_n796_), .A2(new_n798_), .B1(new_n799_), .B2(KEYINPUT51), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(KEYINPUT51), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(G1338gat));
  NAND3_X1  g601(.A1(new_n486_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n784_), .A2(new_n803_), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n804_), .B(KEYINPUT114), .Z(new_n805_));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807_));
  OAI21_X1  g606(.A(G106gat), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n787_), .B2(new_n486_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n806_), .A2(new_n807_), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n810_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n805_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT53), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n805_), .A2(new_n811_), .A3(new_n815_), .A4(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1339gat));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n648_), .A2(new_n818_), .A3(new_n245_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n648_), .B2(new_n245_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n663_), .B2(new_n630_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n630_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n245_), .A2(KEYINPUT116), .A3(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n617_), .A2(KEYINPUT55), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n619_), .A2(new_n582_), .B1(new_n611_), .B2(KEYINPUT67), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n613_), .A4(new_n616_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n610_), .A2(new_n616_), .A3(new_n612_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n620_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n833_), .A2(new_n832_), .A3(new_n620_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n629_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT56), .B1(new_n836_), .B2(new_n627_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(KEYINPUT118), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n833_), .A2(new_n620_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT117), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n833_), .A2(new_n832_), .A3(new_n620_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n843_), .A2(new_n844_), .B1(new_n827_), .B2(new_n830_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT118), .B(new_n837_), .C1(new_n845_), .C2(new_n629_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n826_), .B1(new_n841_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n202_), .B1(new_n219_), .B2(new_n223_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n228_), .A2(new_n229_), .A3(new_n203_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n244_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n661_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT119), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n661_), .A2(new_n854_), .A3(new_n851_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n631_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n848_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n655_), .A2(KEYINPUT57), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n837_), .B1(new_n845_), .B2(new_n629_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n863_));
  INV_X1    g662(.A(new_n838_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n845_), .B2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n836_), .A2(KEYINPUT120), .A3(new_n838_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n862_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n824_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(new_n868_), .A3(KEYINPUT58), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n867_), .A2(new_n868_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n580_), .B(new_n869_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n843_), .A2(new_n844_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n629_), .B1(new_n874_), .B2(new_n831_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(new_n875_), .B2(KEYINPUT56), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n846_), .A3(new_n839_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n856_), .B1(new_n877_), .B2(new_n826_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n657_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n861_), .B(new_n872_), .C1(new_n879_), .C2(KEYINPUT57), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n821_), .B1(new_n880_), .B2(new_n647_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n295_), .A2(new_n650_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n513_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(G113gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n663_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT59), .B1(new_n881_), .B2(new_n883_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n871_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n869_), .A2(new_n580_), .ZN(new_n889_));
  OAI22_X1  g688(.A1(new_n888_), .A2(new_n889_), .B1(new_n878_), .B2(new_n859_), .ZN(new_n890_));
  AOI21_X1  g689(.A(KEYINPUT57), .B1(new_n858_), .B2(new_n655_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n647_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT122), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n880_), .A2(new_n894_), .A3(new_n647_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n821_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n883_), .A2(KEYINPUT59), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n887_), .B(new_n663_), .C1(new_n896_), .C2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n886_), .B1(new_n899_), .B2(new_n885_), .ZN(G1340gat));
  INV_X1    g699(.A(new_n821_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n892_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n903_));
  AOI21_X1  g702(.A(G120gat), .B1(new_n634_), .B2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n903_), .B2(G120gat), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n902_), .A2(new_n513_), .A3(new_n882_), .A4(new_n905_), .ZN(new_n906_));
  XOR2_X1   g705(.A(new_n906_), .B(KEYINPUT123), .Z(new_n907_));
  OAI21_X1  g706(.A(new_n887_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n908_));
  OAI21_X1  g707(.A(G120gat), .B1(new_n908_), .B2(new_n660_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1341gat));
  INV_X1    g709(.A(G127gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n884_), .A2(new_n911_), .A3(new_n646_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n887_), .B(new_n646_), .C1(new_n896_), .C2(new_n897_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n914_), .B2(new_n911_), .ZN(G1342gat));
  INV_X1    g714(.A(G134gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n884_), .A2(new_n916_), .A3(new_n657_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n887_), .B(new_n580_), .C1(new_n896_), .C2(new_n897_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n917_), .B1(new_n919_), .B2(new_n916_), .ZN(G1343gat));
  NOR3_X1   g719(.A1(new_n732_), .A2(new_n687_), .A3(new_n650_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n902_), .A2(new_n671_), .A3(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n245_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(new_n308_), .ZN(G1344gat));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n660_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n309_), .ZN(G1345gat));
  NOR2_X1   g725(.A1(new_n922_), .A2(new_n647_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT61), .B(G155gat), .Z(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1346gat));
  OAI21_X1  g728(.A(G162gat), .B1(new_n922_), .B2(new_n703_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n657_), .A2(new_n317_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n922_), .B2(new_n931_), .ZN(G1347gat));
  XNOR2_X1  g731(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n514_), .A2(new_n512_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n486_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n896_), .A2(new_n245_), .A3(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n933_), .B1(new_n937_), .B2(new_n250_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n933_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n892_), .A2(KEYINPUT122), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n894_), .B1(new_n880_), .B2(new_n647_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n901_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n935_), .ZN(new_n943_));
  OAI211_X1 g742(.A(G169gat), .B(new_n939_), .C1(new_n943_), .C2(new_n245_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n896_), .A2(new_n936_), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n945_), .B(new_n663_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n938_), .A2(new_n944_), .A3(new_n946_), .ZN(G1348gat));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n634_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n881_), .A2(new_n486_), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n660_), .A2(new_n934_), .A3(new_n251_), .ZN(new_n950_));
  AOI22_X1  g749(.A1(new_n948_), .A2(new_n251_), .B1(new_n949_), .B2(new_n950_), .ZN(G1349gat));
  NOR2_X1   g750(.A1(new_n934_), .A2(new_n647_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n274_), .B1(new_n949_), .B2(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n647_), .A2(new_n453_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n953_), .B1(new_n945_), .B2(new_n954_), .ZN(G1350gat));
  OAI21_X1  g754(.A(G190gat), .B1(new_n943_), .B2(new_n703_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n945_), .A2(new_n261_), .A3(new_n657_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1351gat));
  NAND3_X1  g757(.A1(new_n512_), .A2(new_n422_), .A3(new_n295_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n881_), .A2(new_n959_), .ZN(new_n960_));
  OR2_X1    g759(.A1(new_n381_), .A2(KEYINPUT125), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n381_), .A2(KEYINPUT125), .ZN(new_n962_));
  AOI22_X1  g761(.A1(new_n960_), .A2(new_n663_), .B1(new_n961_), .B2(new_n962_), .ZN(new_n963_));
  INV_X1    g762(.A(new_n960_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n964_), .A2(new_n245_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n963_), .B1(new_n965_), .B2(new_n962_), .ZN(G1352gat));
  NAND2_X1  g765(.A1(new_n960_), .A2(new_n634_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g767(.A(KEYINPUT63), .B(G211gat), .C1(new_n960_), .C2(new_n646_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n964_), .A2(new_n647_), .ZN(new_n970_));
  XOR2_X1   g769(.A(KEYINPUT63), .B(G211gat), .Z(new_n971_));
  AOI21_X1  g770(.A(new_n969_), .B1(new_n970_), .B2(new_n971_), .ZN(G1354gat));
  NOR4_X1   g771(.A1(new_n881_), .A2(G218gat), .A3(new_n655_), .A4(new_n959_), .ZN(new_n973_));
  INV_X1    g772(.A(new_n973_), .ZN(new_n974_));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n975_));
  NOR3_X1   g774(.A1(new_n881_), .A2(new_n703_), .A3(new_n959_), .ZN(new_n976_));
  OAI211_X1 g775(.A(new_n974_), .B(new_n975_), .C1(new_n375_), .C2(new_n976_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(new_n976_), .A2(new_n375_), .ZN(new_n978_));
  OAI21_X1  g777(.A(KEYINPUT126), .B1(new_n978_), .B2(new_n973_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n977_), .A2(new_n979_), .ZN(G1355gat));
endmodule


