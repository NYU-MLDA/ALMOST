//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n203_));
  NAND4_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT84), .A4(G183gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT25), .B(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n206_), .A2(KEYINPUT84), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n203_), .A2(G183gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT85), .B1(new_n208_), .B2(KEYINPUT84), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n204_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT23), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT86), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  OR3_X1    g016(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT23), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT87), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n223_), .A2(KEYINPUT24), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n219_), .A2(new_n220_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(KEYINPUT24), .A3(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n212_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n220_), .B1(new_n219_), .B2(new_n224_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n226_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n218_), .A2(new_n215_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n231_), .B1(G183gat), .B2(G190gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n232_), .B2(KEYINPUT90), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(KEYINPUT90), .B2(new_n232_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT22), .B1(new_n221_), .B2(KEYINPUT88), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n222_), .B(new_n235_), .C1(new_n236_), .C2(KEYINPUT88), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT89), .ZN(new_n238_));
  OAI22_X1  g037(.A1(new_n228_), .A2(new_n229_), .B1(new_n234_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G99gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G43gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n239_), .B(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G113gat), .B(G120gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT91), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n245_), .A2(new_n246_), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  NAND2_X1  g049(.A1(G227gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(G15gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT30), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n250_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n244_), .B(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G211gat), .B(G218gat), .Z(new_n257_));
  INV_X1    g056(.A(KEYINPUT21), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G197gat), .B(G204gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n258_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n260_), .B1(new_n262_), .B2(new_n257_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G155gat), .B(G162gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT94), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G141gat), .ZN(new_n267_));
  INV_X1    g066(.A(G148gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n269_), .A2(KEYINPUT2), .B1(KEYINPUT93), .B2(KEYINPUT3), .ZN(new_n270_));
  OR4_X1    g069(.A1(KEYINPUT93), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n268_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(KEYINPUT93), .B2(KEYINPUT3), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT2), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n270_), .A2(new_n271_), .A3(new_n273_), .A4(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n266_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT95), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n280_), .B1(KEYINPUT1), .B2(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n282_), .B1(KEYINPUT1), .B2(new_n281_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n269_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(new_n272_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n279_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n263_), .B1(new_n286_), .B2(KEYINPUT29), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G228gat), .A2(G233gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n287_), .B1(KEYINPUT96), .B2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(KEYINPUT96), .Z(new_n290_));
  OAI21_X1  g089(.A(new_n289_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G78gat), .B(G106gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT97), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n286_), .A2(KEYINPUT29), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G22gat), .B(G50gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT28), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n295_), .B(new_n297_), .Z(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n291_), .B(new_n292_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n300_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n286_), .A2(new_n250_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(KEYINPUT4), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n249_), .A2(new_n247_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT99), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n279_), .A2(new_n285_), .A3(new_n310_), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n304_), .A2(KEYINPUT4), .A3(new_n311_), .ZN(new_n312_));
  OR3_X1    g111(.A1(new_n308_), .A2(new_n312_), .A3(KEYINPUT100), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT100), .B1(new_n308_), .B2(new_n312_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G1gat), .B(G29gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(G85gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT0), .B(G57gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  NAND3_X1  g117(.A1(new_n304_), .A2(new_n311_), .A3(new_n306_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n313_), .A2(new_n314_), .A3(new_n318_), .A4(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT33), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT101), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT19), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n263_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n239_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n219_), .B1(G183gat), .B2(G190gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT22), .B(G169gat), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n230_), .B1(new_n332_), .B2(new_n222_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n211_), .A2(new_n205_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n231_), .A2(new_n224_), .A3(new_n227_), .A4(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT20), .B1(new_n337_), .B2(new_n328_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n327_), .B1(new_n330_), .B2(new_n338_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n239_), .A2(new_n328_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT20), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n337_), .B2(new_n328_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(new_n326_), .A3(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G8gat), .B(G36gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT18), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n339_), .A2(new_n343_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT98), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n351_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT98), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(new_n349_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n318_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n304_), .A2(new_n311_), .A3(new_n307_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n305_), .A2(new_n306_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n356_), .B(new_n357_), .C1(new_n358_), .C2(new_n312_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n352_), .A2(new_n355_), .A3(new_n359_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n320_), .A2(new_n321_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n320_), .A2(KEYINPUT101), .A3(new_n321_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n324_), .A2(new_n360_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n313_), .A2(new_n314_), .A3(new_n319_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n356_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n320_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n339_), .A2(new_n343_), .B1(KEYINPUT32), .B2(new_n347_), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n367_), .B(KEYINPUT102), .Z(new_n368_));
  AOI21_X1  g167(.A(new_n328_), .B1(new_n337_), .B2(KEYINPUT104), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(KEYINPUT104), .B2(new_n337_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT103), .B(KEYINPUT20), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(KEYINPUT105), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n329_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT105), .B1(new_n370_), .B2(new_n371_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n326_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n340_), .A2(new_n327_), .A3(new_n342_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n347_), .A2(KEYINPUT32), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n366_), .B(new_n368_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n303_), .B1(new_n363_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n366_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT27), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n383_));
  OAI211_X1 g182(.A(KEYINPUT27), .B(new_n353_), .C1(new_n377_), .C2(new_n347_), .ZN(new_n384_));
  AND4_X1   g183(.A1(new_n381_), .A2(new_n303_), .A3(new_n383_), .A4(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n256_), .B1(new_n380_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n383_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n303_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n381_), .A2(new_n255_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n386_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT72), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT69), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G99gat), .A2(G106gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT66), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(KEYINPUT6), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n399_), .A2(KEYINPUT66), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n396_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(KEYINPUT66), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n397_), .A2(KEYINPUT6), .ZN(new_n403_));
  AND2_X1   g202(.A1(G99gat), .A2(G106gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT7), .ZN(new_n407_));
  INV_X1    g206(.A(G99gat), .ZN(new_n408_));
  INV_X1    g207(.A(G106gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n401_), .A2(new_n405_), .A3(new_n406_), .A4(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT8), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G85gat), .A2(G92gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G85gat), .A2(G92gat), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT68), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n411_), .A2(new_n412_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n412_), .B1(new_n411_), .B2(new_n416_), .ZN(new_n418_));
  OR2_X1    g217(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n409_), .A3(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n401_), .A2(new_n405_), .A3(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(new_n415_), .B2(KEYINPUT64), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT64), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n425_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n425_), .B1(G85gat), .B2(G92gat), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n427_), .B1(new_n432_), .B2(new_n423_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(KEYINPUT65), .A3(new_n426_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n422_), .B1(new_n431_), .B2(new_n434_), .ZN(new_n435_));
  OAI22_X1  g234(.A1(new_n417_), .A2(new_n418_), .B1(new_n435_), .B2(KEYINPUT67), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n401_), .A2(new_n405_), .A3(new_n421_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n429_), .A2(new_n430_), .ZN(new_n438_));
  AOI21_X1  g237(.A(KEYINPUT65), .B1(new_n433_), .B2(new_n426_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT67), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n395_), .B1(new_n436_), .B2(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n404_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n410_), .A2(new_n406_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n416_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT8), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n411_), .A2(new_n412_), .A3(new_n416_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n440_), .A2(new_n441_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n435_), .A2(KEYINPUT67), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(KEYINPUT69), .A4(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G57gat), .B(G64gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT11), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT70), .ZN(new_n457_));
  XOR2_X1   g256(.A(G71gat), .B(G78gat), .Z(new_n458_));
  OAI21_X1  g257(.A(new_n458_), .B1(KEYINPUT11), .B2(new_n455_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n459_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n443_), .A2(new_n454_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT71), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n436_), .B2(new_n442_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n451_), .A2(new_n452_), .A3(KEYINPUT71), .A4(new_n453_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT12), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n466_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n463_), .B1(new_n443_), .B2(new_n454_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n464_), .B(new_n470_), .C1(new_n471_), .C2(KEYINPUT12), .ZN(new_n472_));
  INV_X1    g271(.A(G230gat), .ZN(new_n473_));
  INV_X1    g272(.A(G233gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n394_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n449_), .A2(new_n450_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT69), .B1(new_n477_), .B2(new_n453_), .ZN(new_n478_));
  AND4_X1   g277(.A1(KEYINPUT69), .A2(new_n451_), .A3(new_n452_), .A4(new_n453_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n462_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n464_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n475_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n464_), .A2(new_n470_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n468_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n475_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(KEYINPUT72), .A4(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n476_), .A2(new_n482_), .A3(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G120gat), .B(G148gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT74), .ZN(new_n489_));
  XOR2_X1   g288(.A(G176gat), .B(G204gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  NAND2_X1  g292(.A1(new_n487_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n493_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n476_), .A2(new_n486_), .A3(new_n482_), .A4(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n494_), .A2(KEYINPUT13), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT13), .B1(new_n494_), .B2(new_n496_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(G1gat), .ZN(new_n501_));
  INV_X1    g300(.A(G8gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT14), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G15gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT78), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT78), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(G15gat), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n505_), .A2(new_n507_), .A3(G22gat), .ZN(new_n508_));
  AOI21_X1  g307(.A(G22gat), .B1(new_n505_), .B2(new_n507_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n503_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G1gat), .B(G8gat), .Z(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G29gat), .B(G36gat), .Z(new_n514_));
  XOR2_X1   g313(.A(G43gat), .B(G50gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n511_), .B(new_n503_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n516_), .B(KEYINPUT15), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n513_), .A2(new_n517_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT82), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT83), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n516_), .B1(new_n513_), .B2(new_n517_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(KEYINPUT81), .A3(new_n518_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT81), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n531_), .B1(new_n519_), .B2(new_n528_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n530_), .A2(new_n532_), .A3(G229gat), .A4(G233gat), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n522_), .A2(KEYINPUT83), .A3(new_n524_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n527_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G113gat), .B(G141gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G169gat), .B(G197gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(new_n537_), .Z(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n527_), .A2(new_n533_), .A3(new_n534_), .A4(new_n538_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n500_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n393_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n521_), .B(KEYINPUT79), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(new_n462_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G127gat), .B(G155gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT16), .ZN(new_n553_));
  XOR2_X1   g352(.A(G183gat), .B(G211gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n550_), .B1(new_n551_), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n551_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n549_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n466_), .A2(new_n520_), .A3(new_n467_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n443_), .A2(new_n516_), .A3(new_n454_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT34), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT35), .Z(new_n565_));
  NAND4_X1  g364(.A1(new_n561_), .A2(new_n562_), .A3(KEYINPUT76), .A4(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n561_), .A2(new_n562_), .A3(new_n565_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT76), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(KEYINPUT35), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n566_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G190gat), .B(G218gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(KEYINPUT75), .B(KEYINPUT36), .Z(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n572_), .A2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n575_), .B(KEYINPUT36), .Z(new_n579_));
  OAI211_X1 g378(.A(new_n566_), .B(new_n579_), .C1(new_n569_), .C2(new_n571_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT77), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n583_), .A3(KEYINPUT37), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT37), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n578_), .B(new_n580_), .C1(new_n582_), .C2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n560_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT80), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n545_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n501_), .A3(new_n366_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT38), .ZN(new_n592_));
  INV_X1    g391(.A(new_n581_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n560_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n545_), .A2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT106), .Z(new_n596_));
  AND2_X1   g395(.A1(new_n596_), .A2(new_n366_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n592_), .B1(new_n597_), .B2(new_n501_), .ZN(G1324gat));
  INV_X1    g397(.A(KEYINPUT40), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n545_), .A2(new_n387_), .A3(new_n594_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(KEYINPUT107), .A3(G8gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT39), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT107), .B1(new_n600_), .B2(G8gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n590_), .A2(new_n502_), .A3(new_n387_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n602_), .A2(new_n603_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n599_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n607_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n609_), .A2(KEYINPUT40), .A3(new_n604_), .A4(new_n605_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(G1325gat));
  NAND3_X1  g410(.A1(new_n590_), .A2(new_n504_), .A3(new_n255_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n596_), .A2(new_n255_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT41), .B1(new_n613_), .B2(G15gat), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT41), .ZN(new_n615_));
  AOI211_X1 g414(.A(new_n615_), .B(new_n504_), .C1(new_n596_), .C2(new_n255_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n612_), .B1(new_n614_), .B2(new_n616_), .ZN(G1326gat));
  INV_X1    g416(.A(G22gat), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n590_), .A2(new_n618_), .A3(new_n303_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT42), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n596_), .A2(new_n303_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n620_), .B1(new_n621_), .B2(G22gat), .ZN(new_n622_));
  AOI211_X1 g421(.A(KEYINPUT42), .B(new_n618_), .C1(new_n596_), .C2(new_n303_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n619_), .B1(new_n622_), .B2(new_n623_), .ZN(G1327gat));
  INV_X1    g423(.A(KEYINPUT43), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n584_), .A2(new_n586_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n625_), .B1(new_n393_), .B2(new_n627_), .ZN(new_n628_));
  AOI211_X1 g427(.A(KEYINPUT43), .B(new_n626_), .C1(new_n386_), .C2(new_n392_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n544_), .A2(new_n560_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT108), .Z(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(KEYINPUT44), .A3(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n632_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT44), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n366_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G29gat), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n559_), .A2(new_n581_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n545_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n381_), .A2(G29gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT109), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n639_), .B1(new_n641_), .B2(new_n643_), .ZN(G1328gat));
  NOR3_X1   g443(.A1(new_n641_), .A2(G36gat), .A3(new_n388_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT45), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n633_), .A2(new_n387_), .A3(new_n636_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G36gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT46), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n647_), .A2(new_n649_), .A3(KEYINPUT46), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1329gat));
  NAND4_X1  g453(.A1(new_n633_), .A2(G43gat), .A3(new_n255_), .A4(new_n636_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n641_), .A2(new_n256_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(G43gat), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g457(.A(G50gat), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n389_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n545_), .A2(new_n303_), .A3(new_n640_), .ZN(new_n661_));
  AOI22_X1  g460(.A1(new_n637_), .A2(new_n660_), .B1(new_n659_), .B2(new_n661_), .ZN(G1331gat));
  NOR2_X1   g461(.A1(new_n499_), .A2(new_n542_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n393_), .A2(new_n663_), .ZN(new_n664_));
  AND4_X1   g463(.A1(G57gat), .A2(new_n664_), .A3(new_n366_), .A4(new_n594_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n588_), .A2(new_n500_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n588_), .A2(KEYINPUT110), .A3(new_n500_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n393_), .A2(new_n668_), .A3(new_n543_), .A4(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT111), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n381_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n672_), .B1(new_n671_), .B2(new_n670_), .ZN(new_n673_));
  INV_X1    g472(.A(G57gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n665_), .B1(new_n673_), .B2(new_n674_), .ZN(G1332gat));
  OR3_X1    g474(.A1(new_n670_), .A2(G64gat), .A3(new_n388_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n664_), .A2(new_n387_), .A3(new_n594_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G64gat), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n678_), .A2(KEYINPUT113), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(KEYINPUT113), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n676_), .B1(new_n682_), .B2(new_n683_), .ZN(G1333gat));
  NAND3_X1  g483(.A1(new_n664_), .A2(new_n255_), .A3(new_n594_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G71gat), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT115), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n670_), .A2(G71gat), .A3(new_n256_), .ZN(new_n690_));
  OR3_X1    g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n689_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1334gat));
  NAND3_X1  g492(.A1(new_n664_), .A2(new_n303_), .A3(new_n594_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G78gat), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT116), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT116), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n694_), .A2(new_n697_), .A3(G78gat), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT50), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n696_), .A2(KEYINPUT50), .A3(new_n698_), .ZN(new_n702_));
  OR3_X1    g501(.A1(new_n670_), .A2(G78gat), .A3(new_n389_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n701_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT117), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT117), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n701_), .A2(new_n702_), .A3(new_n706_), .A4(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1335gat));
  NAND2_X1  g507(.A1(new_n663_), .A2(new_n560_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n630_), .A2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G85gat), .B1(new_n711_), .B2(new_n381_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n664_), .A2(new_n640_), .ZN(new_n713_));
  INV_X1    g512(.A(G85gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n366_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1336gat));
  OAI21_X1  g515(.A(G92gat), .B1(new_n711_), .B2(new_n388_), .ZN(new_n717_));
  INV_X1    g516(.A(G92gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n713_), .A2(new_n718_), .A3(new_n387_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1337gat));
  OAI21_X1  g519(.A(G99gat), .B1(new_n711_), .B2(new_n256_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n713_), .A2(new_n419_), .A3(new_n420_), .A4(new_n255_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g523(.A1(new_n713_), .A2(new_n409_), .A3(new_n303_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n303_), .B(new_n710_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(G106gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n726_), .B2(G106gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g530(.A(KEYINPUT121), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT120), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n530_), .A2(new_n532_), .A3(new_n524_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT119), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(new_n735_), .A3(new_n539_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n524_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n522_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n735_), .B1(new_n734_), .B2(new_n539_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n541_), .B(new_n733_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n541_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT120), .ZN(new_n743_));
  AOI221_X4 g542(.A(new_n732_), .B1(new_n741_), .B2(new_n743_), .C1(new_n494_), .C2(new_n496_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n494_), .A2(new_n496_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n741_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT121), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n744_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n472_), .A2(new_n749_), .A3(new_n475_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n485_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n476_), .A2(new_n749_), .A3(new_n486_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT56), .B1(new_n754_), .B2(new_n493_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  AOI211_X1 g555(.A(new_n756_), .B(new_n495_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n542_), .B(new_n496_), .C1(new_n755_), .C2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n593_), .B1(new_n748_), .B2(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n746_), .A2(new_n496_), .ZN(new_n760_));
  OAI211_X1 g559(.A(KEYINPUT58), .B(new_n760_), .C1(new_n755_), .C2(new_n757_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT58), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n626_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n759_), .A2(KEYINPUT57), .B1(new_n761_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT122), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n766_), .B1(new_n759_), .B2(KEYINPUT57), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n745_), .A2(new_n746_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n732_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n745_), .A2(KEYINPUT121), .A3(new_n746_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n496_), .A2(new_n542_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n754_), .A2(new_n493_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n756_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n754_), .A2(KEYINPUT56), .A3(new_n493_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n772_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n581_), .B1(new_n771_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(KEYINPUT122), .A3(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n765_), .A2(new_n767_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n560_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n497_), .A2(new_n498_), .A3(new_n542_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n587_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n782_), .A2(new_n587_), .A3(KEYINPUT118), .A4(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n782_), .A2(new_n587_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT54), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n786_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n781_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT123), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT123), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n781_), .A2(new_n794_), .A3(new_n791_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n390_), .A2(new_n381_), .A3(new_n256_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n793_), .A2(new_n542_), .A3(new_n795_), .A4(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(G113gat), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT124), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT124), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n797_), .A2(new_n801_), .A3(new_n798_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n796_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n765_), .B1(KEYINPUT57), .B2(new_n759_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n560_), .ZN(new_n805_));
  AOI211_X1 g604(.A(KEYINPUT59), .B(new_n803_), .C1(new_n805_), .C2(new_n791_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n543_), .A2(new_n798_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n794_), .B1(new_n781_), .B2(new_n791_), .ZN(new_n809_));
  AOI211_X1 g608(.A(KEYINPUT123), .B(new_n790_), .C1(new_n780_), .C2(new_n560_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n803_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT59), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n807_), .B(new_n808_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n800_), .A2(new_n802_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT125), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT125), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n800_), .A2(new_n816_), .A3(new_n813_), .A4(new_n802_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1340gat));
  NOR2_X1   g617(.A1(new_n499_), .A2(KEYINPUT60), .ZN(new_n819_));
  INV_X1    g618(.A(G120gat), .ZN(new_n820_));
  MUX2_X1   g619(.A(KEYINPUT60), .B(new_n819_), .S(new_n820_), .Z(new_n821_));
  NAND2_X1  g620(.A1(new_n811_), .A2(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT126), .ZN(new_n823_));
  INV_X1    g622(.A(new_n811_), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n499_), .B(new_n806_), .C1(new_n824_), .C2(KEYINPUT59), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n823_), .B1(new_n825_), .B2(new_n820_), .ZN(G1341gat));
  INV_X1    g625(.A(G127gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n811_), .A2(new_n827_), .A3(new_n559_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n560_), .B(new_n806_), .C1(new_n824_), .C2(KEYINPUT59), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n827_), .ZN(G1342gat));
  INV_X1    g629(.A(G134gat), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n811_), .A2(new_n831_), .A3(new_n593_), .ZN(new_n832_));
  AOI211_X1 g631(.A(new_n626_), .B(new_n806_), .C1(new_n824_), .C2(KEYINPUT59), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n831_), .ZN(G1343gat));
  NOR3_X1   g633(.A1(new_n809_), .A2(new_n810_), .A3(new_n255_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n389_), .A2(new_n387_), .A3(new_n381_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n543_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(new_n267_), .ZN(G1344gat));
  NOR2_X1   g638(.A1(new_n837_), .A2(new_n499_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(new_n268_), .ZN(G1345gat));
  NAND3_X1  g640(.A1(new_n835_), .A2(new_n559_), .A3(new_n836_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT61), .B(G155gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1346gat));
  OAI21_X1  g643(.A(G162gat), .B1(new_n837_), .B2(new_n626_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n581_), .A2(G162gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n837_), .B2(new_n846_), .ZN(G1347gat));
  AOI21_X1  g646(.A(new_n303_), .B1(new_n805_), .B2(new_n791_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n388_), .A2(new_n391_), .ZN(new_n849_));
  XOR2_X1   g648(.A(new_n849_), .B(KEYINPUT127), .Z(new_n850_));
  AND2_X1   g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n221_), .B1(new_n851_), .B2(new_n542_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n852_), .A2(KEYINPUT62), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(KEYINPUT62), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n542_), .A3(new_n332_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(G1348gat));
  AOI21_X1  g655(.A(G176gat), .B1(new_n851_), .B2(new_n500_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n809_), .A2(new_n810_), .A3(new_n303_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n850_), .A2(G176gat), .A3(new_n500_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(G1349gat));
  AND2_X1   g659(.A1(new_n850_), .A2(new_n559_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G183gat), .B1(new_n858_), .B2(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n861_), .A2(new_n206_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n848_), .B2(new_n863_), .ZN(G1350gat));
  NAND3_X1  g663(.A1(new_n851_), .A2(new_n211_), .A3(new_n593_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n851_), .A2(new_n627_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n214_), .ZN(G1351gat));
  NAND4_X1  g666(.A1(new_n835_), .A2(new_n381_), .A3(new_n303_), .A4(new_n387_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n543_), .ZN(new_n869_));
  INV_X1    g668(.A(G197gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1352gat));
  NOR2_X1   g670(.A1(new_n868_), .A2(new_n499_), .ZN(new_n872_));
  INV_X1    g671(.A(G204gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1353gat));
  XNOR2_X1  g673(.A(KEYINPUT63), .B(G211gat), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n868_), .A2(new_n560_), .A3(new_n875_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n868_), .A2(new_n560_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n877_), .B2(new_n878_), .ZN(G1354gat));
  OAI21_X1  g678(.A(G218gat), .B1(new_n868_), .B2(new_n626_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n581_), .A2(G218gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n868_), .B2(new_n881_), .ZN(G1355gat));
endmodule


