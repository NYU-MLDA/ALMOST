//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT4), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT2), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT84), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(new_n209_), .B2(KEYINPUT3), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(KEYINPUT84), .A3(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT85), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT83), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n215_), .A2(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(new_n218_), .B(KEYINPUT1), .Z(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n217_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(new_n208_), .A3(new_n205_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G127gat), .B(G134gat), .ZN(new_n224_));
  INV_X1    g023(.A(G113gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G120gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n220_), .A2(new_n223_), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n220_), .A2(KEYINPUT86), .A3(new_n223_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT86), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n215_), .A2(new_n219_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n223_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n228_), .B1(new_n230_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n229_), .B1(new_n235_), .B2(KEYINPUT94), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n229_), .A2(KEYINPUT94), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n204_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n235_), .A2(KEYINPUT4), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n203_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n236_), .A2(new_n202_), .A3(new_n237_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G57gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G85gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(G1gat), .B(G29gat), .Z(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n240_), .A2(new_n241_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT33), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT26), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G190gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT25), .B(G183gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT79), .B(G190gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n251_), .B(new_n252_), .C1(new_n254_), .C2(new_n250_), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n255_), .B(KEYINPUT80), .Z(new_n256_));
  NAND2_X1  g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT23), .ZN(new_n258_));
  INV_X1    g057(.A(G169gat), .ZN(new_n259_));
  INV_X1    g058(.A(G176gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n261_), .A2(KEYINPUT24), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G169gat), .A2(G176gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(KEYINPUT24), .A3(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n258_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n256_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT22), .B(G169gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n260_), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(KEYINPUT81), .Z(new_n270_));
  OAI21_X1  g069(.A(new_n258_), .B1(new_n254_), .B2(G183gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n263_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G197gat), .B(G204gat), .Z(new_n274_));
  AND2_X1   g073(.A1(new_n274_), .A2(KEYINPUT21), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G211gat), .B(G218gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n276_), .B1(new_n274_), .B2(KEYINPUT21), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n277_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT88), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n273_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT92), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G226gat), .A2(G233gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT19), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n258_), .B1(G183gat), .B2(G190gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(new_n263_), .A3(new_n269_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n250_), .A2(G190gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n252_), .A2(new_n251_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n289_), .B1(new_n292_), .B2(new_n265_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n280_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n287_), .A4(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n280_), .A2(new_n293_), .ZN(new_n296_));
  OAI211_X1 g095(.A(KEYINPUT20), .B(new_n296_), .C1(new_n273_), .C2(new_n282_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n286_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G8gat), .B(G36gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G64gat), .B(G92gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n295_), .A2(new_n298_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n303_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n236_), .A2(new_n237_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n245_), .B1(new_n308_), .B2(new_n202_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT95), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n202_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n312_));
  OAI211_X1 g111(.A(KEYINPUT95), .B(new_n245_), .C1(new_n308_), .C2(new_n202_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT33), .A4(new_n246_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n249_), .A2(new_n307_), .A3(new_n314_), .A4(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n297_), .A2(new_n286_), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n280_), .B(KEYINPUT90), .Z(new_n318_));
  OAI211_X1 g117(.A(new_n318_), .B(new_n289_), .C1(new_n292_), .C2(new_n265_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n317_), .B1(new_n320_), .B2(new_n286_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n303_), .A2(KEYINPUT32), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n295_), .A2(new_n298_), .A3(new_n322_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n247_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n246_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n323_), .B(new_n324_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n316_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(G228gat), .ZN(new_n329_));
  INV_X1    g128(.A(G233gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT89), .B(KEYINPUT29), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n220_), .B2(new_n223_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n318_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n335_), .B1(new_n230_), .B2(new_n234_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n282_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n334_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G78gat), .B(G106gat), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT91), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n230_), .A2(new_n234_), .A3(new_n335_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G22gat), .B(G50gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n344_), .B(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n334_), .B(new_n339_), .C1(new_n336_), .C2(new_n337_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n343_), .A2(new_n348_), .B1(new_n349_), .B2(new_n341_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n341_), .A2(new_n348_), .A3(KEYINPUT91), .A4(new_n349_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G71gat), .B(G99gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n228_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT30), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n267_), .A2(new_n359_), .A3(new_n272_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n267_), .B2(new_n272_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n358_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n362_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(new_n228_), .A3(new_n360_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G15gat), .B(G43gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G227gat), .A2(G233gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n363_), .A2(new_n365_), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n369_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n357_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n363_), .A2(new_n365_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n368_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n363_), .A2(new_n365_), .A3(new_n369_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n356_), .A3(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n328_), .A2(new_n353_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT27), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n380_));
  OAI211_X1 g179(.A(KEYINPUT27), .B(new_n304_), .C1(new_n321_), .C2(new_n303_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n326_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(KEYINPUT96), .A3(new_n247_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n377_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n343_), .A2(new_n348_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n341_), .A2(new_n349_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n372_), .A2(new_n376_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(new_n351_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT96), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n383_), .A2(new_n385_), .A3(new_n392_), .A4(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n378_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT13), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G57gat), .B(G64gat), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n398_), .A2(KEYINPUT11), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(KEYINPUT11), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G71gat), .B(G78gat), .ZN(new_n401_));
  OR3_X1    g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(new_n401_), .A3(KEYINPUT11), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT8), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G99gat), .A2(G106gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT7), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT6), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT65), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT65), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT6), .ZN(new_n412_));
  AND2_X1   g211(.A1(G99gat), .A2(G106gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G99gat), .A2(G106gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n411_), .A2(KEYINPUT6), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n409_), .A2(KEYINPUT65), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n408_), .A2(new_n414_), .A3(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G85gat), .B(G92gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n406_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n410_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n413_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT66), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT66), .B1(new_n418_), .B2(new_n414_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n408_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT8), .B1(new_n428_), .B2(KEYINPUT67), .ZN(new_n429_));
  INV_X1    g228(.A(new_n408_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n425_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n418_), .A2(KEYINPUT66), .A3(new_n414_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n430_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT67), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n420_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n422_), .B1(new_n429_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n431_), .A2(new_n432_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT64), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(G92gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n439_), .A2(KEYINPUT9), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n438_), .A2(G92gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(G85gat), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n421_), .A2(KEYINPUT9), .ZN(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT10), .B(G99gat), .Z(new_n444_));
  INV_X1    g243(.A(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n437_), .A2(new_n442_), .A3(new_n443_), .A4(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n405_), .B1(new_n436_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n422_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n421_), .B1(new_n428_), .B2(KEYINPUT67), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n406_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(new_n447_), .A3(new_n404_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n449_), .A2(KEYINPUT12), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT12), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n456_), .B(new_n405_), .C1(new_n436_), .C2(new_n448_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G230gat), .A2(G233gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n449_), .B2(new_n454_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G120gat), .B(G148gat), .Z(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G176gat), .B(G204gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n460_), .A2(new_n462_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n459_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n470_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n467_), .B1(new_n471_), .B2(new_n461_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n469_), .A2(KEYINPUT69), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT69), .B1(new_n469_), .B2(new_n472_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n397_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT69), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n468_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n471_), .A2(new_n461_), .A3(new_n467_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(KEYINPUT13), .A3(new_n473_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G113gat), .B(G141gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(new_n259_), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n485_), .B(G197gat), .Z(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G29gat), .B(G36gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(G43gat), .ZN(new_n489_));
  INV_X1    g288(.A(G50gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n488_), .A2(G43gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(G43gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(G50gat), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496_));
  INV_X1    g295(.A(G1gat), .ZN(new_n497_));
  INV_X1    g296(.A(G8gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G1gat), .B(G8gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n495_), .A2(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n503_), .A2(KEYINPUT78), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(KEYINPUT78), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n504_), .A2(new_n505_), .B1(new_n502_), .B2(new_n495_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G229gat), .A2(G233gat), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n505_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n491_), .A2(KEYINPUT15), .A3(new_n494_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT15), .B1(new_n491_), .B2(new_n494_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n502_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n510_), .A2(new_n515_), .A3(new_n507_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n487_), .B1(new_n509_), .B2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n516_), .B(new_n487_), .C1(new_n507_), .C2(new_n506_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n483_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n396_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT37), .ZN(new_n523_));
  INV_X1    g322(.A(new_n495_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n453_), .A2(new_n524_), .A3(new_n447_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT70), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n453_), .A2(KEYINPUT70), .A3(new_n524_), .A4(new_n447_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n513_), .B1(new_n453_), .B2(new_n447_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G232gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT34), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(KEYINPUT35), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n529_), .A2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(KEYINPUT35), .B(new_n532_), .C1(new_n530_), .C2(KEYINPUT71), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n529_), .A2(new_n536_), .A3(new_n534_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT72), .B(G190gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(G218gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G134gat), .B(G162gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n544_), .B(KEYINPUT36), .Z(new_n545_));
  AOI21_X1  g344(.A(new_n523_), .B1(new_n540_), .B2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n544_), .A2(KEYINPUT36), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n538_), .A2(new_n547_), .A3(new_n539_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT73), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n538_), .A2(KEYINPUT73), .A3(new_n547_), .A4(new_n539_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n546_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n529_), .A2(new_n536_), .A3(new_n534_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n536_), .B1(new_n534_), .B2(new_n529_), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT74), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT74), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n538_), .A2(new_n557_), .A3(new_n539_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n545_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT37), .B1(new_n559_), .B2(new_n548_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT16), .B(G183gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(G211gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G127gat), .B(G155gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT17), .Z(new_n565_));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT75), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n502_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(new_n405_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT77), .Z(new_n571_));
  INV_X1    g370(.A(new_n564_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n569_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n553_), .A2(new_n560_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n522_), .A2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n394_), .A2(new_n385_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n497_), .A3(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT38), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n559_), .A2(new_n548_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(new_n575_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n396_), .A2(new_n521_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT97), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n396_), .A2(new_n588_), .A3(new_n521_), .A4(new_n585_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(G1gat), .B1(new_n590_), .B2(new_n579_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n582_), .A2(new_n591_), .ZN(G1324gat));
  NAND3_X1  g391(.A1(new_n578_), .A2(new_n498_), .A3(new_n382_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT98), .Z(new_n594_));
  OAI21_X1  g393(.A(G8gat), .B1(new_n586_), .B2(new_n383_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT39), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT40), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n597_), .B(new_n599_), .ZN(G1325gat));
  INV_X1    g399(.A(G15gat), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n578_), .A2(new_n601_), .A3(new_n390_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT101), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n603_), .B(G15gat), .C1(new_n590_), .C2(new_n377_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n377_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT101), .B1(new_n605_), .B2(new_n601_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n604_), .A2(KEYINPUT41), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT41), .B1(new_n604_), .B2(new_n606_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n602_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(KEYINPUT102), .B(new_n602_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1326gat));
  OAI21_X1  g412(.A(G22gat), .B1(new_n590_), .B2(new_n353_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT42), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n353_), .A2(G22gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT103), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n578_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(G1327gat));
  INV_X1    g418(.A(new_n575_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n522_), .A2(new_n620_), .A3(new_n583_), .ZN(new_n621_));
  AOI21_X1  g420(.A(G29gat), .B1(new_n621_), .B2(new_n580_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n553_), .A2(new_n560_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n396_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n396_), .B2(new_n624_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n626_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n631_), .A2(new_n521_), .A3(new_n575_), .A4(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n392_), .A2(new_n385_), .A3(new_n394_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n353_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n316_), .B2(new_n327_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n383_), .A2(new_n635_), .B1(new_n637_), .B2(new_n377_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n628_), .B1(new_n638_), .B2(new_n623_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n396_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n639_), .A2(new_n640_), .A3(new_n521_), .A4(new_n575_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n632_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n634_), .A2(new_n580_), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n622_), .B1(new_n643_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g443(.A1(new_n634_), .A2(new_n382_), .A3(new_n642_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT106), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n634_), .A2(new_n642_), .A3(new_n647_), .A4(new_n382_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(G36gat), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(G36gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n621_), .A2(new_n650_), .A3(new_n382_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT45), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n649_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(KEYINPUT46), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n649_), .B(new_n652_), .C1(new_n654_), .C2(KEYINPUT46), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1329gat));
  NAND3_X1  g457(.A1(new_n634_), .A2(new_n390_), .A3(new_n642_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n377_), .A2(G43gat), .ZN(new_n660_));
  AOI22_X1  g459(.A1(new_n659_), .A2(G43gat), .B1(new_n621_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g461(.A(G50gat), .B1(new_n621_), .B2(new_n636_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n634_), .A2(new_n636_), .A3(new_n642_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(G50gat), .ZN(G1331gat));
  INV_X1    g464(.A(new_n520_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n482_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n638_), .A2(new_n577_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G57gat), .B1(new_n669_), .B2(new_n580_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n638_), .A2(new_n668_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(new_n585_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n580_), .A2(G57gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n670_), .B1(new_n672_), .B2(new_n673_), .ZN(G1332gat));
  INV_X1    g473(.A(G64gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n672_), .B2(new_n382_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT48), .Z(new_n677_));
  NAND2_X1  g476(.A1(new_n382_), .A2(new_n675_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT108), .Z(new_n679_));
  NAND2_X1  g478(.A1(new_n669_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n677_), .A2(new_n680_), .ZN(G1333gat));
  INV_X1    g480(.A(G71gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n672_), .B2(new_n390_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT49), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n669_), .A2(new_n682_), .A3(new_n390_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1334gat));
  INV_X1    g485(.A(G78gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n672_), .B2(new_n636_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT109), .Z(new_n689_));
  INV_X1    g488(.A(KEYINPUT50), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n690_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n669_), .A2(new_n687_), .A3(new_n636_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(G1335gat));
  NOR2_X1   g493(.A1(new_n583_), .A2(new_n620_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n671_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n671_), .A2(KEYINPUT110), .A3(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(G85gat), .B1(new_n700_), .B2(new_n580_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n639_), .A2(new_n640_), .A3(new_n575_), .A4(new_n667_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n580_), .A2(G85gat), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT111), .Z(new_n705_));
  AOI21_X1  g504(.A(new_n701_), .B1(new_n703_), .B2(new_n705_), .ZN(G1336gat));
  AOI21_X1  g505(.A(G92gat), .B1(new_n700_), .B2(new_n382_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n441_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n383_), .B1(new_n708_), .B2(new_n439_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n703_), .B2(new_n709_), .ZN(G1337gat));
  NAND3_X1  g509(.A1(new_n700_), .A2(new_n444_), .A3(new_n390_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G99gat), .B1(new_n702_), .B2(new_n377_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n713_), .B(new_n714_), .Z(G1338gat));
  OAI21_X1  g514(.A(G106gat), .B1(new_n702_), .B2(new_n353_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT52), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n718_), .B(G106gat), .C1(new_n702_), .C2(new_n353_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n636_), .A2(new_n445_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n720_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT113), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT113), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n720_), .A2(new_n726_), .A3(new_n723_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n725_), .A2(KEYINPUT53), .A3(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT53), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n726_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT113), .B(new_n722_), .C1(new_n717_), .C2(new_n719_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n729_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n728_), .A2(new_n732_), .ZN(G1339gat));
  NAND2_X1  g532(.A1(new_n583_), .A2(new_n523_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n734_), .A2(new_n520_), .A3(new_n620_), .A4(new_n552_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT54), .B1(new_n735_), .B2(new_n483_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT54), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n576_), .A2(new_n737_), .A3(new_n520_), .A4(new_n482_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n520_), .A2(new_n479_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n455_), .A2(new_n470_), .A3(new_n457_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT55), .B(new_n470_), .C1(new_n455_), .C2(new_n457_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n741_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n745_), .A2(KEYINPUT56), .A3(new_n467_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT56), .B1(new_n745_), .B2(new_n467_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n740_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n507_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n510_), .A2(new_n515_), .A3(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n750_), .B(new_n486_), .C1(new_n749_), .C2(new_n506_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n518_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n518_), .A2(new_n751_), .A3(KEYINPUT114), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n480_), .A2(new_n473_), .A3(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n480_), .A2(new_n756_), .A3(KEYINPUT115), .A4(new_n473_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n748_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n583_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT57), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n761_), .A2(KEYINPUT57), .A3(new_n583_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n746_), .A2(new_n747_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n766_), .A2(KEYINPUT58), .A3(new_n469_), .A4(new_n756_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n469_), .B(new_n756_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT58), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n624_), .A3(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n764_), .A2(new_n765_), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n739_), .B1(new_n575_), .B2(new_n772_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n579_), .A2(new_n382_), .A3(new_n391_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(G113gat), .B1(new_n776_), .B2(new_n666_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT116), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT59), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n761_), .A2(KEYINPUT57), .A3(new_n583_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT57), .B1(new_n761_), .B2(new_n583_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n620_), .B1(new_n783_), .B2(new_n771_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT59), .B(new_n774_), .C1(new_n784_), .C2(new_n739_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n780_), .A2(new_n785_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n786_), .A2(new_n225_), .A3(new_n520_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n778_), .A2(new_n787_), .ZN(G1340gat));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n780_), .A2(new_n785_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n483_), .ZN(new_n792_));
  AOI211_X1 g591(.A(KEYINPUT118), .B(new_n482_), .C1(new_n780_), .C2(new_n785_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n227_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n227_), .B1(new_n482_), .B2(KEYINPUT60), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n227_), .A2(KEYINPUT60), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n776_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n776_), .A2(KEYINPUT117), .A3(new_n795_), .A4(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n789_), .B1(new_n794_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n792_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n791_), .A2(new_n790_), .A3(new_n483_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(G120gat), .A3(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n801_), .A3(KEYINPUT119), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n803_), .A2(new_n807_), .ZN(G1341gat));
  AOI21_X1  g607(.A(G127gat), .B1(new_n776_), .B2(new_n620_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n620_), .A2(G127gat), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT120), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n809_), .B1(new_n791_), .B2(new_n811_), .ZN(G1342gat));
  AOI21_X1  g611(.A(G134gat), .B1(new_n776_), .B2(new_n584_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n786_), .A2(new_n623_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g614(.A1(new_n773_), .A2(new_n386_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n579_), .A2(new_n382_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT121), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(KEYINPUT121), .A3(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n666_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n483_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT122), .B(G148gat), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n825_), .B(new_n826_), .ZN(G1345gat));
  NAND2_X1  g626(.A1(new_n822_), .A2(new_n620_), .ZN(new_n828_));
  XOR2_X1   g627(.A(KEYINPUT61), .B(G155gat), .Z(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT123), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n828_), .B(new_n830_), .Z(G1346gat));
  AOI21_X1  g630(.A(G162gat), .B1(new_n822_), .B2(new_n584_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n623_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(G162gat), .B2(new_n833_), .ZN(G1347gat));
  NOR2_X1   g633(.A1(new_n580_), .A2(new_n383_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n390_), .ZN(new_n836_));
  XOR2_X1   g635(.A(new_n836_), .B(KEYINPUT124), .Z(new_n837_));
  NOR2_X1   g636(.A1(new_n773_), .A2(new_n636_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n259_), .B1(new_n840_), .B2(new_n666_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n841_), .A2(KEYINPUT62), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n840_), .A2(new_n666_), .A3(new_n268_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(KEYINPUT62), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n842_), .A2(new_n843_), .A3(new_n844_), .ZN(G1348gat));
  NOR2_X1   g644(.A1(new_n839_), .A2(new_n482_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(new_n260_), .ZN(G1349gat));
  INV_X1    g646(.A(KEYINPUT125), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n839_), .A2(new_n575_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n252_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n849_), .A2(G183gat), .ZN(new_n852_));
  NOR4_X1   g651(.A1(new_n839_), .A2(KEYINPUT125), .A3(new_n252_), .A4(new_n575_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n851_), .A2(new_n852_), .A3(new_n853_), .ZN(G1350gat));
  OAI21_X1  g653(.A(G190gat), .B1(new_n839_), .B2(new_n623_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n584_), .A2(new_n251_), .A3(new_n290_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n839_), .B2(new_n856_), .ZN(G1351gat));
  AND2_X1   g656(.A1(new_n816_), .A2(new_n835_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n666_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT126), .B(G197gat), .Z(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1352gat));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n483_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g662(.A1(new_n858_), .A2(new_n620_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n865_));
  AND2_X1   g664(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n864_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n864_), .B2(new_n865_), .ZN(G1354gat));
  AOI21_X1  g667(.A(G218gat), .B1(new_n858_), .B2(new_n584_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n624_), .A2(G218gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n858_), .B2(new_n870_), .ZN(G1355gat));
endmodule


