//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_;
  INV_X1    g000(.A(KEYINPUT22), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G169gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT86), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT22), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT85), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT87), .B(G176gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n204_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT88), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT23), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n213_), .A2(KEYINPUT23), .ZN(new_n215_));
  MUX2_X1   g014(.A(new_n214_), .B(new_n215_), .S(KEYINPUT89), .Z(new_n216_));
  OR2_X1    g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n216_), .A2(new_n217_), .B1(G169gat), .B2(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT25), .B(G183gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  AOI22_X1  g022(.A1(new_n220_), .A2(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G176gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT24), .B1(new_n205_), .B2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n224_), .B(new_n214_), .C1(new_n223_), .C2(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n219_), .A2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G71gat), .B(G99gat), .Z(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G43gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n228_), .B(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G227gat), .A2(G233gat), .ZN(new_n232_));
  INV_X1    g031(.A(G15gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT30), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n231_), .B(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G127gat), .B(G134gat), .Z(new_n237_));
  XOR2_X1   g036(.A(G113gat), .B(G120gat), .Z(new_n238_));
  XOR2_X1   g037(.A(new_n237_), .B(new_n238_), .Z(new_n239_));
  INV_X1    g038(.A(KEYINPUT90), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n241_), .B(KEYINPUT31), .Z(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT91), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n236_), .A2(KEYINPUT92), .A3(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n231_), .A2(new_n235_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n231_), .A2(new_n235_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n242_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT92), .B1(new_n236_), .B2(new_n243_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT93), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n236_), .A2(new_n243_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT92), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT93), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(new_n247_), .A4(new_n244_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G211gat), .B(G218gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT96), .B(G204gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G197gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n259_), .B1(G197gat), .B2(G204gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n257_), .B1(new_n261_), .B2(KEYINPUT21), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT21), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(G197gat), .B2(G204gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(new_n258_), .B2(G197gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT97), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n262_), .A2(new_n266_), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n260_), .A2(new_n263_), .A3(new_n257_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n203_), .A2(new_n206_), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n270_), .B(KEYINPUT100), .Z(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n209_), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n214_), .A2(new_n217_), .B1(G169gat), .B2(G176gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n223_), .B1(new_n226_), .B2(KEYINPUT99), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(KEYINPUT99), .B2(new_n226_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n216_), .A2(new_n224_), .A3(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n269_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n278_), .A2(KEYINPUT101), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G226gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT19), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n282_), .B1(new_n278_), .B2(KEYINPUT101), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT20), .B1(new_n228_), .B2(new_n269_), .ZN(new_n284_));
  OR3_X1    g083(.A1(new_n279_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT20), .ZN(new_n286_));
  INV_X1    g085(.A(new_n269_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n274_), .A2(new_n277_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n286_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n228_), .A2(new_n269_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n282_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G8gat), .B(G36gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT102), .B(KEYINPUT18), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n285_), .A2(new_n292_), .A3(new_n298_), .ZN(new_n299_));
  NOR3_X1   g098(.A1(new_n279_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n297_), .B1(new_n300_), .B2(new_n291_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT27), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G78gat), .B(G106gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT3), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT2), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n312_), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n315_), .B(KEYINPUT94), .Z(new_n316_));
  OAI211_X1 g115(.A(new_n308_), .B(new_n309_), .C1(new_n314_), .C2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n307_), .B1(KEYINPUT1), .B2(new_n309_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(KEYINPUT1), .B2(new_n309_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n310_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n313_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n322_), .A2(KEYINPUT29), .ZN(new_n323_));
  NAND2_X1  g122(.A1(KEYINPUT95), .A2(G233gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(KEYINPUT95), .A2(G233gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(G228gat), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OR3_X1    g127(.A1(new_n323_), .A2(new_n269_), .A3(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n328_), .B1(new_n323_), .B2(new_n269_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n306_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(new_n330_), .A3(new_n306_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n322_), .A2(KEYINPUT29), .ZN(new_n335_));
  XOR2_X1   g134(.A(G22gat), .B(G50gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT28), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n335_), .B(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n331_), .B2(KEYINPUT98), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n332_), .A2(KEYINPUT98), .A3(new_n333_), .A4(new_n338_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n278_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n281_), .B1(new_n284_), .B2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n289_), .A2(new_n290_), .A3(new_n282_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n297_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n299_), .A2(KEYINPUT27), .A3(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n317_), .A2(new_n321_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n241_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n241_), .A2(new_n349_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n322_), .A2(new_n239_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT4), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT103), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n354_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n350_), .A2(new_n360_), .A3(new_n357_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G1gat), .B(G29gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(G85gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT0), .B(G57gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  NAND3_X1  g164(.A1(new_n359_), .A2(new_n361_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n365_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n358_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n361_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n367_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n304_), .A2(new_n342_), .A3(new_n348_), .A4(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n350_), .A2(new_n360_), .A3(new_n358_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n367_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n376_), .B1(new_n357_), .B2(new_n356_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT33), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n366_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n359_), .A2(KEYINPUT33), .A3(new_n361_), .A4(new_n365_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n379_), .A2(new_n299_), .A3(new_n301_), .A4(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n298_), .A2(KEYINPUT32), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n346_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n285_), .A2(new_n292_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n372_), .B(new_n383_), .C1(new_n384_), .C2(new_n382_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n342_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT104), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n374_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  AOI211_X1 g187(.A(KEYINPUT104), .B(new_n342_), .C1(new_n381_), .C2(new_n385_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n256_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT105), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n256_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n304_), .A2(new_n348_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n394_), .A2(new_n342_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n373_), .A3(new_n395_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n256_), .B(KEYINPUT105), .C1(new_n388_), .C2(new_n389_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n392_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G232gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT34), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT35), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n400_), .A2(KEYINPUT35), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT74), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT73), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT7), .ZN(new_n410_));
  INV_X1    g209(.A(G99gat), .ZN(new_n411_));
  INV_X1    g210(.A(G106gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G99gat), .A2(G106gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT6), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(G99gat), .A3(G106gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT8), .ZN(new_n422_));
  XOR2_X1   g221(.A(G85gat), .B(G92gat), .Z(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT64), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n417_), .A2(new_n419_), .A3(KEYINPUT64), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n415_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(KEYINPUT65), .A3(new_n423_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT8), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT65), .B1(new_n428_), .B2(new_n423_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n424_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT10), .B(G99gat), .Z(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n412_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n423_), .A2(KEYINPUT9), .ZN(new_n435_));
  INV_X1    g234(.A(G85gat), .ZN(new_n436_));
  INV_X1    g235(.A(G92gat), .ZN(new_n437_));
  OR3_X1    g236(.A1(new_n436_), .A2(new_n437_), .A3(KEYINPUT9), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n434_), .A2(new_n435_), .A3(new_n438_), .A4(new_n420_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n432_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G29gat), .B(G36gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G43gat), .B(G50gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n409_), .B1(new_n440_), .B2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n432_), .A2(KEYINPUT73), .A3(new_n443_), .A4(new_n439_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n408_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT69), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT68), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n432_), .A2(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(KEYINPUT68), .B(new_n424_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n448_), .B1(new_n452_), .B2(new_n439_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n439_), .ZN(new_n454_));
  AOI211_X1 g253(.A(KEYINPUT69), .B(new_n454_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n443_), .B(KEYINPUT15), .Z(new_n457_));
  OAI211_X1 g256(.A(new_n404_), .B(new_n447_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n451_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT65), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n417_), .A2(new_n419_), .A3(KEYINPUT64), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT64), .B1(new_n417_), .B2(new_n419_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n413_), .A2(new_n414_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n423_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n460_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(KEYINPUT8), .A3(new_n429_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT68), .B1(new_n467_), .B2(new_n424_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n439_), .B1(new_n459_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT69), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n452_), .A2(new_n448_), .A3(new_n439_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n457_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n447_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n403_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT76), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n458_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G190gat), .B(G218gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT75), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G134gat), .B(G162gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n458_), .A2(new_n474_), .A3(new_n480_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n476_), .A2(KEYINPUT36), .A3(new_n481_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n398_), .A2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G120gat), .B(G148gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G176gat), .B(G204gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G57gat), .B(G64gat), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n496_));
  XOR2_X1   g295(.A(G71gat), .B(G78gat), .Z(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n496_), .A2(new_n497_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  OR3_X1    g300(.A1(new_n440_), .A2(KEYINPUT66), .A3(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n500_), .B1(new_n432_), .B2(new_n439_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT66), .B1(new_n440_), .B2(new_n501_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(G230gat), .A2(G233gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT67), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n501_), .A2(KEYINPUT12), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n513_));
  XOR2_X1   g312(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n514_));
  NAND3_X1  g313(.A1(new_n504_), .A2(KEYINPUT71), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT71), .ZN(new_n516_));
  INV_X1    g315(.A(new_n514_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n516_), .B1(new_n503_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n440_), .A2(new_n501_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(new_n507_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n513_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n493_), .B1(new_n510_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n508_), .B(KEYINPUT67), .ZN(new_n525_));
  INV_X1    g324(.A(new_n493_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n522_), .A3(new_n526_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n524_), .A2(KEYINPUT13), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT13), .B1(new_n524_), .B2(new_n527_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT79), .B(G15gat), .ZN(new_n532_));
  INV_X1    g331(.A(G22gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT14), .ZN(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT81), .B(G8gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT80), .B(G1gat), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G1gat), .B(G8gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(new_n457_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT84), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n541_), .B2(new_n443_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n541_), .B(new_n443_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n543_), .A2(new_n546_), .B1(new_n547_), .B2(new_n545_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G113gat), .B(G141gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(G169gat), .B(G197gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n548_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n541_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n500_), .B(KEYINPUT82), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G127gat), .B(G155gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT16), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n561_), .A2(new_n562_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n557_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT83), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n557_), .A2(new_n563_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n565_), .A2(new_n566_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n531_), .A2(new_n553_), .A3(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n488_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n372_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(G1gat), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n398_), .A2(new_n552_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT78), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT37), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n487_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(KEYINPUT78), .A2(KEYINPUT37), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n579_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n485_), .A2(new_n486_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n530_), .A2(new_n580_), .A3(new_n571_), .A4(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n577_), .A2(new_n585_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n586_), .A2(new_n373_), .A3(new_n537_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n576_), .B1(new_n587_), .B2(KEYINPUT38), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(KEYINPUT38), .B2(new_n587_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT106), .ZN(G1324gat));
  NAND2_X1  g389(.A1(new_n574_), .A2(new_n394_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(G8gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT39), .ZN(new_n593_));
  INV_X1    g392(.A(new_n394_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n594_), .A2(new_n536_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n593_), .B1(new_n586_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT40), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(G1325gat));
  AOI21_X1  g397(.A(new_n233_), .B1(new_n574_), .B2(new_n393_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT41), .ZN(new_n600_));
  INV_X1    g399(.A(new_n586_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n233_), .A3(new_n393_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(G1326gat));
  AOI21_X1  g402(.A(new_n533_), .B1(new_n574_), .B2(new_n342_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT42), .Z(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n533_), .A3(new_n342_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(G1327gat));
  NOR2_X1   g406(.A1(new_n487_), .A2(new_n571_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n577_), .A2(new_n530_), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(G29gat), .B1(new_n609_), .B2(new_n372_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n580_), .A2(new_n583_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n398_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT43), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT43), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n398_), .A2(new_n614_), .A3(new_n611_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n531_), .A2(new_n553_), .A3(new_n571_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT44), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(KEYINPUT44), .A3(new_n617_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n372_), .A2(G29gat), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n610_), .B1(new_n622_), .B2(new_n623_), .ZN(G1328gat));
  NAND3_X1  g423(.A1(new_n620_), .A2(new_n394_), .A3(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G36gat), .ZN(new_n626_));
  INV_X1    g425(.A(G36gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n609_), .A2(new_n627_), .A3(new_n394_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT45), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT46), .Z(G1329gat));
  AOI21_X1  g430(.A(G43gat), .B1(new_n609_), .B2(new_n393_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT107), .Z(new_n633_));
  NAND3_X1  g432(.A1(new_n622_), .A2(G43gat), .A3(new_n393_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g435(.A(G50gat), .B1(new_n609_), .B2(new_n342_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n342_), .A2(G50gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n622_), .B2(new_n638_), .ZN(G1331gat));
  NAND4_X1  g438(.A1(new_n488_), .A2(new_n553_), .A3(new_n531_), .A4(new_n571_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(G57gat), .A3(new_n372_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT108), .Z(new_n643_));
  AND3_X1   g442(.A1(new_n398_), .A2(new_n553_), .A3(new_n531_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n580_), .A2(new_n571_), .A3(new_n583_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(G57gat), .B1(new_n646_), .B2(new_n372_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n643_), .A2(new_n647_), .ZN(G1332gat));
  OAI21_X1  g447(.A(G64gat), .B1(new_n640_), .B2(new_n594_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT48), .ZN(new_n650_));
  INV_X1    g449(.A(G64gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n646_), .A2(new_n651_), .A3(new_n394_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(G1333gat));
  OAI21_X1  g452(.A(G71gat), .B1(new_n640_), .B2(new_n256_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT49), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n256_), .A2(G71gat), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT109), .Z(new_n657_));
  NAND2_X1  g456(.A1(new_n646_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(G1334gat));
  INV_X1    g458(.A(new_n342_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G78gat), .B1(new_n640_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT50), .ZN(new_n662_));
  INV_X1    g461(.A(G78gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n646_), .A2(new_n663_), .A3(new_n342_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1335gat));
  AND2_X1   g464(.A1(new_n644_), .A2(new_n608_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G85gat), .B1(new_n666_), .B2(new_n372_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT110), .Z(new_n668_));
  NOR3_X1   g467(.A1(new_n530_), .A2(new_n552_), .A3(new_n571_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n373_), .A2(new_n436_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(G1336gat));
  NAND2_X1  g472(.A1(new_n616_), .A2(new_n669_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G92gat), .B1(new_n674_), .B2(new_n594_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n666_), .A2(new_n437_), .A3(new_n394_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT111), .Z(G1337gat));
  AOI21_X1  g477(.A(new_n411_), .B1(new_n671_), .B2(new_n393_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n393_), .A2(new_n433_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n666_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT112), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT51), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n681_), .B(new_n683_), .ZN(G1338gat));
  INV_X1    g483(.A(KEYINPUT114), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n671_), .A2(KEYINPUT113), .A3(new_n342_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G106gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT113), .B1(new_n671_), .B2(new_n342_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n685_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT113), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n690_), .B1(new_n674_), .B2(new_n660_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n691_), .A2(new_n686_), .A3(KEYINPUT114), .A4(G106gat), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n689_), .A2(KEYINPUT52), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT52), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n685_), .B(new_n694_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n666_), .A2(new_n412_), .A3(new_n342_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT53), .B1(new_n693_), .B2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n689_), .A2(KEYINPUT52), .A3(new_n692_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT53), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n695_), .A4(new_n696_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(G1339gat));
  AOI21_X1  g501(.A(new_n544_), .B1(new_n541_), .B2(new_n443_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n543_), .A2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n551_), .B1(new_n547_), .B2(new_n544_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n548_), .A2(new_n551_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n527_), .A2(new_n706_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n513_), .A2(new_n519_), .A3(new_n505_), .A4(new_n502_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n522_), .A2(KEYINPUT55), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT55), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n513_), .A2(new_n710_), .A3(new_n519_), .A4(new_n521_), .ZN(new_n711_));
  AOI221_X4 g510(.A(KEYINPUT116), .B1(new_n708_), .B2(new_n507_), .C1(new_n709_), .C2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT116), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n709_), .A2(new_n711_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n708_), .A2(new_n507_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n713_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n493_), .B1(new_n712_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT56), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n470_), .A2(new_n471_), .ZN(new_n720_));
  AOI22_X1  g519(.A1(new_n720_), .A2(new_n512_), .B1(new_n518_), .B2(new_n515_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n710_), .B1(new_n721_), .B2(new_n521_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n711_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n715_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT116), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n714_), .A2(new_n713_), .A3(new_n715_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(KEYINPUT56), .A3(new_n493_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n707_), .B1(new_n719_), .B2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT58), .B1(new_n729_), .B2(KEYINPUT117), .ZN(new_n730_));
  INV_X1    g529(.A(new_n707_), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT56), .B1(new_n727_), .B2(new_n493_), .ZN(new_n732_));
  AOI211_X1 g531(.A(new_n718_), .B(new_n526_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT117), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT58), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n730_), .A2(new_n737_), .A3(new_n611_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n527_), .A2(new_n552_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT115), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n527_), .A2(new_n552_), .A3(KEYINPUT115), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n719_), .B2(new_n728_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n524_), .A2(new_n527_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n706_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n487_), .B1(new_n744_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT57), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT57), .B(new_n487_), .C1(new_n744_), .C2(new_n747_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n738_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n572_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT54), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n645_), .A2(new_n754_), .A3(new_n553_), .A4(new_n530_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT54), .B1(new_n584_), .B2(new_n552_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n753_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT59), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n393_), .A2(new_n372_), .A3(new_n395_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(KEYINPUT121), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(KEYINPUT121), .B2(new_n760_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n758_), .A2(KEYINPUT122), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT122), .B1(new_n758_), .B2(new_n762_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT120), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n741_), .A2(new_n742_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n767_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n746_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT57), .B1(new_n769_), .B2(new_n487_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n751_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n571_), .B1(new_n772_), .B2(new_n738_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n757_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT118), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n753_), .A2(new_n776_), .A3(new_n757_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n760_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n766_), .B1(new_n778_), .B2(new_n759_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n760_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n776_), .B1(new_n753_), .B2(new_n757_), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT118), .B(new_n774_), .C1(new_n752_), .C2(new_n572_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n780_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n765_), .B1(new_n779_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(G113gat), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n553_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n778_), .A2(KEYINPUT119), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n783_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(new_n552_), .A3(new_n790_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n785_), .A2(new_n787_), .B1(new_n791_), .B2(new_n786_), .ZN(G1340gat));
  INV_X1    g591(.A(KEYINPUT60), .ZN(new_n793_));
  AOI21_X1  g592(.A(G120gat), .B1(new_n531_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n793_), .B2(G120gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n788_), .A2(new_n790_), .A3(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n531_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n779_), .B2(new_n784_), .ZN(new_n798_));
  INV_X1    g597(.A(G120gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n796_), .B1(new_n798_), .B2(new_n799_), .ZN(G1341gat));
  INV_X1    g599(.A(G127gat), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n572_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n788_), .A2(new_n571_), .A3(new_n790_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n785_), .A2(new_n802_), .B1(new_n803_), .B2(new_n801_), .ZN(G1342gat));
  INV_X1    g603(.A(new_n611_), .ZN(new_n805_));
  INV_X1    g604(.A(G134gat), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n487_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n788_), .A2(new_n808_), .A3(new_n790_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n785_), .A2(new_n807_), .B1(new_n809_), .B2(new_n806_), .ZN(G1343gat));
  NAND2_X1  g609(.A1(new_n775_), .A2(new_n777_), .ZN(new_n811_));
  NOR4_X1   g610(.A1(new_n393_), .A2(new_n660_), .A3(new_n373_), .A4(new_n394_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT123), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(KEYINPUT123), .B(new_n812_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(G141gat), .B1(new_n816_), .B2(new_n553_), .ZN(new_n817_));
  INV_X1    g616(.A(G141gat), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n552_), .C1(new_n813_), .C2(new_n815_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1344gat));
  OAI21_X1  g619(.A(G148gat), .B1(new_n816_), .B2(new_n530_), .ZN(new_n821_));
  INV_X1    g620(.A(G148gat), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(new_n531_), .C1(new_n813_), .C2(new_n815_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1345gat));
  XNOR2_X1  g623(.A(KEYINPUT61), .B(G155gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n816_), .B2(new_n572_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n825_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n571_), .B(new_n827_), .C1(new_n813_), .C2(new_n815_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1346gat));
  OAI21_X1  g628(.A(G162gat), .B1(new_n816_), .B2(new_n805_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n487_), .A2(G162gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1347gat));
  AOI21_X1  g632(.A(new_n342_), .B1(new_n753_), .B2(new_n757_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n256_), .A2(new_n372_), .A3(new_n594_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  AOI211_X1 g636(.A(KEYINPUT62), .B(new_n205_), .C1(new_n837_), .C2(new_n552_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT62), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n552_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(G169gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n837_), .A2(new_n271_), .A3(new_n552_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n838_), .B1(new_n841_), .B2(new_n842_), .ZN(G1348gat));
  NAND2_X1  g642(.A1(new_n837_), .A2(new_n531_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n342_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n835_), .A2(G176gat), .A3(new_n531_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n844_), .A2(new_n209_), .B1(new_n845_), .B2(new_n846_), .ZN(G1349gat));
  AND2_X1   g646(.A1(new_n835_), .A2(new_n571_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G183gat), .B1(new_n845_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n220_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n834_), .B2(new_n851_), .ZN(G1350gat));
  OAI21_X1  g651(.A(G190gat), .B1(new_n836_), .B2(new_n805_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n808_), .A2(new_n221_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n836_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1351gat));
  NOR4_X1   g656(.A1(new_n393_), .A2(new_n594_), .A3(new_n660_), .A4(new_n372_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n552_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G197gat), .ZN(G1352gat));
  OAI211_X1 g661(.A(new_n531_), .B(new_n858_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G204gat), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n530_), .A2(new_n258_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT125), .B1(new_n860_), .B2(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n858_), .B(new_n865_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n864_), .B1(new_n866_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT126), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT126), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n872_), .B(new_n864_), .C1(new_n866_), .C2(new_n869_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(G1353gat));
  NAND2_X1  g673(.A1(new_n860_), .A2(new_n571_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n876_));
  AND2_X1   g675(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n875_), .B2(new_n876_), .ZN(G1354gat));
  NAND2_X1  g678(.A1(new_n860_), .A2(new_n808_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G218gat), .B1(new_n881_), .B2(KEYINPUT127), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT127), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n883_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n611_), .A2(G218gat), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n882_), .A2(new_n884_), .B1(new_n860_), .B2(new_n885_), .ZN(G1355gat));
endmodule


