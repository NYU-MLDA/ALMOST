//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n798_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n828_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_;
  XOR2_X1   g000(.A(G120gat), .B(G148gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G176gat), .B(G204gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT75), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G57gat), .B(G64gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT11), .ZN(new_n209_));
  XOR2_X1   g008(.A(G71gat), .B(G78gat), .Z(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n208_), .A2(KEYINPUT11), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n210_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n211_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT12), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT73), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT72), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT69), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n221_));
  NAND2_X1  g020(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n222_));
  INV_X1    g021(.A(G99gat), .ZN(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n221_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n226_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n228_), .A2(KEYINPUT68), .A3(new_n222_), .A4(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT6), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT6), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(G99gat), .A3(G106gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n233_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n231_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G85gat), .ZN(new_n240_));
  INV_X1    g039(.A(G92gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT8), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G85gat), .A2(G92gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n220_), .B1(new_n239_), .B2(new_n246_), .ZN(new_n247_));
  AOI211_X1 g046(.A(KEYINPUT69), .B(new_n245_), .C1(new_n231_), .C2(new_n238_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT70), .B(KEYINPUT71), .Z(new_n250_));
  NAND2_X1  g049(.A1(new_n235_), .A2(new_n237_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n233_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n231_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n242_), .A2(new_n244_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n243_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n219_), .B1(new_n249_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n251_), .A2(new_n232_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(new_n227_), .B2(new_n230_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT69), .B1(new_n261_), .B2(new_n245_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n239_), .A2(new_n220_), .A3(new_n246_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n255_), .A2(new_n257_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT8), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n266_), .A3(KEYINPUT72), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n259_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT10), .B(G99gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT64), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT65), .B(G106gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT9), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n273_), .B(new_n242_), .C1(new_n256_), .C2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n257_), .A2(KEYINPUT66), .A3(KEYINPUT9), .ZN(new_n276_));
  AND4_X1   g075(.A1(new_n272_), .A2(new_n275_), .A3(new_n251_), .A4(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n218_), .B1(new_n268_), .B2(new_n278_), .ZN(new_n279_));
  AOI211_X1 g078(.A(KEYINPUT73), .B(new_n277_), .C1(new_n259_), .C2(new_n267_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n217_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n277_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n282_), .A2(new_n214_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(new_n215_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n214_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G230gat), .A2(G233gat), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n281_), .A2(new_n284_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n286_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n207_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT76), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n283_), .A2(new_n215_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n264_), .A2(KEYINPUT72), .A3(new_n266_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT72), .B1(new_n264_), .B2(new_n266_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n278_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT73), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n268_), .A2(new_n218_), .A3(new_n278_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n294_), .B1(new_n300_), .B2(new_n217_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n289_), .B1(new_n301_), .B2(new_n287_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n293_), .B1(new_n302_), .B2(new_n206_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n288_), .A2(new_n293_), .A3(new_n290_), .A4(new_n206_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n292_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT77), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n288_), .A2(new_n290_), .A3(new_n206_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT76), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n304_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(KEYINPUT77), .A3(new_n292_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n308_), .A2(KEYINPUT13), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT13), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT77), .B1(new_n311_), .B2(new_n292_), .ZN(new_n315_));
  AOI211_X1 g114(.A(new_n307_), .B(new_n291_), .C1(new_n310_), .C2(new_n304_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G29gat), .B(G36gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G43gat), .B(G50gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n321_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT15), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G15gat), .B(G22gat), .ZN(new_n326_));
  INV_X1    g125(.A(G1gat), .ZN(new_n327_));
  INV_X1    g126(.A(G8gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT14), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G1gat), .B(G8gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n325_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n332_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n324_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G229gat), .A2(G233gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT84), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n324_), .A2(new_n334_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n321_), .B(new_n322_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n340_), .A2(new_n332_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n338_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n332_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n335_), .A2(new_n343_), .A3(KEYINPUT84), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n336_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT85), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT85), .ZN(new_n348_));
  AOI211_X1 g147(.A(new_n348_), .B(new_n336_), .C1(new_n342_), .C2(new_n344_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n337_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G113gat), .B(G141gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G169gat), .B(G197gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n350_), .A2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n337_), .B(new_n353_), .C1(new_n347_), .C2(new_n349_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n356_), .A2(KEYINPUT86), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(KEYINPUT86), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n355_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT87), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n356_), .B(KEYINPUT86), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(KEYINPUT87), .A3(new_n355_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n318_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT19), .ZN(new_n368_));
  INV_X1    g167(.A(G197gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(G204gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT95), .ZN(new_n371_));
  INV_X1    g170(.A(G204gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(G197gat), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT94), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(KEYINPUT94), .A3(G197gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT96), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(G211gat), .B(G218gat), .Z(new_n380_));
  NAND4_X1  g179(.A1(new_n371_), .A2(KEYINPUT96), .A3(new_n375_), .A4(new_n376_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n379_), .A2(KEYINPUT21), .A3(new_n380_), .A4(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n370_), .A2(new_n373_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(KEYINPUT21), .B2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n384_), .B1(new_n377_), .B2(KEYINPUT21), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G183gat), .A2(G190gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n387_), .B(KEYINPUT23), .Z(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT26), .B(G190gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT25), .B(G183gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n392_), .B1(G169gat), .B2(G176gat), .ZN(new_n393_));
  NOR3_X1   g192(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n387_), .B(KEYINPUT23), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(G183gat), .B2(G190gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(G169gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n386_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT99), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT90), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n398_), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT90), .B1(G183gat), .B2(G190gat), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n406_), .B(new_n400_), .C1(new_n388_), .C2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT25), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(G183gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT89), .ZN(new_n411_));
  OR3_X1    g210(.A1(new_n409_), .A2(KEYINPUT88), .A3(G183gat), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT88), .B1(new_n409_), .B2(G183gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n389_), .A3(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n395_), .B(new_n397_), .C1(new_n411_), .C2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n408_), .A2(new_n415_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n386_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n404_), .A2(KEYINPUT20), .A3(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n403_), .A2(KEYINPUT99), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n368_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n386_), .A2(new_n402_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n386_), .A2(new_n416_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(KEYINPUT20), .A3(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n423_), .A2(new_n368_), .ZN(new_n424_));
  XOR2_X1   g223(.A(G8gat), .B(G36gat), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT101), .ZN(new_n426_));
  XOR2_X1   g225(.A(G64gat), .B(G92gat), .Z(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n420_), .A2(new_n424_), .A3(new_n430_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n431_), .A2(KEYINPUT106), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT20), .B1(new_n386_), .B2(new_n416_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(KEYINPUT99), .B2(new_n403_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n368_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n419_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n423_), .A2(new_n368_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n430_), .B(KEYINPUT105), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n433_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n431_), .A2(KEYINPUT106), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n432_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT107), .ZN(new_n445_));
  INV_X1    g244(.A(new_n430_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n436_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n423_), .A2(new_n368_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n431_), .A3(KEYINPUT102), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT102), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n451_), .B(new_n446_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n445_), .B1(new_n453_), .B2(KEYINPUT27), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n450_), .A2(KEYINPUT107), .A3(new_n433_), .A4(new_n452_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n444_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G141gat), .ZN(new_n457_));
  INV_X1    g256(.A(G148gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G141gat), .A2(G148gat), .ZN(new_n460_));
  INV_X1    g259(.A(G155gat), .ZN(new_n461_));
  INV_X1    g260(.A(G162gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT1), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n463_), .B1(G155gat), .B2(G162gat), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT1), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n459_), .B(new_n460_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G155gat), .B(G162gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n467_), .B(KEYINPUT92), .Z(new_n468_));
  OAI21_X1  g267(.A(new_n459_), .B1(KEYINPUT91), .B2(KEYINPUT3), .ZN(new_n469_));
  OR4_X1    g268(.A1(KEYINPUT91), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT2), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n460_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n473_));
  AND4_X1   g272(.A1(new_n469_), .A2(new_n470_), .A3(new_n472_), .A4(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n466_), .B1(new_n468_), .B2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G127gat), .B(G134gat), .Z(new_n476_));
  XNOR2_X1  g275(.A(G113gat), .B(G120gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n478_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G225gat), .A2(G233gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  OR3_X1    g283(.A1(new_n480_), .A2(KEYINPUT103), .A3(KEYINPUT4), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n479_), .A2(KEYINPUT4), .A3(new_n480_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT103), .B1(new_n480_), .B2(KEYINPUT4), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n484_), .B1(new_n483_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G1gat), .B(G29gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(G85gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT0), .B(G57gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n489_), .A2(new_n494_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  OR3_X1    g297(.A1(new_n475_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT28), .B1(new_n475_), .B2(KEYINPUT29), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G22gat), .B(G50gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT93), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n475_), .A2(KEYINPUT29), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n386_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G228gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G78gat), .B(G106gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT97), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n509_), .A2(new_n511_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT97), .B1(new_n509_), .B2(new_n511_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n505_), .B(new_n514_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n510_), .A2(KEYINPUT98), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n509_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n509_), .A2(new_n518_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n503_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G71gat), .B(G99gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(G43gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n416_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(new_n478_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G227gat), .A2(G233gat), .ZN(new_n528_));
  INV_X1    g327(.A(G15gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT30), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT31), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n527_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n456_), .A2(new_n498_), .A3(new_n523_), .A4(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT104), .B1(new_n489_), .B2(new_n494_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n536_), .A2(KEYINPUT33), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n488_), .A2(new_n483_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n493_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n536_), .A2(KEYINPUT33), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n453_), .A2(new_n537_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n430_), .A2(KEYINPUT32), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n420_), .A2(new_n424_), .A3(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n440_), .A2(KEYINPUT32), .A3(new_n430_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n497_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n522_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n523_), .A2(new_n497_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n456_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n535_), .B1(new_n548_), .B2(new_n534_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n366_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G134gat), .B(G162gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(KEYINPUT36), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n300_), .A2(new_n325_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT35), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT34), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  AOI22_X1  g359(.A1(new_n282_), .A2(new_n324_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n560_), .A2(new_n557_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n556_), .B(new_n561_), .C1(new_n557_), .C2(new_n560_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n555_), .B1(new_n566_), .B2(KEYINPUT80), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT80), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n564_), .A2(new_n568_), .A3(new_n565_), .A4(new_n554_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n553_), .A2(KEYINPUT36), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n566_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT37), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(KEYINPUT81), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(KEYINPUT81), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n573_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n567_), .A2(new_n569_), .B1(new_n566_), .B2(new_n571_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(KEYINPUT81), .A3(new_n574_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n332_), .B(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(new_n214_), .Z(new_n583_));
  OR2_X1    g382(.A1(new_n583_), .A2(KEYINPUT82), .ZN(new_n584_));
  XOR2_X1   g383(.A(G127gat), .B(G155gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT16), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT17), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n583_), .A2(KEYINPUT82), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n584_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT83), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n588_), .A2(new_n589_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n583_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n580_), .A2(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n550_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(new_n327_), .A3(new_n497_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT108), .B(KEYINPUT38), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n600_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n596_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n549_), .A2(new_n603_), .A3(new_n578_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n366_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G1gat), .B1(new_n605_), .B2(new_n498_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n601_), .A2(new_n602_), .A3(new_n606_), .ZN(G1324gat));
  OAI21_X1  g406(.A(G8gat), .B1(new_n605_), .B2(new_n456_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT39), .ZN(new_n609_));
  INV_X1    g408(.A(new_n456_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n598_), .A2(new_n328_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n612_), .B(new_n614_), .ZN(G1325gat));
  OAI21_X1  g414(.A(G15gat), .B1(new_n605_), .B2(new_n533_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT41), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n598_), .A2(new_n529_), .A3(new_n534_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT110), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(G1326gat));
  OAI21_X1  g421(.A(G22gat), .B1(new_n605_), .B2(new_n523_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT42), .ZN(new_n624_));
  INV_X1    g423(.A(G22gat), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n598_), .A2(new_n625_), .A3(new_n522_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(G1327gat));
  NOR2_X1   g426(.A1(new_n578_), .A2(new_n603_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT112), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n550_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(G29gat), .B1(new_n630_), .B2(new_n497_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n549_), .A2(new_n580_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n580_), .A2(KEYINPUT111), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(KEYINPUT43), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT43), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n549_), .B(new_n580_), .C1(KEYINPUT111), .C2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n318_), .A2(new_n603_), .A3(new_n365_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n637_), .A2(KEYINPUT44), .A3(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT44), .B1(new_n637_), .B2(new_n638_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n497_), .A2(G29gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n631_), .B1(new_n641_), .B2(new_n642_), .ZN(G1328gat));
  INV_X1    g442(.A(KEYINPUT46), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n639_), .A2(new_n640_), .A3(new_n456_), .ZN(new_n645_));
  INV_X1    g444(.A(G36gat), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n630_), .A2(new_n646_), .A3(new_n610_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT45), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n644_), .B1(new_n647_), .B2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n648_), .B(KEYINPUT45), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n652_), .B(KEYINPUT46), .C1(new_n646_), .C2(new_n645_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1329gat));
  XOR2_X1   g453(.A(KEYINPUT113), .B(G43gat), .Z(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n630_), .B2(new_n534_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n534_), .A2(G43gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n641_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT47), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(G1330gat));
  AOI21_X1  g459(.A(G50gat), .B1(new_n630_), .B2(new_n522_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n522_), .A2(G50gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n641_), .B2(new_n662_), .ZN(G1331gat));
  INV_X1    g462(.A(new_n318_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(new_n364_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n604_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(G57gat), .A3(new_n497_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT114), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(G57gat), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n665_), .A2(new_n549_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n597_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n672_), .B2(new_n498_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n669_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT115), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n669_), .A2(KEYINPUT115), .A3(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1332gat));
  INV_X1    g477(.A(G64gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n666_), .B2(new_n610_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT48), .Z(new_n681_));
  INV_X1    g480(.A(new_n672_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n679_), .A3(new_n610_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1333gat));
  INV_X1    g483(.A(G71gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n666_), .B2(new_n534_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT49), .Z(new_n687_));
  NAND3_X1  g486(.A1(new_n682_), .A2(new_n685_), .A3(new_n534_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1334gat));
  INV_X1    g488(.A(G78gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n666_), .B2(new_n522_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT50), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n682_), .A2(new_n690_), .A3(new_n522_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1335gat));
  NAND2_X1  g493(.A1(new_n665_), .A2(new_n596_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n636_), .B2(new_n634_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G85gat), .B1(new_n697_), .B2(new_n498_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n671_), .A2(new_n629_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n497_), .A2(new_n240_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(G1336gat));
  OAI21_X1  g500(.A(new_n241_), .B1(new_n699_), .B2(new_n456_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n610_), .A2(G92gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT116), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n697_), .B2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT117), .ZN(G1337gat));
  OAI21_X1  g505(.A(G99gat), .B1(new_n697_), .B2(new_n533_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n534_), .A2(new_n270_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n699_), .B2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g509(.A1(new_n671_), .A2(new_n271_), .A3(new_n522_), .A4(new_n629_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n224_), .B1(new_n696_), .B2(new_n522_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT52), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n712_), .A2(new_n713_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n711_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT53), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT53), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n718_), .B(new_n711_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1339gat));
  XNOR2_X1  g519(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n364_), .A2(new_n596_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n313_), .A2(new_n317_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT118), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n313_), .A2(new_n317_), .A3(new_n723_), .A4(KEYINPUT118), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n580_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n722_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  AOI211_X1 g529(.A(new_n580_), .B(new_n721_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n346_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n341_), .A2(new_n336_), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n353_), .B(new_n733_), .C1(new_n333_), .C2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n311_), .A2(new_n362_), .A3(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n281_), .A2(new_n285_), .A3(new_n284_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(G230gat), .A3(G233gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n301_), .A2(KEYINPUT55), .A3(new_n287_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT55), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n288_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n739_), .A2(new_n740_), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n207_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT56), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT56), .B1(new_n743_), .B2(new_n744_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n737_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT58), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n737_), .B(KEYINPUT58), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n580_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n745_), .A2(KEYINPUT120), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT121), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT120), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n743_), .A2(new_n756_), .A3(new_n744_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n754_), .A2(new_n755_), .A3(new_n746_), .A4(new_n757_), .ZN(new_n758_));
  AOI22_X1  g557(.A1(new_n361_), .A2(new_n363_), .B1(new_n310_), .B2(new_n304_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n743_), .A2(new_n756_), .A3(new_n744_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n756_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(KEYINPUT56), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT121), .B1(new_n745_), .B2(new_n746_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n758_), .B(new_n759_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n362_), .B(new_n736_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n573_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n753_), .B1(new_n766_), .B2(KEYINPUT57), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n768_), .B(new_n573_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n596_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n732_), .A2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n456_), .A2(new_n497_), .A3(new_n523_), .A4(new_n534_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT122), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(G113gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n364_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT59), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n774_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n771_), .A2(KEYINPUT59), .A3(new_n773_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n365_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n781_), .B2(new_n776_), .ZN(G1340gat));
  INV_X1    g581(.A(KEYINPUT60), .ZN(new_n783_));
  AOI21_X1  g582(.A(G120gat), .B1(new_n318_), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT123), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n783_), .B2(G120gat), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n771_), .A2(new_n786_), .A3(new_n773_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT124), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n664_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n789_));
  INV_X1    g588(.A(G120gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n788_), .B1(new_n789_), .B2(new_n790_), .ZN(G1341gat));
  INV_X1    g590(.A(G127gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n775_), .A2(new_n792_), .A3(new_n603_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n596_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(new_n792_), .ZN(G1342gat));
  INV_X1    g594(.A(G134gat), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n775_), .A2(new_n796_), .A3(new_n573_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n729_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(new_n796_), .ZN(G1343gat));
  NOR3_X1   g598(.A1(new_n523_), .A2(new_n498_), .A3(new_n534_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n771_), .A2(new_n456_), .A3(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(new_n365_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(new_n457_), .ZN(G1344gat));
  NOR2_X1   g602(.A1(new_n801_), .A2(new_n664_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(new_n458_), .ZN(G1345gat));
  NOR2_X1   g604(.A1(new_n801_), .A2(new_n596_), .ZN(new_n806_));
  XOR2_X1   g605(.A(KEYINPUT61), .B(G155gat), .Z(new_n807_));
  XNOR2_X1  g606(.A(new_n806_), .B(new_n807_), .ZN(G1346gat));
  OAI21_X1  g607(.A(G162gat), .B1(new_n801_), .B2(new_n729_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n573_), .A2(new_n462_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n801_), .B2(new_n810_), .ZN(G1347gat));
  NOR3_X1   g610(.A1(new_n522_), .A2(new_n497_), .A3(new_n533_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n771_), .A2(new_n364_), .A3(new_n610_), .A4(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT62), .ZN(new_n814_));
  AND4_X1   g613(.A1(KEYINPUT125), .A2(new_n813_), .A3(new_n814_), .A4(G169gat), .ZN(new_n815_));
  INV_X1    g614(.A(G169gat), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT125), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(KEYINPUT62), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n813_), .A2(new_n818_), .B1(KEYINPUT125), .B2(new_n814_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n456_), .B1(new_n732_), .B2(new_n770_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n812_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT22), .B(G169gat), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n364_), .A2(new_n822_), .ZN(new_n823_));
  XOR2_X1   g622(.A(new_n823_), .B(KEYINPUT126), .Z(new_n824_));
  OAI22_X1  g623(.A1(new_n815_), .A2(new_n819_), .B1(new_n821_), .B2(new_n824_), .ZN(G1348gat));
  NAND3_X1  g624(.A1(new_n820_), .A2(new_n318_), .A3(new_n812_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g626(.A1(new_n820_), .A2(new_n603_), .A3(new_n812_), .ZN(new_n828_));
  MUX2_X1   g627(.A(new_n390_), .B(G183gat), .S(new_n828_), .Z(G1350gat));
  OAI21_X1  g628(.A(G190gat), .B1(new_n821_), .B2(new_n729_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n573_), .A2(new_n389_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n821_), .B2(new_n831_), .ZN(G1351gat));
  NAND2_X1  g631(.A1(new_n547_), .A2(new_n533_), .ZN(new_n833_));
  AOI211_X1 g632(.A(new_n456_), .B(new_n833_), .C1(new_n732_), .C2(new_n770_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n364_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n318_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g637(.A1(new_n834_), .A2(new_n603_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT63), .B(G211gat), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n839_), .B2(new_n842_), .ZN(G1354gat));
  INV_X1    g642(.A(G218gat), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n834_), .B2(new_n580_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n833_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n578_), .A2(G218gat), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n820_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT127), .B1(new_n845_), .B2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n820_), .A2(new_n580_), .A3(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(G218gat), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT127), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n834_), .A2(new_n847_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n851_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n849_), .A2(new_n854_), .ZN(G1355gat));
endmodule


