//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n904_, new_n905_, new_n907_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(G127gat), .A2(G134gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G127gat), .A2(G134gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G113gat), .ZN(new_n206_));
  INV_X1    g005(.A(G120gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G113gat), .A2(G120gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n205_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n205_), .A2(new_n210_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT87), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT87), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(new_n217_), .B(KEYINPUT31), .Z(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT85), .B(G99gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G15gat), .B(G43gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT84), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G71gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n222_), .A2(G71gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n220_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n225_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n220_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n223_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G227gat), .ZN(new_n231_));
  INV_X1    g030(.A(G233gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n226_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(G169gat), .B(G176gat), .Z(new_n239_));
  AOI21_X1  g038(.A(new_n238_), .B1(new_n239_), .B2(KEYINPUT24), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT25), .B(G183gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT26), .B(G190gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(G183gat), .A3(G190gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G183gat), .ZN(new_n248_));
  INV_X1    g047(.A(G190gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT23), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n244_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n247_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n240_), .A2(new_n243_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n244_), .B1(G183gat), .B2(G190gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n245_), .A2(KEYINPUT83), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT83), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n257_), .A2(new_n244_), .A3(G183gat), .A4(G190gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n255_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n254_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  OR2_X1    g060(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G176gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT82), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT82), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n268_), .A3(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n253_), .B1(new_n261_), .B2(new_n270_), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n271_), .A2(KEYINPUT30), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(KEYINPUT30), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT86), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT88), .B1(new_n237_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n274_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT88), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n236_), .A4(new_n235_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n272_), .A2(KEYINPUT86), .A3(new_n273_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n279_), .B1(new_n275_), .B2(new_n278_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n219_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n275_), .A2(new_n278_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n279_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(new_n218_), .A3(new_n280_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n283_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G204gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G197gat), .ZN(new_n290_));
  INV_X1    g089(.A(G197gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G204gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT21), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT94), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n290_), .A2(new_n292_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT21), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G211gat), .B(G218gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT94), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n290_), .A2(new_n292_), .A3(new_n299_), .A4(new_n293_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n295_), .A2(new_n297_), .A3(new_n298_), .A4(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT95), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n297_), .A2(new_n298_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n293_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(KEYINPUT94), .B2(new_n294_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n300_), .A2(new_n298_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT95), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n302_), .A2(new_n303_), .A3(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT90), .ZN(new_n311_));
  OR2_X1    g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  AND3_X1   g111(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT89), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT89), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G141gat), .A3(G148gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n311_), .A2(new_n315_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT91), .B(KEYINPUT2), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT92), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n310_), .A2(KEYINPUT3), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n328_), .B1(G141gat), .B2(G148gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n316_), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n327_), .A2(new_n329_), .B1(new_n330_), .B2(KEYINPUT2), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n320_), .A2(KEYINPUT92), .A3(new_n323_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n326_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n312_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n322_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n309_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G228gat), .A2(G233gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(G78gat), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n309_), .B(new_n340_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n343_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n346_));
  INV_X1    g145(.A(G106gat), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n320_), .A2(KEYINPUT92), .A3(new_n323_), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT92), .B1(new_n320_), .B2(new_n323_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n327_), .A2(new_n329_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n330_), .A2(KEYINPUT2), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n349_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n321_), .B1(new_n354_), .B2(new_n335_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT29), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n340_), .B1(new_n356_), .B2(new_n309_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n344_), .ZN(new_n358_));
  OAI21_X1  g157(.A(G78gat), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n360_));
  AOI21_X1  g159(.A(G106gat), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT96), .B1(new_n348_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n347_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT96), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(G106gat), .A3(new_n360_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n337_), .A2(new_n338_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G22gat), .B(G50gat), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n362_), .A2(new_n366_), .A3(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n371_), .A2(new_n364_), .A3(new_n363_), .A4(new_n365_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n213_), .B(new_n321_), .C1(new_n354_), .C2(new_n335_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n376_), .B(KEYINPUT4), .C1(new_n217_), .C2(new_n337_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT100), .B(KEYINPUT4), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n355_), .A2(new_n214_), .A3(new_n216_), .A4(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n379_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT101), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n337_), .A2(new_n217_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(new_n213_), .B2(new_n337_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n378_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT101), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n377_), .A2(new_n387_), .A3(new_n379_), .A4(new_n381_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n383_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G1gat), .B(G29gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(G85gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT0), .ZN(new_n392_));
  INV_X1    g191(.A(G57gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n389_), .A2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n383_), .A2(new_n394_), .A3(new_n386_), .A4(new_n388_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT104), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(KEYINPUT104), .A3(new_n397_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT18), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(G64gat), .ZN(new_n404_));
  INV_X1    g203(.A(G92gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n301_), .A2(KEYINPUT95), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n307_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n260_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n252_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT98), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT98), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n252_), .A2(new_n413_), .A3(new_n410_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n264_), .A2(KEYINPUT97), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT97), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n265_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n412_), .A2(new_n254_), .A3(new_n414_), .A4(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n240_), .A2(new_n243_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n420_), .A2(new_n259_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n409_), .A2(new_n303_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT20), .B1(new_n309_), .B2(new_n271_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G226gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT19), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n422_), .A2(new_n423_), .A3(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n409_), .A2(new_n421_), .A3(new_n419_), .A4(new_n303_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT20), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n309_), .B2(new_n271_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n425_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n406_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n428_), .A2(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n426_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n419_), .A2(new_n421_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n309_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n309_), .A2(new_n271_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(KEYINPUT20), .A4(new_n425_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n406_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n434_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n432_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT27), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n422_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n426_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n432_), .B(KEYINPUT27), .C1(new_n446_), .C2(new_n406_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n400_), .A2(new_n401_), .A3(new_n443_), .A4(new_n447_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n288_), .A2(new_n375_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n375_), .A2(new_n448_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n373_), .A2(new_n374_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n432_), .A2(new_n440_), .A3(KEYINPUT99), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT99), .B1(new_n432_), .B2(new_n440_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n397_), .A2(KEYINPUT102), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT33), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT33), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n397_), .A2(KEYINPUT102), .A3(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n377_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT103), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n461_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n385_), .A2(new_n379_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n462_), .A2(new_n395_), .A3(new_n463_), .A4(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n455_), .A2(new_n457_), .A3(new_n459_), .A4(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n406_), .A2(KEYINPUT32), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n398_), .B(new_n468_), .C1(new_n446_), .C2(new_n467_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n452_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n470_));
  AND4_X1   g269(.A1(KEYINPUT105), .A2(new_n451_), .A3(new_n288_), .A4(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n283_), .A2(new_n287_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(new_n375_), .B2(new_n448_), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT105), .B1(new_n473_), .B2(new_n470_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n450_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G232gat), .A2(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT34), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G29gat), .B(G36gat), .ZN(new_n478_));
  INV_X1    g277(.A(G43gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(G50gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n478_), .B(G43gat), .ZN(new_n482_));
  INV_X1    g281(.A(G50gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G85gat), .B(G92gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT9), .ZN(new_n488_));
  XOR2_X1   g287(.A(KEYINPUT10), .B(G99gat), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n347_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT6), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT9), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(G85gat), .A3(G92gat), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n488_), .A2(new_n490_), .A3(new_n495_), .A4(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT8), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(KEYINPUT64), .ZN(new_n500_));
  NOR2_X1   g299(.A1(G99gat), .A2(G106gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT7), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT64), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n492_), .A2(new_n494_), .A3(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n499_), .B1(new_n505_), .B2(new_n487_), .ZN(new_n506_));
  AOI211_X1 g305(.A(KEYINPUT8), .B(new_n486_), .C1(new_n502_), .C2(new_n495_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n498_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT65), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(KEYINPUT65), .B(new_n498_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n485_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n481_), .A2(new_n484_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT15), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT15), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n485_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n502_), .A2(new_n495_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(new_n499_), .A3(new_n487_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n492_), .A2(new_n494_), .A3(new_n503_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n503_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n486_), .B1(new_n521_), .B2(new_n502_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n518_), .B1(new_n522_), .B2(new_n499_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n514_), .A2(new_n516_), .B1(new_n523_), .B2(new_n498_), .ZN(new_n524_));
  OAI211_X1 g323(.A(KEYINPUT35), .B(new_n477_), .C1(new_n512_), .C2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT65), .B1(new_n523_), .B2(new_n498_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n511_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n513_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n477_), .A2(KEYINPUT35), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n477_), .A2(KEYINPUT35), .ZN(new_n530_));
  INV_X1    g329(.A(new_n516_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n485_), .A2(new_n515_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n508_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .A4(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n525_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G190gat), .B(G218gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(G134gat), .ZN(new_n537_));
  INV_X1    g336(.A(G162gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n540_), .A2(KEYINPUT36), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(KEYINPUT36), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n525_), .A2(new_n534_), .A3(new_n541_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n475_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT106), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G127gat), .B(G155gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT16), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(new_n248_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(G211gat), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G1gat), .B(G8gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT75), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G15gat), .B(G22gat), .ZN(new_n557_));
  INV_X1    g356(.A(G8gat), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n556_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n560_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n563_), .B(new_n564_), .Z(new_n565_));
  XNOR2_X1  g364(.A(G57gat), .B(G64gat), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n566_), .A2(KEYINPUT11), .ZN(new_n567_));
  XOR2_X1   g366(.A(G71gat), .B(G78gat), .Z(new_n568_));
  OR2_X1    g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n568_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n569_), .B(new_n570_), .C1(KEYINPUT11), .C2(new_n566_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT68), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n565_), .B(new_n572_), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n571_), .B(KEYINPUT66), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n565_), .B(new_n574_), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n552_), .B(new_n553_), .ZN(new_n576_));
  OAI22_X1  g375(.A1(new_n554_), .A2(new_n573_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT76), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n548_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G230gat), .A2(G233gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n510_), .A2(new_n511_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n574_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT67), .Z(new_n583_));
  OR2_X1    g382(.A1(new_n581_), .A2(new_n574_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n580_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT12), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n572_), .A2(KEYINPUT12), .A3(new_n508_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n588_), .A2(KEYINPUT69), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(KEYINPUT69), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n582_), .A2(new_n580_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT70), .Z(new_n593_));
  AOI21_X1  g392(.A(new_n585_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT5), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G176gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(G204gat), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(KEYINPUT71), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n599_), .B1(new_n594_), .B2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n602_), .A2(KEYINPUT13), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(KEYINPUT13), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n563_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT78), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n563_), .A2(new_n513_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT79), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n563_), .B(new_n513_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(G229gat), .A3(G233gat), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT77), .Z(new_n616_));
  NAND2_X1  g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G113gat), .B(G141gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT80), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(G169gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(new_n291_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n621_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n613_), .A2(new_n616_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n605_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n579_), .A2(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n396_), .A2(KEYINPUT104), .A3(new_n397_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT104), .B1(new_n396_), .B2(new_n397_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n202_), .B1(new_n627_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT107), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT105), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n443_), .A2(new_n447_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n628_), .A2(new_n629_), .A3(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n288_), .B1(new_n636_), .B2(new_n452_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n452_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n473_), .A2(KEYINPUT105), .A3(new_n470_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n449_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n626_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n545_), .A2(KEYINPUT72), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT72), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n525_), .A2(new_n534_), .A3(new_n644_), .A4(new_n541_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n544_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT37), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT73), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n546_), .A2(KEYINPUT37), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT73), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n646_), .A2(new_n650_), .A3(KEYINPUT37), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n649_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT74), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n648_), .A2(KEYINPUT74), .A3(new_n649_), .A4(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n578_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n642_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n202_), .A3(new_n631_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT38), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n633_), .A2(new_n662_), .ZN(G1324gat));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n664_));
  INV_X1    g463(.A(new_n626_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n548_), .A2(new_n665_), .A3(new_n578_), .A4(new_n635_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n666_), .A2(G8gat), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(new_n668_), .B2(new_n667_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n660_), .A2(new_n558_), .A3(new_n635_), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n667_), .A2(new_n668_), .A3(KEYINPUT39), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n670_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT109), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT109), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n670_), .A2(new_n675_), .A3(new_n671_), .A4(new_n672_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n674_), .A2(KEYINPUT40), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT40), .B1(new_n674_), .B2(new_n676_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1325gat));
  INV_X1    g478(.A(G15gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n627_), .B2(new_n472_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT41), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n660_), .A2(new_n680_), .A3(new_n472_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1326gat));
  INV_X1    g483(.A(G22gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n627_), .B2(new_n375_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT42), .Z(new_n687_));
  NAND3_X1  g486(.A1(new_n660_), .A2(new_n685_), .A3(new_n375_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1327gat));
  NOR2_X1   g488(.A1(new_n578_), .A2(new_n546_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n642_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n631_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT111), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n639_), .A2(new_n640_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n656_), .B1(new_n695_), .B2(new_n450_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n694_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NOR4_X1   g497(.A1(new_n641_), .A2(KEYINPUT110), .A3(KEYINPUT43), .A4(new_n656_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n475_), .B2(new_n657_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n626_), .A2(new_n578_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n693_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n475_), .A2(new_n697_), .A3(new_n657_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT110), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n641_), .B2(new_n656_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n696_), .A2(new_n694_), .A3(new_n697_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(KEYINPUT111), .A3(new_n702_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n704_), .A2(new_n705_), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n704_), .A2(KEYINPUT112), .A3(new_n705_), .A4(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n710_), .A2(KEYINPUT44), .A3(new_n702_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n717_), .A2(G29gat), .A3(new_n631_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n692_), .B1(new_n716_), .B2(new_n718_), .ZN(G1328gat));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n635_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n710_), .A2(KEYINPUT111), .A3(new_n702_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT111), .B1(new_n710_), .B2(new_n702_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT112), .B1(new_n724_), .B2(new_n705_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n715_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n721_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT113), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n728_), .A3(G36gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n720_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT113), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n691_), .A2(new_n731_), .A3(new_n635_), .ZN(new_n733_));
  XOR2_X1   g532(.A(KEYINPUT114), .B(KEYINPUT45), .Z(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n729_), .A2(new_n732_), .A3(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT115), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n737_), .A3(KEYINPUT46), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT46), .B1(new_n736_), .B2(new_n737_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1329gat));
  NAND4_X1  g539(.A1(new_n716_), .A2(G43gat), .A3(new_n472_), .A4(new_n717_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n691_), .A2(new_n472_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(G43gat), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g543(.A(G50gat), .B1(new_n691_), .B2(new_n375_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n716_), .A2(G50gat), .A3(new_n717_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(new_n375_), .ZN(G1331gat));
  NOR2_X1   g546(.A1(new_n605_), .A2(new_n625_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n641_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n659_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G57gat), .B1(new_n751_), .B2(new_n631_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n579_), .A2(new_n749_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n630_), .A2(new_n393_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(G1332gat));
  INV_X1    g554(.A(G64gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n753_), .B2(new_n635_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT48), .Z(new_n758_));
  NAND3_X1  g557(.A1(new_n751_), .A2(new_n756_), .A3(new_n635_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1333gat));
  INV_X1    g559(.A(G71gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n753_), .B2(new_n472_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT49), .Z(new_n763_));
  NAND3_X1  g562(.A1(new_n751_), .A2(new_n761_), .A3(new_n472_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1334gat));
  AOI21_X1  g564(.A(new_n343_), .B1(new_n753_), .B2(new_n375_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT50), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n751_), .A2(new_n343_), .A3(new_n375_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1335gat));
  NAND3_X1  g568(.A1(new_n710_), .A2(new_n658_), .A3(new_n748_), .ZN(new_n770_));
  INV_X1    g569(.A(G85gat), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n770_), .A2(new_n771_), .A3(new_n630_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n750_), .A2(new_n690_), .ZN(new_n773_));
  AOI21_X1  g572(.A(G85gat), .B1(new_n773_), .B2(new_n631_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1336gat));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n405_), .A3(new_n635_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n770_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(new_n405_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT116), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n770_), .B2(new_n288_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n773_), .A2(new_n489_), .A3(new_n472_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g582(.A(G106gat), .B1(new_n770_), .B2(new_n452_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT52), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n785_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n786_), .B(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n773_), .A2(new_n347_), .A3(new_n375_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT117), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g591(.A1(new_n593_), .A2(new_n591_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n580_), .B1(new_n591_), .B2(new_n583_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n600_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT56), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n614_), .A2(new_n611_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n610_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n621_), .B(new_n799_), .C1(new_n800_), .C2(new_n611_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n624_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n803_), .B(new_n600_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n798_), .A2(new_n802_), .A3(new_n599_), .A4(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT58), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT121), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n806_), .A2(KEYINPUT121), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n657_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT122), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(KEYINPUT122), .A3(new_n657_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n812_), .B(new_n813_), .C1(new_n806_), .C2(new_n805_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n802_), .A2(new_n602_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n798_), .A2(new_n599_), .A3(new_n804_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n625_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(KEYINPUT57), .A3(new_n546_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n546_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT119), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n818_), .A2(new_n823_), .A3(new_n546_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(new_n822_), .A3(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n814_), .A2(new_n819_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n658_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n659_), .A2(new_n817_), .A3(new_n605_), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT54), .Z(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n630_), .A2(new_n635_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n452_), .A3(new_n472_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(KEYINPUT59), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n825_), .A2(KEYINPUT120), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n821_), .A2(new_n837_), .A3(new_n822_), .A4(new_n824_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n836_), .A2(new_n819_), .A3(new_n814_), .A4(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n829_), .B1(new_n839_), .B2(new_n658_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n833_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n835_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n843_), .A2(new_n206_), .A3(new_n817_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n840_), .A2(new_n817_), .A3(new_n833_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(G113gat), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(KEYINPUT123), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n845_), .A2(new_n848_), .A3(G113gat), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n844_), .A2(new_n847_), .A3(new_n849_), .ZN(G1340gat));
  OAI21_X1  g649(.A(G120gat), .B1(new_n843_), .B2(new_n605_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n207_), .B1(new_n605_), .B2(KEYINPUT60), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n841_), .B(new_n852_), .C1(KEYINPUT60), .C2(new_n207_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1341gat));
  AOI21_X1  g653(.A(G127gat), .B1(new_n841_), .B2(new_n578_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n843_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n578_), .A2(G127gat), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(G1342gat));
  INV_X1    g657(.A(new_n546_), .ZN(new_n859_));
  AOI21_X1  g658(.A(G134gat), .B1(new_n841_), .B2(new_n859_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n657_), .A2(G134gat), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n856_), .B2(new_n861_), .ZN(G1343gat));
  NOR3_X1   g661(.A1(new_n840_), .A2(new_n452_), .A3(new_n472_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(new_n625_), .A3(new_n832_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g664(.A(new_n605_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n863_), .A2(new_n866_), .A3(new_n832_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g667(.A1(new_n863_), .A2(new_n578_), .A3(new_n832_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT61), .B(G155gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1346gat));
  AND2_X1   g670(.A1(new_n863_), .A2(new_n832_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n859_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n656_), .A2(new_n538_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n873_), .A2(new_n538_), .B1(new_n872_), .B2(new_n874_), .ZN(G1347gat));
  AND2_X1   g674(.A1(new_n630_), .A2(new_n635_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n472_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n827_), .B2(new_n830_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n452_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT124), .B1(new_n879_), .B2(new_n817_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n878_), .A2(new_n881_), .A3(new_n625_), .A4(new_n452_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(G169gat), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n879_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n886_), .B(new_n625_), .C1(new_n417_), .C2(new_n415_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n880_), .A2(new_n882_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n885_), .A2(new_n887_), .A3(new_n888_), .ZN(G1348gat));
  INV_X1    g688(.A(KEYINPUT126), .ZN(new_n890_));
  OR3_X1    g689(.A1(new_n840_), .A2(new_n890_), .A3(new_n375_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n877_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n840_), .B2(new_n375_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n891_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n605_), .A2(new_n265_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n265_), .B1(new_n879_), .B2(new_n605_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  OAI211_X1 g697(.A(KEYINPUT125), .B(new_n265_), .C1(new_n879_), .C2(new_n605_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n894_), .A2(new_n895_), .B1(new_n898_), .B2(new_n899_), .ZN(G1349gat));
  NOR3_X1   g699(.A1(new_n879_), .A2(new_n658_), .A3(new_n241_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n891_), .A2(new_n578_), .A3(new_n892_), .A4(new_n893_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n248_), .ZN(G1350gat));
  OAI21_X1  g702(.A(G190gat), .B1(new_n879_), .B2(new_n656_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n859_), .A2(new_n242_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n879_), .B2(new_n905_), .ZN(G1351gat));
  NAND3_X1  g705(.A1(new_n863_), .A2(new_n625_), .A3(new_n876_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g707(.A1(new_n863_), .A2(new_n866_), .A3(new_n876_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n909_), .B(new_n910_), .Z(G1353gat));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n863_), .A2(new_n876_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n658_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT63), .B(G211gat), .Z(new_n915_));
  NAND4_X1  g714(.A1(new_n863_), .A2(new_n578_), .A3(new_n876_), .A4(new_n915_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1354gat));
  INV_X1    g716(.A(G218gat), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n913_), .A2(new_n918_), .A3(new_n656_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n863_), .A2(new_n859_), .A3(new_n876_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n918_), .B2(new_n920_), .ZN(G1355gat));
endmodule


