//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_;
  XNOR2_X1  g000(.A(KEYINPUT86), .B(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G228gat), .ZN(new_n204_));
  INV_X1    g003(.A(G233gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT85), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G22gat), .B(G50gat), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n208_), .B(new_n209_), .Z(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G155gat), .B(G162gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n216_), .A2(KEYINPUT2), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n217_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n220_), .B2(KEYINPUT81), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n215_), .B(KEYINPUT80), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n219_), .B(new_n221_), .C1(new_n222_), .C2(KEYINPUT2), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT82), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n214_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(new_n215_), .B(KEYINPUT80), .Z(new_n226_));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n228_), .A2(KEYINPUT82), .A3(new_n221_), .A4(new_n219_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n217_), .B1(new_n231_), .B2(KEYINPUT1), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n226_), .B(new_n232_), .C1(KEYINPUT1), .C2(new_n214_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n213_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(new_n233_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n237_), .A2(KEYINPUT29), .A3(new_n212_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n211_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n234_), .A2(new_n235_), .A3(new_n213_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n212_), .B1(new_n237_), .B2(KEYINPUT29), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n241_), .A3(new_n210_), .ZN(new_n242_));
  INV_X1    g041(.A(G78gat), .ZN(new_n243_));
  INV_X1    g042(.A(G197gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(G204gat), .ZN(new_n245_));
  INV_X1    g044(.A(G204gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(G197gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT21), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G211gat), .B(G218gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT84), .B1(new_n244_), .B2(G204gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT84), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(new_n246_), .A3(G197gat), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n250_), .B(new_n252_), .C1(G197gat), .C2(new_n246_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n248_), .B(new_n249_), .C1(new_n253_), .C2(KEYINPUT21), .ZN(new_n254_));
  INV_X1    g053(.A(new_n249_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(KEYINPUT21), .A3(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(new_n207_), .B2(new_n206_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n243_), .B(new_n258_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n235_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n257_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n206_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n261_), .B1(KEYINPUT85), .B2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(G78gat), .B1(new_n260_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n264_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n239_), .A2(new_n242_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n265_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n203_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n239_), .A2(new_n242_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n265_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n239_), .A2(new_n242_), .A3(new_n265_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n202_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n268_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT27), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT19), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT23), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT24), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT25), .B(G183gat), .ZN(new_n285_));
  INV_X1    g084(.A(G190gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT78), .B1(new_n286_), .B2(KEYINPUT26), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G190gat), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n285_), .B(new_n287_), .C1(new_n288_), .C2(KEYINPUT78), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT24), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n284_), .B(new_n289_), .C1(new_n291_), .C2(new_n281_), .ZN(new_n292_));
  INV_X1    g091(.A(G183gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n286_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n280_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT22), .B(G169gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT79), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G169gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n297_), .B1(new_n299_), .B2(KEYINPUT22), .ZN(new_n300_));
  INV_X1    g099(.A(G176gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n295_), .B(new_n290_), .C1(new_n298_), .C2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n257_), .A2(new_n292_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT87), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(KEYINPUT20), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n305_), .B1(new_n304_), .B2(KEYINPUT20), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n296_), .A2(new_n301_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n290_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT89), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n295_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n280_), .A2(KEYINPUT89), .A3(new_n294_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT90), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n315_), .A2(new_n316_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n291_), .A2(KEYINPUT88), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n291_), .A2(KEYINPUT88), .ZN(new_n321_));
  NOR3_X1   g120(.A1(new_n320_), .A2(new_n321_), .A3(new_n281_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n288_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n285_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n284_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  OAI22_X1  g124(.A1(new_n318_), .A2(new_n319_), .B1(new_n322_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n261_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n278_), .B1(new_n309_), .B2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G8gat), .B(G36gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n292_), .A2(new_n303_), .ZN(new_n334_));
  OAI211_X1 g133(.A(KEYINPUT20), .B(new_n278_), .C1(new_n334_), .C2(new_n257_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n325_), .A2(new_n322_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n315_), .A2(new_n316_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(new_n317_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n335_), .B1(new_n338_), .B2(new_n257_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n328_), .A2(new_n333_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n333_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n304_), .A2(KEYINPUT20), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT87), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n343_), .B(new_n306_), .C1(new_n338_), .C2(new_n257_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n277_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n339_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n341_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n275_), .B1(new_n340_), .B2(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G127gat), .B(G134gat), .Z(new_n349_));
  XOR2_X1   g148(.A(G113gat), .B(G120gat), .Z(new_n350_));
  XOR2_X1   g149(.A(new_n349_), .B(new_n350_), .Z(new_n351_));
  NAND2_X1  g150(.A1(new_n237_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n351_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n230_), .A2(new_n353_), .A3(new_n233_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(KEYINPUT4), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n353_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n354_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n361_), .A2(new_n357_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n356_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G1gat), .B(G29gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G57gat), .B(G85gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n369_), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n355_), .A2(new_n359_), .B1(new_n362_), .B2(new_n356_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n369_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G227gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(G15gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT30), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT31), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n292_), .A2(new_n303_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G71gat), .B(G99gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G43gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n381_), .B(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n353_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n384_), .A2(new_n353_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n380_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n387_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n379_), .A3(new_n385_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n374_), .A2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT20), .B1(new_n334_), .B2(new_n257_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n261_), .A2(new_n336_), .A3(new_n315_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n277_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n344_), .B2(new_n277_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n333_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n345_), .A2(new_n341_), .A3(new_n346_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(KEYINPUT27), .A3(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n274_), .A2(new_n348_), .A3(new_n392_), .A4(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT96), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n348_), .A2(new_n399_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n403_), .A2(new_n374_), .A3(new_n274_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT95), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n333_), .B1(new_n328_), .B2(new_n339_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT33), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n407_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n408_));
  AND4_X1   g207(.A1(new_n407_), .A2(new_n360_), .A3(new_n363_), .A4(new_n372_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n406_), .B(new_n398_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT93), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n361_), .B2(new_n357_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n352_), .A2(KEYINPUT93), .A3(new_n354_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n356_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(KEYINPUT94), .A3(new_n369_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT94), .B1(new_n415_), .B2(new_n369_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n414_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n355_), .A2(new_n419_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n417_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n405_), .B1(new_n410_), .B2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n418_), .A2(new_n420_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n416_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n373_), .A2(KEYINPUT33), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n371_), .A2(new_n407_), .A3(new_n372_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n340_), .A2(new_n347_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n424_), .A2(new_n427_), .A3(new_n428_), .A4(KEYINPUT95), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n396_), .A2(KEYINPUT32), .A3(new_n341_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n341_), .A2(KEYINPUT32), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n345_), .A2(new_n346_), .A3(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n374_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n422_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n404_), .B1(new_n434_), .B2(new_n274_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n391_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n402_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G190gat), .B(G218gat), .Z(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT70), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G134gat), .B(G162gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT36), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G99gat), .A2(G106gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT6), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(G99gat), .A3(G106gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  OR2_X1    g247(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n449_));
  INV_X1    g248(.A(G106gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G85gat), .ZN(new_n453_));
  INV_X1    g252(.A(G92gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G85gat), .A2(G92gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(KEYINPUT9), .A3(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n456_), .A2(KEYINPUT9), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n448_), .A2(new_n452_), .A3(new_n457_), .A4(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G99gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n450_), .A3(KEYINPUT64), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT7), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT7), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n464_), .A2(new_n461_), .A3(new_n450_), .A4(KEYINPUT64), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n448_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n455_), .A2(new_n456_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n466_), .A2(new_n470_), .A3(new_n468_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n460_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G29gat), .B(G36gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  XOR2_X1   g275(.A(G43gat), .B(G50gat), .Z(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G43gat), .B(G50gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT35), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G232gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT34), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n474_), .A2(new_n481_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n481_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n478_), .A2(KEYINPUT15), .A3(new_n480_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n474_), .A2(new_n490_), .A3(KEYINPUT69), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT69), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n488_), .A2(new_n489_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n466_), .A2(new_n470_), .A3(new_n468_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n470_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n459_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n492_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n486_), .B1(new_n491_), .B2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n485_), .A2(new_n482_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT69), .B1(new_n474_), .B2(new_n490_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n493_), .A2(new_n496_), .A3(new_n492_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n499_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n504_), .A3(new_n486_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n443_), .B1(new_n500_), .B2(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n506_), .A2(KEYINPUT72), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT36), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n500_), .A2(new_n508_), .A3(new_n505_), .A4(new_n441_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(KEYINPUT72), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n507_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n437_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G230gat), .A2(G233gat), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT11), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n243_), .A2(G71gat), .ZN(new_n515_));
  INV_X1    g314(.A(G71gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(G78gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(G57gat), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(G64gat), .ZN(new_n520_));
  INV_X1    g319(.A(G64gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(G57gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT66), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(G57gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n519_), .A2(G64gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT66), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  AOI211_X1 g326(.A(new_n514_), .B(new_n518_), .C1(new_n523_), .C2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n518_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n523_), .A2(new_n527_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n529_), .B1(new_n530_), .B2(KEYINPUT11), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n523_), .A2(new_n514_), .A3(new_n527_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n528_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n496_), .A2(new_n533_), .B1(KEYINPUT67), .B2(KEYINPUT12), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n526_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT11), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(new_n532_), .A3(new_n518_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n530_), .A2(KEYINPUT11), .A3(new_n529_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n496_), .B(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(KEYINPUT67), .B(KEYINPUT12), .Z(new_n543_));
  OAI211_X1 g342(.A(new_n513_), .B(new_n535_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n496_), .A2(new_n533_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n472_), .A2(new_n473_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(new_n541_), .A3(new_n459_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n513_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G120gat), .B(G148gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT5), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G176gat), .B(G204gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n544_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT68), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n545_), .A2(new_n547_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n543_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n534_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n548_), .B1(new_n560_), .B2(new_n513_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(KEYINPUT68), .A3(new_n554_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n561_), .A2(new_n554_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n563_), .A2(KEYINPUT13), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT13), .B1(new_n563_), .B2(new_n565_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G15gat), .B(G22gat), .ZN(new_n570_));
  INV_X1    g369(.A(G1gat), .ZN(new_n571_));
  INV_X1    g370(.A(G8gat), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT14), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n570_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n573_), .A2(new_n574_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G1gat), .B(G8gat), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n577_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n481_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT76), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n481_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n583_));
  OR3_X1    g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n582_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n584_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n578_), .A2(new_n579_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n493_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n585_), .A3(new_n580_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G113gat), .B(G141gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT77), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G169gat), .B(G197gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n592_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n588_), .A2(new_n591_), .A3(new_n596_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n569_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n589_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(new_n533_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT75), .ZN(new_n607_));
  XOR2_X1   g406(.A(G127gat), .B(G155gat), .Z(new_n608_));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n607_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n606_), .A2(new_n612_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT17), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT17), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n617_), .B1(new_n618_), .B2(new_n614_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n603_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n512_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n374_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT97), .Z(new_n625_));
  AND2_X1   g424(.A1(new_n437_), .A2(new_n600_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT37), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n507_), .A2(new_n510_), .A3(new_n627_), .A4(new_n509_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT71), .ZN(new_n629_));
  INV_X1    g428(.A(new_n505_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n504_), .B1(new_n503_), .B2(new_n486_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n442_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n509_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n629_), .B1(new_n633_), .B2(KEYINPUT37), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT71), .B(new_n627_), .C1(new_n632_), .C2(new_n509_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n628_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n619_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(new_n569_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n626_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n571_), .A3(new_n374_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT38), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n625_), .A2(new_n642_), .ZN(G1324gat));
  INV_X1    g442(.A(new_n403_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G8gat), .B1(new_n622_), .B2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT39), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n640_), .A2(new_n572_), .A3(new_n403_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g448(.A(G15gat), .B1(new_n622_), .B2(new_n391_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT41), .Z(new_n651_));
  NAND3_X1  g450(.A1(new_n640_), .A2(new_n376_), .A3(new_n436_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1326gat));
  OAI21_X1  g452(.A(G22gat), .B1(new_n622_), .B2(new_n274_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT42), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n274_), .A2(G22gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n639_), .B2(new_n656_), .ZN(G1327gat));
  NOR2_X1   g456(.A1(new_n619_), .A2(new_n511_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n568_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n626_), .A2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G29gat), .B1(new_n660_), .B2(new_n374_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n662_));
  INV_X1    g461(.A(new_n636_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n437_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT98), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n437_), .A2(new_n666_), .A3(new_n662_), .A4(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n437_), .A2(new_n663_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT43), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n665_), .A2(new_n667_), .A3(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n603_), .A2(new_n619_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n670_), .A2(KEYINPUT44), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT44), .B1(new_n670_), .B2(new_n671_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n374_), .A2(G29gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n661_), .B1(new_n674_), .B2(new_n675_), .ZN(G1328gat));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT100), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n644_), .A2(G36gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n626_), .A2(new_n659_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT99), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT99), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n626_), .A2(new_n683_), .A3(new_n659_), .A4(new_n679_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n681_), .A2(new_n682_), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n682_), .B1(new_n681_), .B2(new_n684_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n678_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n674_), .A2(new_n403_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(G36gat), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n677_), .A2(KEYINPUT100), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1329gat));
  AOI21_X1  g490(.A(G43gat), .B1(new_n660_), .B2(new_n436_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT102), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n694_));
  INV_X1    g493(.A(G43gat), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n391_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n674_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n696_), .ZN(new_n698_));
  NOR4_X1   g497(.A1(new_n672_), .A2(new_n673_), .A3(KEYINPUT101), .A4(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n693_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT47), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n702_), .B(new_n693_), .C1(new_n697_), .C2(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1330gat));
  INV_X1    g503(.A(G50gat), .ZN(new_n705_));
  INV_X1    g504(.A(new_n274_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n660_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n674_), .A2(new_n706_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n708_), .A2(KEYINPUT103), .A3(G50gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT103), .B1(new_n708_), .B2(G50gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n709_), .B2(new_n710_), .ZN(G1331gat));
  AND2_X1   g510(.A1(new_n437_), .A2(new_n601_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n637_), .A2(new_n568_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT104), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n716_), .A2(KEYINPUT105), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(KEYINPUT105), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n717_), .A2(new_n519_), .A3(new_n374_), .A4(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n568_), .A2(new_n600_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n512_), .A2(new_n619_), .A3(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G57gat), .B1(new_n721_), .B2(new_n623_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n719_), .A2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT106), .ZN(G1332gat));
  OAI21_X1  g523(.A(G64gat), .B1(new_n721_), .B2(new_n644_), .ZN(new_n725_));
  XOR2_X1   g524(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n716_), .A2(new_n521_), .A3(new_n403_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1333gat));
  OAI21_X1  g528(.A(G71gat), .B1(new_n721_), .B2(new_n391_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT109), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n716_), .A2(new_n516_), .A3(new_n436_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1334gat));
  OAI21_X1  g534(.A(G78gat), .B1(new_n721_), .B2(new_n274_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT50), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n716_), .A2(new_n243_), .A3(new_n706_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1335gat));
  AND3_X1   g538(.A1(new_n712_), .A2(new_n569_), .A3(new_n658_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(new_n453_), .A3(new_n374_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n665_), .A2(new_n669_), .A3(new_n743_), .A4(new_n667_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n568_), .A2(new_n619_), .A3(new_n600_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n662_), .B1(new_n437_), .B2(new_n663_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(KEYINPUT98), .B2(new_n664_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n743_), .B1(new_n748_), .B2(new_n667_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n742_), .B1(new_n746_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n670_), .A2(KEYINPUT110), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n751_), .A2(KEYINPUT111), .A3(new_n745_), .A4(new_n744_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n750_), .A2(new_n374_), .A3(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n741_), .B1(new_n753_), .B2(new_n453_), .ZN(G1336gat));
  NAND3_X1  g553(.A1(new_n740_), .A2(new_n454_), .A3(new_n403_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n750_), .A2(new_n403_), .A3(new_n752_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(new_n454_), .ZN(G1337gat));
  NAND3_X1  g556(.A1(new_n750_), .A2(new_n436_), .A3(new_n752_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G99gat), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n740_), .A2(new_n436_), .A3(new_n449_), .A4(new_n451_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT51), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n759_), .A2(new_n763_), .A3(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1338gat));
  NAND3_X1  g564(.A1(new_n740_), .A2(new_n450_), .A3(new_n706_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT112), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n670_), .A2(new_n706_), .A3(new_n745_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(G106gat), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n767_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR4_X1   g573(.A1(new_n706_), .A2(new_n403_), .A3(new_n623_), .A4(new_n391_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n584_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n581_), .A2(new_n585_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n596_), .B1(new_n778_), .B2(new_n590_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n599_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT68), .B1(new_n561_), .B2(new_n554_), .ZN(new_n782_));
  AND4_X1   g581(.A1(KEYINPUT68), .A2(new_n544_), .A3(new_n549_), .A4(new_n554_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n781_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n544_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT114), .B1(new_n560_), .B2(new_n513_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n560_), .A2(KEYINPUT55), .A3(new_n513_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789_));
  INV_X1    g588(.A(new_n513_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n543_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n789_), .B(new_n790_), .C1(new_n791_), .C2(new_n534_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .A4(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n553_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n553_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n784_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT58), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n599_), .A2(new_n780_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n557_), .B2(new_n562_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n553_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT56), .B1(new_n793_), .B2(new_n553_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n802_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT58), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(KEYINPUT115), .A3(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n800_), .A2(new_n663_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n563_), .A2(new_n600_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n801_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n511_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT57), .B(new_n511_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n808_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n620_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n568_), .A2(new_n636_), .A3(new_n619_), .A4(new_n601_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(KEYINPUT113), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(KEYINPUT113), .B2(new_n819_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n819_), .A2(KEYINPUT113), .A3(new_n818_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  AND4_X1   g622(.A1(new_n776_), .A2(new_n817_), .A3(new_n821_), .A4(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n822_), .B1(new_n816_), .B2(new_n620_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n776_), .B1(new_n825_), .B2(new_n821_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n775_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT59), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n821_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n775_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G113gat), .B1(new_n832_), .B2(new_n601_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n827_), .A2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT117), .B(new_n775_), .C1(new_n824_), .C2(new_n826_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n601_), .A2(G113gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n833_), .B1(new_n837_), .B2(new_n838_), .ZN(G1340gat));
  INV_X1    g638(.A(KEYINPUT60), .ZN(new_n840_));
  AOI21_X1  g639(.A(G120gat), .B1(new_n569_), .B2(new_n840_), .ZN(new_n841_));
  XOR2_X1   g640(.A(new_n841_), .B(KEYINPUT118), .Z(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n840_), .B2(G120gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n835_), .A2(new_n836_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n835_), .A2(KEYINPUT119), .A3(new_n836_), .A4(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G120gat), .B1(new_n832_), .B2(new_n568_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT120), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n848_), .A2(new_n852_), .A3(new_n849_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1341gat));
  OAI21_X1  g653(.A(G127gat), .B1(new_n832_), .B2(new_n620_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n620_), .A2(G127gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n837_), .B2(new_n856_), .ZN(G1342gat));
  OAI21_X1  g656(.A(G134gat), .B1(new_n832_), .B2(new_n636_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n511_), .A2(G134gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n837_), .B2(new_n859_), .ZN(G1343gat));
  INV_X1    g659(.A(new_n826_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n825_), .A2(new_n776_), .A3(new_n821_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NOR4_X1   g662(.A1(new_n403_), .A2(new_n274_), .A3(new_n623_), .A4(new_n436_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n601_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT121), .B(G141gat), .Z(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1344gat));
  NOR2_X1   g667(.A1(new_n865_), .A2(new_n568_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT122), .B(G148gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1345gat));
  NOR2_X1   g670(.A1(new_n865_), .A2(new_n620_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT61), .B(G155gat), .Z(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  OAI21_X1  g673(.A(G162gat), .B1(new_n865_), .B2(new_n636_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n511_), .A2(G162gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n865_), .B2(new_n876_), .ZN(G1347gat));
  AND2_X1   g676(.A1(new_n403_), .A2(new_n392_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n878_), .A2(new_n600_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT123), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n879_), .A2(KEYINPUT123), .ZN(new_n881_));
  AND4_X1   g680(.A1(new_n274_), .A2(new_n829_), .A3(new_n880_), .A4(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n299_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n883_), .B2(new_n882_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT62), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n829_), .A2(new_n274_), .A3(new_n878_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(new_n296_), .A3(new_n600_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1348gat));
  AOI21_X1  g688(.A(new_n706_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n890_), .A2(G176gat), .A3(new_n569_), .A4(new_n878_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n887_), .A2(new_n569_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(G176gat), .B2(new_n892_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT125), .ZN(G1349gat));
  NAND3_X1  g693(.A1(new_n890_), .A2(new_n619_), .A3(new_n878_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n620_), .A2(new_n285_), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n895_), .A2(new_n293_), .B1(new_n887_), .B2(new_n896_), .ZN(G1350gat));
  NOR2_X1   g696(.A1(new_n511_), .A2(new_n323_), .ZN(new_n898_));
  XOR2_X1   g697(.A(new_n898_), .B(KEYINPUT126), .Z(new_n899_));
  NAND2_X1  g698(.A1(new_n887_), .A2(new_n899_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n887_), .A2(new_n663_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n286_), .ZN(G1351gat));
  NOR4_X1   g701(.A1(new_n644_), .A2(new_n374_), .A3(new_n274_), .A4(new_n436_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n863_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n600_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n569_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g707(.A1(new_n904_), .A2(new_n619_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  AND2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n910_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n913_), .A2(KEYINPUT127), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(KEYINPUT127), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n912_), .B1(new_n914_), .B2(new_n915_), .ZN(G1354gat));
  INV_X1    g715(.A(new_n904_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G218gat), .B1(new_n917_), .B2(new_n636_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n511_), .A2(G218gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n917_), .B2(new_n919_), .ZN(G1355gat));
endmodule


