//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_, new_n968_;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT37), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G29gat), .B(G36gat), .ZN(new_n204_));
  AND2_X1   g003(.A1(new_n204_), .A2(KEYINPUT74), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(KEYINPUT74), .ZN(new_n206_));
  XOR2_X1   g005(.A(G43gat), .B(G50gat), .Z(new_n207_));
  OR3_X1    g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n207_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT15), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G85gat), .ZN(new_n220_));
  INV_X1    g019(.A(G92gat), .ZN(new_n221_));
  NOR3_X1   g020(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT9), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT10), .B(G99gat), .Z(new_n224_));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225_));
  INV_X1    g024(.A(G106gat), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n225_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n213_), .B(new_n223_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n219_), .A2(KEYINPUT66), .ZN(new_n231_));
  NOR4_X1   g030(.A1(KEYINPUT65), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  NOR2_X1   g032(.A1(KEYINPUT65), .A2(G99gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n233_), .B1(new_n234_), .B2(new_n226_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT66), .B1(new_n215_), .B2(new_n217_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n231_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n230_), .B1(new_n239_), .B2(new_n212_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n236_), .A2(new_n218_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(new_n230_), .A3(new_n212_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n229_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n212_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n237_), .A2(new_n235_), .A3(new_n232_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n248_), .B2(new_n231_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n242_), .B1(new_n249_), .B2(new_n230_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(KEYINPUT70), .A3(new_n229_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n211_), .A2(new_n246_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n244_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT35), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G232gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT34), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n253_), .A2(new_n210_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT75), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n254_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n210_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n260_), .B(new_n261_), .C1(new_n244_), .C2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n257_), .A2(new_n254_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n259_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n264_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(new_n258_), .A3(new_n252_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT77), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G190gat), .B(G218gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G134gat), .B(G162gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n273_), .B(KEYINPUT36), .Z(new_n274_));
  NAND3_X1  g073(.A1(new_n269_), .A2(new_n270_), .A3(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n273_), .A2(KEYINPUT36), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n266_), .A2(new_n268_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n270_), .B1(new_n269_), .B2(new_n274_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n203_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n274_), .B(KEYINPUT76), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n269_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(KEYINPUT37), .A3(new_n277_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G57gat), .B(G64gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G64gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G57gat), .ZN(new_n288_));
  INV_X1    g087(.A(G57gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G64gat), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n288_), .A2(new_n290_), .A3(new_n285_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT11), .B1(new_n286_), .B2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT67), .B(G71gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(G78gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n288_), .A2(new_n290_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT68), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n284_), .A2(new_n285_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT11), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n292_), .A2(new_n294_), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n301_));
  INV_X1    g100(.A(G78gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n293_), .B(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n300_), .A2(new_n304_), .A3(KEYINPUT69), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT69), .B1(new_n300_), .B2(new_n304_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G15gat), .B(G22gat), .ZN(new_n309_));
  INV_X1    g108(.A(G1gat), .ZN(new_n310_));
  INV_X1    g109(.A(G8gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT14), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G1gat), .B(G8gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G231gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT78), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n315_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n308_), .B(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(G127gat), .B(G155gat), .Z(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G183gat), .B(G211gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n324_), .A2(KEYINPUT17), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(KEYINPUT17), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n319_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT80), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n300_), .A2(new_n304_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n318_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n318_), .A2(new_n330_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n325_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n280_), .A2(new_n283_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT69), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n330_), .A2(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n339_), .A2(new_n250_), .A3(new_n229_), .A4(new_n305_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G230gat), .A2(G233gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT72), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(KEYINPUT72), .A3(new_n341_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT12), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n330_), .A2(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n246_), .A2(new_n347_), .A3(new_n251_), .A4(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n244_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n348_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n246_), .A2(new_n251_), .A3(new_n349_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT71), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n346_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(new_n340_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n341_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G120gat), .B(G148gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT5), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G176gat), .B(G204gat), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n356_), .A2(new_n359_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n364_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT73), .ZN(new_n368_));
  OAI22_X1  g167(.A1(new_n366_), .A2(new_n367_), .B1(new_n368_), .B2(KEYINPUT13), .ZN(new_n369_));
  INV_X1    g168(.A(new_n367_), .ZN(new_n370_));
  XOR2_X1   g169(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n365_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n202_), .B1(new_n337_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT23), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(G183gat), .A3(G190gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT23), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT89), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT89), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n382_), .A3(KEYINPUT23), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n378_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G169gat), .A2(G176gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT24), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n387_), .B1(new_n389_), .B2(new_n385_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n384_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT25), .B(G183gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G183gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n395_), .B2(KEYINPUT25), .ZN(new_n396_));
  INV_X1    g195(.A(G190gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT26), .B1(new_n397_), .B2(KEYINPUT88), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT88), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT26), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(G190gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n396_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n394_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n388_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT22), .B(G169gat), .ZN(new_n405_));
  INV_X1    g204(.A(G176gat), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT90), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n380_), .A2(new_n377_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(G183gat), .A2(G190gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n414_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n415_));
  OAI22_X1  g214(.A1(new_n391_), .A2(new_n403_), .B1(new_n410_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G227gat), .A2(G233gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G15gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n416_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT91), .B(KEYINPUT30), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G113gat), .B(G120gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(G134gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G127gat), .ZN(new_n425_));
  INV_X1    g224(.A(G127gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(G134gat), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n425_), .A2(new_n427_), .A3(KEYINPUT92), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT92), .B1(new_n425_), .B2(new_n427_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n423_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT92), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n426_), .A2(G134gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n424_), .A2(G127gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n425_), .A2(new_n427_), .A3(KEYINPUT92), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n422_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n430_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n421_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n421_), .A2(new_n438_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G71gat), .B(G99gat), .Z(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(G43gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT31), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n441_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n439_), .A2(new_n444_), .A3(new_n440_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G226gat), .A2(G233gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT19), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G211gat), .B(G218gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G197gat), .B(G204gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT21), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n452_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT96), .ZN(new_n458_));
  AND2_X1   g257(.A1(G197gat), .A2(G204gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G197gat), .A2(G204gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n458_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n454_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n458_), .B(KEYINPUT21), .C1(new_n459_), .C2(new_n460_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n457_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT97), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  AOI211_X1 g265(.A(KEYINPUT97), .B(new_n457_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n456_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT20), .B1(new_n468_), .B2(new_n416_), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT21), .B1(new_n453_), .B2(new_n458_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n463_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n452_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT97), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n464_), .A2(new_n465_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT100), .B1(new_n384_), .B2(new_n412_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n379_), .A2(new_n382_), .A3(KEYINPUT23), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n382_), .B1(new_n379_), .B2(KEYINPUT23), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n377_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT100), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n413_), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT22), .B(G169gat), .Z(new_n482_));
  INV_X1    g281(.A(KEYINPUT99), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n405_), .A2(KEYINPUT99), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n406_), .A3(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n476_), .A2(new_n388_), .A3(new_n481_), .A4(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(KEYINPUT26), .B(G190gat), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n392_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n385_), .B1(new_n389_), .B2(KEYINPUT98), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n491_), .B1(KEYINPUT98), .B2(new_n389_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n490_), .A2(new_n492_), .A3(new_n411_), .A4(new_n387_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n475_), .A2(new_n456_), .B1(new_n487_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n451_), .B1(new_n469_), .B2(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G8gat), .B(G36gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G64gat), .B(G92gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n468_), .A2(new_n416_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT20), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n451_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n487_), .A2(new_n493_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n501_), .B(new_n503_), .C1(new_n468_), .C2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n495_), .A2(new_n500_), .A3(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n506_), .A2(KEYINPUT27), .ZN(new_n507_));
  XOR2_X1   g306(.A(KEYINPUT106), .B(KEYINPUT20), .Z(new_n508_));
  NAND2_X1  g307(.A1(new_n501_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n504_), .A2(new_n468_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n451_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n455_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n415_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n403_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n384_), .A2(new_n390_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n513_), .A2(new_n409_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n502_), .B1(new_n512_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n451_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n504_), .A2(new_n468_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n511_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n500_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT108), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT108), .ZN(new_n524_));
  AOI211_X1 g323(.A(new_n524_), .B(new_n500_), .C1(new_n511_), .C2(new_n520_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n507_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n518_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n503_), .B1(new_n512_), .B2(new_n516_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(new_n510_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n522_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(KEYINPUT102), .A3(new_n506_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT27), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT102), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n533_), .B(new_n522_), .C1(new_n527_), .C2(new_n529_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n531_), .A2(new_n532_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n526_), .A2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G141gat), .B(G148gat), .Z(new_n537_));
  INV_X1    g336(.A(G155gat), .ZN(new_n538_));
  INV_X1    g337(.A(G162gat), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(KEYINPUT93), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT93), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n541_), .B1(G155gat), .B2(G162gat), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT1), .B1(new_n538_), .B2(new_n539_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT1), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(G155gat), .A3(G162gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n537_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT2), .ZN(new_n549_));
  INV_X1    g348(.A(G141gat), .ZN(new_n550_));
  INV_X1    g349(.A(G148gat), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n549_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT3), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n552_), .A2(new_n554_), .A3(new_n555_), .A4(new_n556_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n540_), .A2(new_n542_), .B1(G155gat), .B2(G162gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n548_), .A2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n512_), .B1(KEYINPUT29), .B2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G22gat), .B(G50gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n548_), .A2(new_n559_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT29), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT28), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT94), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT28), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n567_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT94), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(KEYINPUT95), .A2(G228gat), .ZN(new_n574_));
  NOR2_X1   g373(.A1(KEYINPUT95), .A2(G228gat), .ZN(new_n575_));
  OAI21_X1  g374(.A(G233gat), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(new_n302_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n226_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n569_), .A2(new_n573_), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n564_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n569_), .A2(new_n573_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n578_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n569_), .A2(new_n573_), .A3(new_n579_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n563_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n536_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n560_), .A2(new_n437_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT103), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n548_), .A2(new_n430_), .A3(new_n436_), .A4(new_n559_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n438_), .A2(new_n565_), .A3(KEYINPUT103), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n592_), .A2(new_n593_), .B1(G225gat), .B2(G233gat), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n589_), .A2(KEYINPUT4), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n593_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n595_), .B1(new_n596_), .B2(KEYINPUT4), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G225gat), .A2(G233gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT104), .Z(new_n599_));
  AOI21_X1  g398(.A(new_n594_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G1gat), .B(G29gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(G85gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT0), .B(G57gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  OR3_X1    g404(.A1(new_n600_), .A2(KEYINPUT107), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT4), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n599_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n608_), .A2(new_n609_), .A3(new_n595_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n604_), .B1(new_n610_), .B2(new_n594_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n596_), .A2(KEYINPUT4), .ZN(new_n612_));
  INV_X1    g411(.A(new_n595_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n599_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n594_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(new_n605_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n611_), .A2(new_n616_), .A3(KEYINPUT107), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n606_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n449_), .A2(new_n588_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n587_), .A2(new_n618_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n536_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n531_), .A2(new_n534_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n597_), .A2(new_n598_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n605_), .B1(new_n596_), .B2(new_n599_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n600_), .B2(new_n605_), .ZN(new_n627_));
  NOR4_X1   g426(.A1(new_n610_), .A2(KEYINPUT33), .A3(new_n594_), .A4(new_n604_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n625_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT105), .B1(new_n622_), .B2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n531_), .A2(new_n534_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n616_), .A2(KEYINPUT33), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n600_), .A2(new_n626_), .A3(new_n605_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT105), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n631_), .A2(new_n634_), .A3(new_n635_), .A4(new_n625_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n500_), .A2(KEYINPUT32), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n527_), .A2(new_n529_), .A3(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n521_), .B2(new_n637_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n606_), .A3(new_n617_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n630_), .A2(new_n636_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n587_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n621_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n619_), .B1(new_n643_), .B2(new_n449_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n336_), .A2(KEYINPUT81), .A3(new_n373_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n315_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n210_), .A2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT82), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n211_), .A2(new_n315_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(G229gat), .A2(G233gat), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT84), .Z(new_n652_));
  NAND3_X1  g451(.A1(new_n649_), .A2(new_n650_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n262_), .A2(new_n315_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT83), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n648_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n656_), .B2(new_n651_), .ZN(new_n657_));
  XOR2_X1   g456(.A(G113gat), .B(G141gat), .Z(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT86), .ZN(new_n659_));
  XOR2_X1   g458(.A(G169gat), .B(G197gat), .Z(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(KEYINPUT85), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n657_), .B(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n375_), .A2(new_n644_), .A3(new_n645_), .A4(new_n663_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT109), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(KEYINPUT109), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT38), .ZN(new_n668_));
  INV_X1    g467(.A(new_n618_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n310_), .ZN(new_n670_));
  OR3_X1    g469(.A1(new_n667_), .A2(new_n668_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n269_), .A2(new_n274_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT77), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(new_n277_), .A3(new_n275_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n644_), .A2(new_n335_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n663_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n374_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G1gat), .B1(new_n678_), .B2(new_n618_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n668_), .B1(new_n667_), .B2(new_n670_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n671_), .A2(new_n679_), .A3(new_n680_), .ZN(G1324gat));
  NAND4_X1  g480(.A1(new_n665_), .A2(new_n311_), .A3(new_n536_), .A4(new_n666_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n683_));
  INV_X1    g482(.A(new_n536_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G8gat), .B1(new_n678_), .B2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(KEYINPUT39), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(KEYINPUT39), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n682_), .B(new_n683_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n685_), .B(KEYINPUT39), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n683_), .B1(new_n690_), .B2(new_n682_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1325gat));
  OAI21_X1  g491(.A(G15gat), .B1(new_n678_), .B2(new_n448_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT41), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n667_), .A2(G15gat), .A3(new_n448_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1326gat));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n697_));
  INV_X1    g496(.A(new_n678_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n587_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n699_), .B2(G22gat), .ZN(new_n700_));
  INV_X1    g499(.A(G22gat), .ZN(new_n701_));
  AOI211_X1 g500(.A(KEYINPUT42), .B(new_n701_), .C1(new_n698_), .C2(new_n587_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n587_), .A2(new_n701_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n667_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT111), .B1(new_n703_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n707_));
  OAI221_X1 g506(.A(new_n707_), .B1(new_n667_), .B2(new_n704_), .C1(new_n700_), .C2(new_n702_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1327gat));
  NAND2_X1  g508(.A1(new_n644_), .A2(new_n663_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n674_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n334_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n710_), .A2(new_n374_), .A3(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G29gat), .B1(new_n713_), .B2(new_n669_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n677_), .A2(new_n334_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n717_));
  INV_X1    g516(.A(new_n283_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n674_), .B2(new_n203_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n644_), .A2(new_n717_), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n717_), .B1(new_n644_), .B2(new_n720_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n716_), .B(KEYINPUT44), .C1(new_n721_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n644_), .A2(new_n720_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT43), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n644_), .A2(new_n717_), .A3(new_n720_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n729_), .A2(KEYINPUT112), .A3(KEYINPUT44), .A4(new_n716_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n725_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n716_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n669_), .A2(G29gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n714_), .B1(new_n736_), .B2(new_n737_), .ZN(G1328gat));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739_));
  INV_X1    g538(.A(G36gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n713_), .A2(new_n740_), .A3(new_n536_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT45), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n684_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n740_), .B1(new_n731_), .B2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n739_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n715_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n536_), .B1(new_n747_), .B2(KEYINPUT44), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n725_), .B2(new_n730_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n742_), .B(KEYINPUT46), .C1(new_n749_), .C2(new_n740_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(new_n750_), .ZN(G1329gat));
  NAND2_X1  g550(.A1(new_n449_), .A2(G43gat), .ZN(new_n752_));
  AOI221_X4 g551(.A(new_n752_), .B1(new_n733_), .B2(new_n732_), .C1(new_n725_), .C2(new_n730_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G43gat), .B1(new_n713_), .B2(new_n449_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT47), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n756_));
  INV_X1    g555(.A(new_n754_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n756_), .B(new_n757_), .C1(new_n735_), .C2(new_n752_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(new_n758_), .ZN(G1330gat));
  AOI21_X1  g558(.A(G50gat), .B1(new_n713_), .B2(new_n587_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n587_), .A2(G50gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n736_), .B2(new_n761_), .ZN(G1331gat));
  NOR2_X1   g561(.A1(new_n373_), .A2(new_n663_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n675_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G57gat), .B1(new_n765_), .B2(new_n618_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n644_), .A2(new_n676_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n767_), .A2(new_n374_), .A3(new_n336_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n289_), .A3(new_n669_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n766_), .A2(new_n769_), .ZN(G1332gat));
  AOI21_X1  g569(.A(new_n287_), .B1(new_n764_), .B2(new_n536_), .ZN(new_n771_));
  XOR2_X1   g570(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n768_), .A2(new_n287_), .A3(new_n536_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1333gat));
  INV_X1    g574(.A(G71gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n764_), .B2(new_n449_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT49), .Z(new_n778_));
  NAND3_X1  g577(.A1(new_n768_), .A2(new_n776_), .A3(new_n449_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1334gat));
  AOI21_X1  g579(.A(new_n302_), .B1(new_n764_), .B2(new_n587_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT50), .Z(new_n782_));
  NAND3_X1  g581(.A1(new_n768_), .A2(new_n302_), .A3(new_n587_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1335gat));
  AND4_X1   g583(.A1(new_n374_), .A2(new_n767_), .A3(new_n334_), .A4(new_n711_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n220_), .A3(new_n669_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n373_), .A2(new_n663_), .A3(new_n335_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n729_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n669_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n790_), .B2(new_n220_), .ZN(G1336gat));
  NAND3_X1  g590(.A1(new_n785_), .A2(new_n221_), .A3(new_n536_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n788_), .A2(new_n536_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n792_), .B1(new_n794_), .B2(new_n221_), .ZN(G1337gat));
  NAND2_X1  g594(.A1(new_n788_), .A2(new_n449_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n449_), .A2(new_n224_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n796_), .A2(G99gat), .B1(new_n785_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT51), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n798_), .B(new_n800_), .ZN(G1338gat));
  OAI211_X1 g600(.A(new_n587_), .B(new_n787_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(G106gat), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(KEYINPUT115), .A3(G106gat), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(KEYINPUT52), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT115), .B1(new_n802_), .B2(G106gat), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n642_), .A2(G106gat), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n808_), .A2(new_n809_), .B1(new_n785_), .B2(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n807_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n807_), .B2(new_n811_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1339gat));
  INV_X1    g614(.A(new_n652_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n649_), .A2(new_n650_), .A3(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n656_), .B2(new_n816_), .ZN(new_n818_));
  MUX2_X1   g617(.A(new_n818_), .B(new_n657_), .S(new_n661_), .Z(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n365_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n355_), .A2(new_n352_), .A3(new_n350_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n345_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT72), .B1(new_n340_), .B2(new_n341_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n821_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n346_), .A2(new_n353_), .A3(KEYINPUT55), .A4(new_n355_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n355_), .A2(new_n340_), .A3(new_n352_), .A4(new_n350_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n358_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n826_), .A2(new_n827_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n363_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n363_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n820_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT58), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n363_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT56), .B1(new_n830_), .B2(new_n363_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT118), .B(new_n838_), .C1(new_n841_), .C2(new_n820_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n837_), .A2(new_n842_), .A3(new_n720_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n663_), .A2(new_n365_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n370_), .A2(new_n365_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n819_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT57), .B(new_n674_), .C1(new_n845_), .C2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT119), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n674_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n847_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(KEYINPUT57), .A4(new_n674_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n843_), .A2(new_n850_), .A3(new_n853_), .A4(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n334_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n719_), .A2(new_n373_), .A3(new_n676_), .A4(new_n335_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n336_), .A2(KEYINPUT117), .A3(new_n676_), .A4(new_n373_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(KEYINPUT54), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n859_), .A2(new_n860_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n858_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n449_), .A2(new_n588_), .A3(new_n669_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n868_), .B(new_n870_), .C1(KEYINPUT120), .C2(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n866_), .B1(new_n857_), .B2(new_n334_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n869_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n872_), .A2(new_n663_), .A3(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G113gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n875_), .A2(new_n869_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  OR3_X1    g679(.A1(new_n880_), .A2(G113gat), .A3(new_n676_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n881_), .ZN(G1340gat));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n373_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n879_), .B(new_n884_), .C1(KEYINPUT60), .C2(new_n883_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n872_), .A2(new_n374_), .A3(new_n876_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n883_), .ZN(G1341gat));
  OAI21_X1  g686(.A(new_n426_), .B1(new_n880_), .B2(new_n334_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n426_), .B1(new_n335_), .B2(KEYINPUT121), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(KEYINPUT121), .B2(new_n426_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n872_), .A2(new_n876_), .A3(new_n890_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n888_), .A2(new_n891_), .ZN(G1342gat));
  OAI21_X1  g691(.A(new_n424_), .B1(new_n880_), .B2(new_n674_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n720_), .A2(G134gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT122), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n872_), .A2(new_n876_), .A3(new_n895_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n893_), .A2(new_n896_), .ZN(G1343gat));
  NOR4_X1   g696(.A1(new_n449_), .A2(new_n536_), .A3(new_n618_), .A4(new_n642_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n868_), .A2(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT124), .B1(new_n899_), .B2(new_n676_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n898_), .ZN(new_n901_));
  NOR4_X1   g700(.A1(new_n875_), .A2(KEYINPUT124), .A3(new_n676_), .A4(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT123), .B(G141gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n900_), .A2(new_n903_), .A3(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n904_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n875_), .A2(new_n901_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n663_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n906_), .B1(new_n909_), .B2(new_n902_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n905_), .A2(new_n910_), .ZN(G1344gat));
  NAND2_X1  g710(.A1(new_n908_), .A2(new_n374_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g712(.A1(new_n908_), .A2(new_n335_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT61), .B(G155gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1346gat));
  OAI21_X1  g715(.A(G162gat), .B1(new_n899_), .B2(new_n719_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n908_), .A2(new_n539_), .A3(new_n711_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1347gat));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  NOR4_X1   g719(.A1(new_n448_), .A2(new_n684_), .A3(new_n669_), .A4(new_n587_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n868_), .A2(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n676_), .ZN(new_n923_));
  INV_X1    g722(.A(G169gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n920_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n926_));
  OAI211_X1 g725(.A(KEYINPUT62), .B(G169gat), .C1(new_n922_), .C2(new_n676_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n925_), .A2(new_n926_), .A3(new_n927_), .ZN(G1348gat));
  NOR2_X1   g727(.A1(new_n922_), .A2(new_n373_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(new_n406_), .ZN(G1349gat));
  INV_X1    g729(.A(new_n392_), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n868_), .A2(new_n931_), .A3(new_n335_), .A4(new_n921_), .ZN(new_n932_));
  OR2_X1    g731(.A1(new_n932_), .A2(KEYINPUT125), .ZN(new_n933_));
  INV_X1    g732(.A(new_n922_), .ZN(new_n934_));
  AOI21_X1  g733(.A(G183gat), .B1(new_n934_), .B2(new_n335_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n932_), .A2(KEYINPUT125), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n933_), .B1(new_n935_), .B2(new_n936_), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n922_), .B2(new_n719_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n711_), .A2(new_n489_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n922_), .B2(new_n939_), .ZN(G1351gat));
  NOR3_X1   g739(.A1(new_n449_), .A2(new_n620_), .A3(new_n684_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n868_), .A2(KEYINPUT126), .A3(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943_));
  INV_X1    g742(.A(new_n941_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n875_), .B2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n942_), .A2(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(G197gat), .B1(new_n946_), .B2(new_n663_), .ZN(new_n947_));
  INV_X1    g746(.A(G197gat), .ZN(new_n948_));
  AOI211_X1 g747(.A(new_n948_), .B(new_n676_), .C1(new_n942_), .C2(new_n945_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n947_), .A2(new_n949_), .ZN(G1352gat));
  AOI21_X1  g749(.A(KEYINPUT126), .B1(new_n868_), .B2(new_n941_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n875_), .A2(new_n943_), .A3(new_n944_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n374_), .B1(new_n951_), .B2(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(G204gat), .ZN(new_n954_));
  INV_X1    g753(.A(G204gat), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n946_), .A2(new_n955_), .A3(new_n374_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n954_), .A2(new_n956_), .ZN(G1353gat));
  AOI21_X1  g756(.A(new_n334_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n958_), .B1(new_n951_), .B2(new_n952_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(KEYINPUT127), .ZN(new_n961_));
  INV_X1    g760(.A(new_n961_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n959_), .A2(new_n962_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n946_), .A2(new_n958_), .A3(new_n961_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n963_), .A2(new_n964_), .ZN(G1354gat));
  INV_X1    g764(.A(G218gat), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n946_), .A2(new_n966_), .A3(new_n711_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n719_), .B1(new_n942_), .B2(new_n945_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n967_), .B1(new_n966_), .B2(new_n968_), .ZN(G1355gat));
endmodule


