//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n789_, new_n790_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT80), .ZN(new_n204_));
  INV_X1    g003(.A(G155gat), .ZN(new_n205_));
  INV_X1    g004(.A(G162gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT80), .B1(G155gat), .B2(G162gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n203_), .A2(new_n207_), .A3(new_n208_), .A4(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n207_), .A2(new_n208_), .A3(new_n202_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT81), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n214_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n219_), .A2(new_n221_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n216_), .A2(new_n217_), .A3(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n217_), .B1(new_n216_), .B2(new_n224_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n215_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT29), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT21), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G197gat), .B(G204gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(G211gat), .A2(G218gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT21), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G211gat), .A2(G218gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n230_), .A2(new_n232_), .A3(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n229_), .A2(new_n231_), .A3(KEYINPUT21), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n228_), .A2(KEYINPUT83), .A3(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT82), .Z(new_n241_));
  AND2_X1   g040(.A1(G228gat), .A2(G233gat), .ZN(new_n242_));
  OR3_X1    g041(.A1(new_n227_), .A2(KEYINPUT29), .A3(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n242_), .B1(new_n227_), .B2(KEYINPUT29), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G22gat), .B(G50gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n247_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n241_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G78gat), .B(G106gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT28), .ZN(new_n253_));
  INV_X1    g052(.A(new_n248_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n240_), .B(KEYINPUT82), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n249_), .A3(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n251_), .A2(new_n253_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n253_), .B1(new_n251_), .B2(new_n256_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT92), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G127gat), .A2(G134gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G127gat), .A2(G134gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(G113gat), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G127gat), .ZN(new_n265_));
  INV_X1    g064(.A(G134gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G113gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n261_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n264_), .A2(new_n269_), .A3(G120gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(G120gat), .B1(new_n264_), .B2(new_n269_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n227_), .A2(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n272_), .B(new_n215_), .C1(new_n226_), .C2(new_n225_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n274_), .A2(KEYINPUT4), .A3(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(KEYINPUT91), .B(KEYINPUT4), .Z(new_n277_));
  NAND3_X1  g076(.A1(new_n227_), .A2(new_n273_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G225gat), .A2(G233gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n260_), .B1(new_n276_), .B2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n274_), .A2(new_n275_), .A3(new_n279_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n274_), .A2(KEYINPUT4), .A3(new_n275_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n284_), .A2(KEYINPUT92), .A3(new_n280_), .A4(new_n278_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT0), .B(G57gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(G85gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(G1gat), .B(G29gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n282_), .A2(new_n283_), .A3(new_n285_), .A4(new_n290_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G15gat), .B(G43gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT79), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n272_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G227gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT30), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT31), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n297_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT23), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(G183gat), .A3(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G183gat), .ZN(new_n307_));
  INV_X1    g106(.A(G190gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G176gat), .ZN(new_n311_));
  AND2_X1   g110(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT78), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n310_), .A2(new_n314_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G169gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n311_), .ZN(new_n322_));
  AND3_X1   g121(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n324_));
  OAI211_X1 g123(.A(KEYINPUT24), .B(new_n322_), .C1(new_n323_), .C2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n326_));
  AND2_X1   g125(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n329_));
  OAI22_X1  g128(.A1(new_n326_), .A2(new_n327_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  OR3_X1    g129(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n325_), .A2(new_n330_), .A3(new_n306_), .A4(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n320_), .A2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G71gat), .B(G99gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n301_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n301_), .A2(new_n335_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n259_), .A2(new_n294_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n340_), .B(KEYINPUT84), .Z(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT19), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n333_), .A2(new_n239_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT20), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n330_), .A2(new_n306_), .A3(new_n331_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n322_), .A2(KEYINPUT24), .A3(new_n315_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT86), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n314_), .A2(new_n319_), .A3(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n349_), .B1(new_n314_), .B2(new_n319_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n310_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT87), .ZN(new_n353_));
  OR2_X1    g152(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n355_));
  AOI21_X1  g154(.A(G176gat), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n323_), .A2(new_n324_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT86), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n314_), .A2(new_n319_), .A3(new_n349_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT87), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n310_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n348_), .B1(new_n353_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n239_), .ZN(new_n364_));
  AOI211_X1 g163(.A(new_n343_), .B(new_n345_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT88), .ZN(new_n367_));
  INV_X1    g166(.A(new_n348_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n361_), .B1(new_n360_), .B2(new_n310_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n303_), .A2(new_n305_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n370_));
  AOI211_X1 g169(.A(KEYINPUT87), .B(new_n370_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n368_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n239_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n320_), .A2(new_n332_), .A3(new_n238_), .A4(new_n237_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n374_), .A2(KEYINPUT85), .A3(KEYINPUT20), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT85), .B1(new_n374_), .B2(KEYINPUT20), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  AOI211_X1 g176(.A(new_n367_), .B(new_n342_), .C1(new_n373_), .C2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT20), .B1(new_n333_), .B2(new_n239_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT85), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n374_), .A2(KEYINPUT85), .A3(KEYINPUT20), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n381_), .B(new_n382_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT88), .B1(new_n383_), .B2(new_n343_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n366_), .B1(new_n378_), .B2(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G8gat), .B(G36gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(G64gat), .B(G92gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n388_), .B(new_n389_), .Z(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n385_), .A2(new_n391_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n390_), .B(new_n366_), .C1(new_n378_), .C2(new_n384_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(KEYINPUT90), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT27), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT90), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n385_), .A2(new_n396_), .A3(new_n391_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n394_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n368_), .A2(new_n364_), .A3(new_n352_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n343_), .B1(new_n399_), .B2(new_n345_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n383_), .B2(new_n343_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n391_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n393_), .A2(KEYINPUT27), .A3(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n339_), .A2(new_n398_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT97), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n398_), .A2(new_n403_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(KEYINPUT97), .A3(new_n339_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n257_), .A2(new_n258_), .A3(new_n294_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n407_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n401_), .A2(KEYINPUT32), .A3(new_n390_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n390_), .A2(KEYINPUT32), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n294_), .B(new_n414_), .C1(new_n385_), .C2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT96), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n274_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n275_), .ZN(new_n421_));
  OR3_X1    g220(.A1(new_n420_), .A2(new_n421_), .A3(KEYINPUT94), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT94), .B1(new_n420_), .B2(new_n421_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n279_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n284_), .A2(new_n279_), .A3(new_n278_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n424_), .A2(new_n425_), .A3(new_n290_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n293_), .A2(KEYINPUT93), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n293_), .A2(KEYINPUT93), .A3(KEYINPUT33), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n426_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n393_), .A2(KEYINPUT90), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n353_), .A2(new_n362_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n364_), .B1(new_n433_), .B2(new_n368_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n381_), .A2(new_n382_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n343_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n367_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n383_), .A2(KEYINPUT88), .A3(new_n343_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n390_), .B1(new_n439_), .B2(new_n366_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n432_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n397_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n431_), .B(KEYINPUT95), .C1(new_n441_), .C2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n394_), .A2(new_n397_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT95), .B1(new_n445_), .B2(new_n431_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n419_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n259_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n413_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n338_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n410_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(G99gat), .A2(G106gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT7), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT8), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(KEYINPUT10), .B(G99gat), .Z(new_n457_));
  INV_X1    g256(.A(G106gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n459_), .B(KEYINPUT65), .Z(new_n460_));
  INV_X1    g259(.A(KEYINPUT66), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(G92gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(KEYINPUT9), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n461_), .A2(G92gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(G85gat), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT9), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G85gat), .B(G92gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n465_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n456_), .B1(new_n460_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G99gat), .A2(G106gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT67), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT6), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n467_), .A2(new_n455_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n470_), .B(KEYINPUT69), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT68), .B(KEYINPUT6), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n467_), .B1(new_n477_), .B2(new_n454_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT8), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n473_), .A2(new_n474_), .A3(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G57gat), .B(G64gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT70), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT11), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G71gat), .B(G78gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  OR3_X1    g284(.A1(new_n482_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n482_), .B(new_n483_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n486_), .B1(new_n487_), .B2(new_n484_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n480_), .A2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(KEYINPUT71), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT12), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G230gat), .A2(G233gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT64), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n480_), .A2(new_n488_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n493_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n494_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n496_), .B1(new_n497_), .B2(new_n489_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G120gat), .B(G148gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(G204gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT5), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(new_n311_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n495_), .A2(new_n498_), .A3(new_n503_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n507_), .B(KEYINPUT13), .Z(new_n508_));
  XNOR2_X1  g307(.A(G29gat), .B(G36gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(G43gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(G50gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT15), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513_));
  INV_X1    g312(.A(G1gat), .ZN(new_n514_));
  INV_X1    g313(.A(G8gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT14), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G1gat), .B(G8gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n517_), .B(new_n518_), .Z(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n512_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n511_), .A2(new_n519_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n511_), .B(new_n519_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(G229gat), .A3(G233gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G113gat), .B(G141gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(new_n321_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(G197gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n528_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT77), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n452_), .A2(new_n508_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n480_), .A2(new_n511_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G232gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT34), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n538_), .A2(KEYINPUT35), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n473_), .A2(new_n474_), .A3(new_n479_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n512_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n536_), .A2(KEYINPUT73), .A3(new_n539_), .A4(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n538_), .A2(KEYINPUT35), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G190gat), .B(G218gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(G134gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(new_n206_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT36), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n548_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n544_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT74), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n550_), .B(KEYINPUT72), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n544_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT74), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n544_), .A2(new_n555_), .A3(new_n549_), .A4(new_n550_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT75), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n557_), .A2(new_n558_), .A3(KEYINPUT37), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n558_), .B1(new_n557_), .B2(KEYINPUT37), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n554_), .A2(new_n551_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(KEYINPUT37), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n559_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n519_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n488_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT16), .B(G183gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(G211gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(G127gat), .B(G155gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT17), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n566_), .B2(KEYINPUT76), .ZN(new_n573_));
  MUX2_X1   g372(.A(new_n572_), .B(KEYINPUT17), .S(new_n573_), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n563_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n535_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT98), .Z(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(new_n514_), .A3(new_n294_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT38), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n575_), .B1(new_n554_), .B2(new_n551_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n535_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n294_), .ZN(new_n583_));
  OAI21_X1  g382(.A(G1gat), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(G1324gat));
  OAI21_X1  g384(.A(G8gat), .B1(new_n582_), .B2(new_n408_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT39), .Z(new_n587_));
  NOR2_X1   g386(.A1(new_n408_), .A2(G8gat), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n587_), .B1(new_n578_), .B2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g389(.A(G15gat), .B1(new_n582_), .B2(new_n338_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT99), .Z(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT41), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n338_), .A2(G15gat), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n593_), .B1(new_n577_), .B2(new_n594_), .ZN(G1326gat));
  OAI21_X1  g394(.A(G22gat), .B1(new_n582_), .B2(new_n448_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT100), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT42), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n535_), .A2(new_n259_), .A3(new_n576_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n598_), .B1(G22gat), .B2(new_n599_), .ZN(G1327gat));
  NOR2_X1   g399(.A1(new_n561_), .A2(new_n574_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT105), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n535_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(G29gat), .B1(new_n604_), .B2(new_n294_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT104), .ZN(new_n606_));
  INV_X1    g405(.A(new_n508_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(new_n575_), .A3(new_n533_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT102), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n451_), .A2(new_n609_), .ZN(new_n610_));
  OAI211_X1 g409(.A(KEYINPUT102), .B(new_n410_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(new_n563_), .A3(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT103), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n612_), .A2(KEYINPUT103), .A3(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n563_), .ZN(new_n619_));
  OR3_X1    g418(.A1(new_n619_), .A2(new_n452_), .A3(KEYINPUT43), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n608_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n606_), .B1(new_n621_), .B2(KEYINPUT44), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n612_), .A2(KEYINPUT103), .A3(new_n613_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT103), .B1(new_n612_), .B2(new_n613_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n620_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n608_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT44), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(KEYINPUT104), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n622_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n625_), .A2(KEYINPUT44), .A3(new_n626_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n630_), .A2(new_n294_), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n605_), .B1(new_n632_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g432(.A(G36gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n604_), .A2(new_n634_), .A3(new_n407_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT45), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n407_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n622_), .B2(new_n629_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT106), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n634_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n408_), .B1(new_n621_), .B2(KEYINPUT44), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT104), .B1(new_n627_), .B2(new_n628_), .ZN(new_n642_));
  AOI211_X1 g441(.A(new_n606_), .B(KEYINPUT44), .C1(new_n625_), .C2(new_n626_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n641_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT106), .B1(new_n644_), .B2(G36gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n636_), .B1(new_n640_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n647_), .B(new_n636_), .C1(new_n640_), .C2(new_n645_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1329gat));
  NAND4_X1  g450(.A1(new_n630_), .A2(G43gat), .A3(new_n450_), .A4(new_n631_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n603_), .A2(new_n338_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(G43gat), .B2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g454(.A1(new_n630_), .A2(new_n259_), .A3(new_n631_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G50gat), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n448_), .A2(G50gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT108), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n657_), .B1(new_n603_), .B2(new_n659_), .ZN(G1331gat));
  NAND2_X1  g459(.A1(new_n508_), .A2(new_n534_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(new_n452_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n576_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT109), .ZN(new_n664_));
  AOI21_X1  g463(.A(G57gat), .B1(new_n664_), .B2(new_n294_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n581_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT110), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(new_n583_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n665_), .B1(new_n669_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g469(.A(G64gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n667_), .B2(new_n407_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT48), .Z(new_n673_));
  NAND3_X1  g472(.A1(new_n664_), .A2(new_n671_), .A3(new_n407_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1333gat));
  NAND2_X1  g474(.A1(new_n667_), .A2(new_n450_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT111), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(new_n677_), .A3(G71gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT49), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n677_), .B1(new_n676_), .B2(G71gat), .ZN(new_n681_));
  OR3_X1    g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n680_), .B1(new_n679_), .B2(new_n681_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n664_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n338_), .A2(G71gat), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT112), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n682_), .B(new_n683_), .C1(new_n684_), .C2(new_n686_), .ZN(G1334gat));
  OAI21_X1  g486(.A(G78gat), .B1(new_n668_), .B2(new_n448_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT50), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n448_), .A2(G78gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n684_), .B2(new_n690_), .ZN(G1335gat));
  OR2_X1    g490(.A1(new_n625_), .A2(KEYINPUT113), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n661_), .A2(new_n574_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n625_), .A2(KEYINPUT113), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G85gat), .B1(new_n695_), .B2(new_n583_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n662_), .A2(new_n602_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n697_), .A2(G85gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n583_), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT114), .ZN(G1336gat));
  INV_X1    g499(.A(new_n697_), .ZN(new_n701_));
  AOI21_X1  g500(.A(G92gat), .B1(new_n701_), .B2(new_n407_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n695_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n464_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n408_), .B1(new_n704_), .B2(new_n462_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n702_), .B1(new_n703_), .B2(new_n705_), .ZN(G1337gat));
  OAI21_X1  g505(.A(G99gat), .B1(new_n695_), .B2(new_n338_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n701_), .A2(new_n457_), .A3(new_n450_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g509(.A1(new_n625_), .A2(new_n259_), .A3(new_n693_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G106gat), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT52), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n697_), .A2(G106gat), .A3(new_n448_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT115), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g516(.A1(new_n259_), .A2(new_n338_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n407_), .A2(new_n583_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n533_), .A2(new_n506_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT55), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n491_), .A2(new_n494_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n496_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n495_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n722_), .A2(new_n721_), .A3(new_n496_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n504_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT56), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT56), .B(new_n504_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n720_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n531_), .B1(new_n526_), .B2(new_n524_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT116), .Z(new_n733_));
  INV_X1    g532(.A(new_n523_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n524_), .B2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n525_), .A2(new_n527_), .A3(new_n531_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n561_), .B1(new_n731_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT57), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT117), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n739_), .B(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n729_), .A2(new_n730_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n743_), .A2(new_n736_), .A3(new_n506_), .A4(new_n735_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT58), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n745_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n563_), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n574_), .B1(new_n742_), .B2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n576_), .A2(new_n607_), .A3(new_n534_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT54), .Z(new_n751_));
  OAI211_X1 g550(.A(new_n718_), .B(new_n719_), .C1(new_n749_), .C2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G113gat), .B1(new_n753_), .B2(new_n533_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n742_), .A2(new_n748_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n575_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n751_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n758_), .A2(KEYINPUT59), .A3(new_n718_), .A4(new_n719_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT59), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n752_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n534_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n754_), .B1(new_n762_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g562(.A(G120gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n764_), .B1(new_n607_), .B2(KEYINPUT60), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n753_), .B(new_n765_), .C1(KEYINPUT60), .C2(new_n764_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n607_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(new_n764_), .ZN(G1341gat));
  NAND3_X1  g567(.A1(new_n753_), .A2(new_n265_), .A3(new_n574_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n575_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(new_n265_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT118), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT118), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(new_n769_), .C1(new_n770_), .C2(new_n265_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1342gat));
  OAI21_X1  g574(.A(new_n266_), .B1(new_n752_), .B2(new_n561_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT119), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n776_), .A2(new_n777_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n619_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n778_), .B(new_n779_), .C1(G134gat), .C2(new_n780_), .ZN(G1343gat));
  NAND3_X1  g580(.A1(new_n719_), .A2(new_n259_), .A3(new_n338_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT120), .Z(new_n783_));
  NAND2_X1  g582(.A1(new_n758_), .A2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n784_), .A2(new_n534_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(new_n211_), .ZN(G1344gat));
  NOR2_X1   g585(.A1(new_n784_), .A2(new_n607_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(new_n212_), .ZN(G1345gat));
  NOR2_X1   g587(.A1(new_n784_), .A2(new_n575_), .ZN(new_n789_));
  XOR2_X1   g588(.A(KEYINPUT61), .B(G155gat), .Z(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(G1346gat));
  NOR3_X1   g590(.A1(new_n784_), .A2(new_n206_), .A3(new_n619_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n784_), .A2(new_n561_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n206_), .B2(new_n793_), .ZN(G1347gat));
  AOI21_X1  g593(.A(new_n408_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n339_), .ZN(new_n796_));
  OAI21_X1  g595(.A(G169gat), .B1(new_n796_), .B2(new_n534_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(KEYINPUT62), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(KEYINPUT62), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n533_), .B1(new_n313_), .B2(new_n312_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT121), .ZN(new_n801_));
  OAI22_X1  g600(.A1(new_n798_), .A2(new_n799_), .B1(new_n796_), .B2(new_n801_), .ZN(G1348gat));
  NOR2_X1   g601(.A1(new_n796_), .A2(new_n607_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(new_n311_), .ZN(G1349gat));
  NOR2_X1   g603(.A1(new_n327_), .A2(new_n326_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n795_), .A2(new_n574_), .A3(new_n805_), .A4(new_n339_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n806_), .A2(KEYINPUT122), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n307_), .B1(new_n796_), .B2(new_n575_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(KEYINPUT122), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(G1350gat));
  OAI21_X1  g609(.A(G190gat), .B1(new_n796_), .B2(new_n619_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n554_), .B(new_n551_), .C1(new_n329_), .C2(new_n328_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n796_), .B2(new_n812_), .ZN(G1351gat));
  NOR2_X1   g612(.A1(new_n412_), .A2(new_n450_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n795_), .A2(KEYINPUT123), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT123), .B1(new_n795_), .B2(new_n814_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n533_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g618(.A1(new_n795_), .A2(new_n814_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT123), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n607_), .B1(new_n822_), .B2(new_n815_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT124), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(G204gat), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n824_), .A2(G204gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n823_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n823_), .B2(new_n825_), .ZN(G1353gat));
  INV_X1    g627(.A(KEYINPUT63), .ZN(new_n829_));
  INV_X1    g628(.A(G211gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n574_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT125), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n822_), .B2(new_n815_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT126), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n829_), .A2(new_n830_), .A3(KEYINPUT126), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n835_), .B2(new_n833_), .ZN(G1354gat));
  OAI211_X1 g637(.A(G218gat), .B(new_n563_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n561_), .B1(new_n822_), .B2(new_n815_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(G218gat), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(G1355gat));
endmodule


