//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n947_, new_n948_, new_n950_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n983_, new_n984_, new_n985_,
    new_n987_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n995_, new_n996_;
  INV_X1    g000(.A(KEYINPUT12), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G71gat), .B(G78gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT11), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n206_));
  INV_X1    g005(.A(new_n204_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n205_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT6), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT10), .B(G99gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n214_), .B1(G106gat), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT64), .B(G85gat), .ZN(new_n219_));
  INV_X1    g018(.A(G92gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n216_), .B1(new_n217_), .B2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G85gat), .B(G92gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT66), .ZN(new_n224_));
  OR4_X1    g023(.A1(KEYINPUT65), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n225_));
  OAI22_X1  g024(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n214_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT8), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n224_), .A2(new_n230_), .A3(new_n227_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n222_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n202_), .B1(new_n212_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G230gat), .A2(G233gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n229_), .A2(new_n231_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n210_), .A2(KEYINPUT67), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n210_), .A2(KEYINPUT67), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n221_), .A2(new_n217_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n238_), .B(new_n214_), .C1(G106gat), .C2(new_n215_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .A4(new_n239_), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n224_), .A2(new_n230_), .A3(new_n227_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n230_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n239_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  OAI211_X1 g042(.A(KEYINPUT12), .B(new_n205_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n233_), .A2(new_n234_), .A3(new_n240_), .A4(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n210_), .B(KEYINPUT67), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(new_n243_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n244_), .B1(new_n235_), .B2(new_n239_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n253_), .A2(KEYINPUT68), .A3(new_n234_), .A4(new_n233_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n234_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n212_), .A2(new_n232_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n255_), .B1(new_n256_), .B2(new_n251_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n249_), .A2(new_n254_), .A3(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G120gat), .B(G148gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT5), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G176gat), .B(G204gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(new_n261_), .Z(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n262_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n249_), .A2(new_n254_), .A3(new_n257_), .A4(new_n264_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n263_), .A2(KEYINPUT13), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT13), .B1(new_n263_), .B2(new_n265_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT69), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G232gat), .A2(G233gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n274_), .B(KEYINPUT34), .Z(new_n275_));
  INV_X1    g074(.A(KEYINPUT35), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n277_), .B(KEYINPUT71), .Z(new_n278_));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n275_), .A2(new_n276_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G29gat), .B(G36gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G43gat), .B(G50gat), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n283_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT70), .B(KEYINPUT15), .Z(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n243_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n286_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n281_), .B(new_n289_), .C1(new_n290_), .C2(new_n243_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n280_), .A2(new_n279_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n292_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT36), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G190gat), .B(G218gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT72), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G134gat), .B(G162gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n298_), .B(new_n299_), .Z(new_n300_));
  NAND3_X1  g099(.A1(new_n295_), .A2(new_n296_), .A3(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(KEYINPUT36), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n293_), .A2(new_n294_), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT37), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT37), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(new_n306_), .A3(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G15gat), .B(G22gat), .ZN(new_n310_));
  INV_X1    g109(.A(G1gat), .ZN(new_n311_));
  INV_X1    g110(.A(G8gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT14), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G1gat), .B(G8gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G231gat), .A2(G233gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  XOR2_X1   g117(.A(new_n318_), .B(KEYINPUT76), .Z(new_n319_));
  OR2_X1    g118(.A1(new_n319_), .A2(new_n250_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n250_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G127gat), .B(G155gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G183gat), .B(G211gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT17), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT77), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n320_), .A2(new_n321_), .A3(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n210_), .B(KEYINPUT74), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n331_), .A2(new_n318_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT17), .ZN(new_n333_));
  NOR3_X1   g132(.A1(new_n332_), .A2(new_n333_), .A3(new_n326_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(new_n318_), .B2(new_n331_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n329_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n309_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n273_), .A2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n338_), .B(KEYINPUT78), .Z(new_n339_));
  INV_X1    g138(.A(KEYINPUT27), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT20), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(G183gat), .A3(G190gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n344_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT81), .B1(new_n344_), .B2(KEYINPUT23), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n343_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G183gat), .A2(G190gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT22), .B(G169gat), .ZN(new_n353_));
  INV_X1    g152(.A(G176gat), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n352_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(G169gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n354_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n357_), .A2(KEYINPUT24), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(KEYINPUT24), .A3(new_n351_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G183gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT25), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(G183gat), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT26), .B(G190gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n344_), .A2(KEYINPUT23), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n365_), .A2(new_n366_), .B1(new_n343_), .B2(new_n367_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n350_), .A2(new_n355_), .B1(new_n360_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G204gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(G197gat), .ZN(new_n371_));
  INV_X1    g170(.A(G197gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(G204gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT21), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G211gat), .B(G218gat), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT89), .B1(new_n372_), .B2(G204gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT89), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n370_), .A3(G197gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n380_), .A3(new_n373_), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n381_), .A2(KEYINPUT21), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT21), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n376_), .A2(new_n383_), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n377_), .A2(new_n382_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n341_), .B1(new_n369_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT19), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n367_), .A2(new_n343_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n349_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n392_));
  AOI21_X1  g191(.A(G176gat), .B1(new_n392_), .B2(KEYINPUT22), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n393_), .A2(new_n356_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n356_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n347_), .A2(new_n358_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n399_));
  INV_X1    g198(.A(G190gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT26), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT26), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G190gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n363_), .A2(G183gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n401_), .B(new_n403_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT79), .B1(new_n362_), .B2(new_n364_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n359_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n398_), .B1(new_n399_), .B2(new_n408_), .ZN(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT80), .B(new_n359_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n397_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n386_), .B(new_n389_), .C1(new_n411_), .C2(new_n385_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT91), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n408_), .A2(new_n399_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n347_), .A2(new_n358_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n410_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n385_), .B1(new_n417_), .B2(new_n396_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n419_), .A2(KEYINPUT91), .A3(new_n389_), .A4(new_n386_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n417_), .A2(new_n385_), .A3(new_n396_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n343_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT81), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n367_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n344_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n428_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n355_), .B1(new_n432_), .B2(new_n348_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n365_), .A2(new_n366_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n434_), .A2(new_n359_), .A3(new_n358_), .A4(new_n390_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n384_), .A2(new_n381_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n375_), .A2(new_n376_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n381_), .A2(KEYINPUT21), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n341_), .B1(new_n436_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n427_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n388_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n414_), .A2(new_n420_), .A3(new_n426_), .A4(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n389_), .B1(new_n427_), .B2(new_n441_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n426_), .B1(new_n447_), .B2(new_n420_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n340_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT102), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT20), .B1(new_n436_), .B2(new_n440_), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n418_), .A2(new_n452_), .A3(new_n388_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n443_), .B1(new_n453_), .B2(KEYINPUT91), .ZN(new_n454_));
  INV_X1    g253(.A(new_n420_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n425_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n444_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(KEYINPUT102), .A3(new_n340_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n427_), .A2(new_n441_), .A3(new_n389_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT98), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n427_), .A2(new_n441_), .A3(KEYINPUT98), .A4(new_n389_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n388_), .B1(new_n418_), .B2(new_n452_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n425_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(KEYINPUT27), .A3(new_n444_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT101), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT101), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n465_), .A2(new_n468_), .A3(new_n444_), .A4(KEYINPUT27), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n451_), .A2(new_n458_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT100), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G1gat), .B(G29gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G57gat), .B(G85gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G134gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(G127gat), .ZN(new_n479_));
  INV_X1    g278(.A(G127gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(G134gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G120gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G113gat), .ZN(new_n484_));
  INV_X1    g283(.A(G113gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(G120gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n482_), .A2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n479_), .A2(new_n481_), .A3(new_n484_), .A4(new_n486_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT93), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n490_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G141gat), .A2(G148gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT85), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(G141gat), .A2(G148gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G155gat), .A2(G162gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT86), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(G155gat), .A3(G162gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT1), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(G155gat), .A2(G162gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n505_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n506_), .B(new_n507_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n510_));
  AOI211_X1 g309(.A(KEYINPUT87), .B(new_n505_), .C1(new_n502_), .C2(new_n504_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n500_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT88), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n499_), .B(KEYINPUT3), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n514_), .B(new_n515_), .C1(KEYINPUT2), .C2(new_n498_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n502_), .A2(new_n504_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n507_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n493_), .A2(new_n512_), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n492_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n512_), .B2(new_n520_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT4), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G225gat), .A2(G233gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n512_), .A2(new_n520_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n488_), .A2(new_n489_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT94), .B(KEYINPUT4), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n524_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n525_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n477_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT4), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n527_), .A2(new_n492_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n493_), .A2(new_n512_), .A3(new_n520_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n517_), .A2(KEYINPUT1), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT87), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n506_), .A2(new_n507_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n508_), .A2(new_n509_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n543_), .A2(new_n500_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n529_), .A2(new_n530_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n526_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n533_), .B(new_n477_), .C1(new_n538_), .C2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n471_), .B1(new_n534_), .B2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n538_), .A2(new_n546_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n533_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n476_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(KEYINPUT100), .A3(new_n547_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G71gat), .B(G99gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(G43gat), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n417_), .B2(new_n396_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n411_), .A2(new_n557_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G227gat), .A2(G233gat), .ZN(new_n561_));
  INV_X1    g360(.A(G15gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT30), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT31), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n559_), .A2(new_n560_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n565_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n417_), .A2(new_n396_), .A3(new_n557_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n567_), .B1(new_n568_), .B2(new_n558_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT83), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n528_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n566_), .A2(new_n569_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT83), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(new_n529_), .A3(new_n571_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n555_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n440_), .A2(KEYINPUT90), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(G228gat), .A3(G233gat), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT29), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n512_), .B2(new_n520_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G78gat), .B1(new_n585_), .B2(new_n385_), .ZN(new_n586_));
  INV_X1    g385(.A(G78gat), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n587_), .B(new_n440_), .C1(new_n544_), .C2(new_n584_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n586_), .A2(new_n588_), .A3(G106gat), .ZN(new_n589_));
  AOI21_X1  g388(.A(G106gat), .B1(new_n586_), .B2(new_n588_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n583_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(G106gat), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n498_), .A2(new_n499_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n509_), .B1(new_n517_), .B2(KEYINPUT1), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n506_), .A2(new_n507_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n593_), .B1(new_n596_), .B2(new_n542_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT3), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n499_), .B(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT2), .B1(new_n496_), .B2(new_n497_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n518_), .B1(new_n601_), .B2(new_n514_), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT29), .B1(new_n597_), .B2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n587_), .B1(new_n603_), .B2(new_n440_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n585_), .A2(G78gat), .A3(new_n385_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n592_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n586_), .A2(new_n588_), .A3(G106gat), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(new_n607_), .A3(new_n582_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT28), .B1(new_n527_), .B2(KEYINPUT29), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT28), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n544_), .A2(new_n610_), .A3(new_n584_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G22gat), .B(G50gat), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n609_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n591_), .A2(new_n608_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n616_), .B1(new_n591_), .B2(new_n608_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n470_), .A2(new_n580_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT103), .ZN(new_n623_));
  INV_X1    g422(.A(new_n616_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n589_), .A2(new_n590_), .A3(new_n583_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n582_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n624_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n627_), .A2(new_n617_), .B1(new_n549_), .B2(new_n553_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n525_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(new_n631_), .A3(new_n476_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n524_), .A2(new_n525_), .A3(new_n531_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT97), .B1(new_n629_), .B2(new_n477_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n532_), .A2(KEYINPUT33), .A3(new_n533_), .A4(new_n477_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n456_), .A2(new_n635_), .A3(new_n444_), .A4(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n547_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n547_), .A2(KEYINPUT96), .A3(new_n638_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n426_), .A2(KEYINPUT32), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n464_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n447_), .A2(new_n420_), .A3(new_n645_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n647_), .B(new_n648_), .C1(new_n534_), .C2(new_n548_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n644_), .B1(new_n464_), .B2(new_n646_), .ZN(new_n650_));
  OAI22_X1  g449(.A1(new_n637_), .A2(new_n643_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  AOI22_X1  g450(.A1(new_n470_), .A2(new_n628_), .B1(new_n620_), .B2(new_n651_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n574_), .A2(KEYINPUT84), .A3(new_n577_), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT84), .B1(new_n574_), .B2(new_n577_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n623_), .B1(new_n652_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n467_), .A2(new_n469_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT102), .B1(new_n457_), .B2(new_n340_), .ZN(new_n658_));
  AOI211_X1 g457(.A(new_n450_), .B(KEYINPUT27), .C1(new_n456_), .C2(new_n444_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n628_), .B(new_n657_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n651_), .A2(new_n620_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n655_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(KEYINPUT103), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n622_), .B1(new_n656_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n288_), .A2(new_n316_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n290_), .A2(new_n316_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(G229gat), .A2(G233gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n290_), .B(new_n316_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n668_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n669_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(G113gat), .B(G141gat), .ZN(new_n675_));
  XNOR2_X1  g474(.A(G169gat), .B(G197gat), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n675_), .B(new_n676_), .Z(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n677_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n673_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n665_), .A2(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n339_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n311_), .A3(new_n555_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT38), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n304_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n665_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n336_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT104), .B1(new_n272_), .B2(new_n682_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n273_), .A2(new_n692_), .A3(new_n681_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n689_), .A2(new_n690_), .A3(new_n691_), .A4(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G1gat), .B1(new_n694_), .B2(new_n554_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n685_), .A2(new_n686_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n687_), .A2(new_n695_), .A3(new_n696_), .ZN(G1324gat));
  OAI21_X1  g496(.A(G8gat), .B1(new_n694_), .B2(new_n470_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(KEYINPUT105), .A2(KEYINPUT39), .ZN(new_n699_));
  AND2_X1   g498(.A1(KEYINPUT105), .A2(KEYINPUT39), .ZN(new_n700_));
  OR3_X1    g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n470_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n684_), .A2(new_n312_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n698_), .A2(new_n699_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n701_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT40), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n701_), .A2(new_n703_), .A3(KEYINPUT40), .A4(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1325gat));
  OAI21_X1  g508(.A(G15gat), .B1(new_n694_), .B2(new_n663_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT41), .Z(new_n711_));
  NAND3_X1  g510(.A1(new_n684_), .A2(new_n562_), .A3(new_n655_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1326gat));
  INV_X1    g512(.A(G22gat), .ZN(new_n714_));
  INV_X1    g513(.A(new_n620_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n684_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n694_), .A2(new_n620_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(new_n714_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n718_), .A2(new_n719_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n716_), .B1(new_n720_), .B2(new_n721_), .ZN(G1327gat));
  NOR2_X1   g521(.A1(new_n690_), .A2(new_n304_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT107), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(new_n272_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n683_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G29gat), .B1(new_n727_), .B2(new_n555_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n693_), .A2(new_n336_), .A3(new_n691_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n665_), .B2(new_n308_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT103), .B1(new_n662_), .B2(new_n663_), .ZN(new_n731_));
  AOI211_X1 g530(.A(new_n623_), .B(new_n655_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n621_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n309_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n729_), .B1(new_n730_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT44), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n737_), .A2(G29gat), .A3(new_n555_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n665_), .A2(KEYINPUT43), .A3(new_n308_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n734_), .B1(new_n733_), .B2(new_n309_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n739_), .B1(new_n742_), .B2(new_n729_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n728_), .B1(new_n738_), .B2(new_n743_), .ZN(G1328gat));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n748_));
  INV_X1    g547(.A(G36gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n470_), .B1(new_n736_), .B2(KEYINPUT44), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(new_n743_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n683_), .A2(new_n749_), .A3(new_n702_), .A4(new_n725_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT45), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n747_), .B(new_n748_), .C1(new_n751_), .C2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n750_), .A2(new_n743_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(G36gat), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n757_), .A2(new_n745_), .A3(new_n746_), .A4(new_n753_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n755_), .A2(new_n758_), .ZN(G1329gat));
  INV_X1    g558(.A(G43gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(new_n726_), .B2(new_n663_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT109), .ZN(new_n762_));
  INV_X1    g561(.A(new_n743_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n737_), .A2(G43gat), .A3(new_n578_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n762_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT47), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n762_), .B(new_n767_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1330gat));
  AOI21_X1  g568(.A(G50gat), .B1(new_n727_), .B2(new_n715_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n737_), .A2(G50gat), .A3(new_n715_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n743_), .ZN(G1331gat));
  NAND3_X1  g571(.A1(new_n329_), .A2(new_n682_), .A3(new_n335_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n273_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n689_), .A2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G57gat), .B1(new_n775_), .B2(new_n554_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n665_), .A2(new_n681_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n337_), .A2(new_n272_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n554_), .A2(G57gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n776_), .B1(new_n780_), .B2(new_n781_), .ZN(G1332gat));
  NAND3_X1  g581(.A1(new_n689_), .A2(new_n702_), .A3(new_n774_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT48), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n783_), .A2(new_n784_), .A3(G64gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n783_), .B2(G64gat), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n470_), .A2(G64gat), .ZN(new_n787_));
  OAI22_X1  g586(.A1(new_n785_), .A2(new_n786_), .B1(new_n780_), .B2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT110), .ZN(G1333gat));
  OAI21_X1  g588(.A(G71gat), .B1(new_n775_), .B2(new_n663_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT49), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n663_), .A2(G71gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n780_), .B2(new_n792_), .ZN(G1334gat));
  NAND3_X1  g592(.A1(new_n779_), .A2(new_n587_), .A3(new_n715_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n733_), .A2(new_n774_), .A3(new_n715_), .A4(new_n304_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(G78gat), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n796_), .A2(KEYINPUT112), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(KEYINPUT112), .ZN(new_n798_));
  XOR2_X1   g597(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n799_));
  AND3_X1   g598(.A1(new_n797_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n794_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT113), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n804_), .B(new_n794_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1335gat));
  NOR2_X1   g605(.A1(new_n554_), .A2(new_n219_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n730_), .A2(new_n735_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n272_), .A2(new_n682_), .A3(new_n336_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n808_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  AOI211_X1 g611(.A(KEYINPUT114), .B(new_n810_), .C1(new_n730_), .C2(new_n735_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n812_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n811_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT114), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n809_), .A2(new_n808_), .A3(new_n811_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT115), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n807_), .B1(new_n815_), .B2(new_n819_), .ZN(new_n820_));
  NOR4_X1   g619(.A1(new_n665_), .A2(new_n681_), .A3(new_n273_), .A4(new_n724_), .ZN(new_n821_));
  AOI21_X1  g620(.A(G85gat), .B1(new_n821_), .B2(new_n555_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(KEYINPUT116), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825_));
  INV_X1    g624(.A(new_n807_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n814_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n817_), .A2(KEYINPUT115), .A3(new_n818_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n826_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n825_), .B1(new_n829_), .B2(new_n822_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n824_), .A2(new_n830_), .ZN(G1336gat));
  NAND3_X1  g630(.A1(new_n821_), .A2(new_n220_), .A3(new_n702_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n470_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n220_), .ZN(G1337gat));
  INV_X1    g633(.A(new_n215_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n821_), .A2(new_n578_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n663_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n837_));
  INV_X1    g636(.A(G99gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT51), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n841_), .B(new_n836_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1338gat));
  NAND3_X1  g642(.A1(new_n821_), .A2(new_n592_), .A3(new_n715_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n809_), .A2(new_n715_), .A3(new_n811_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n845_), .A2(new_n846_), .A3(G106gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n845_), .B2(G106gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n844_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n773_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n268_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n853_), .B2(new_n268_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n263_), .A2(new_n265_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n666_), .A2(new_n667_), .A3(new_n671_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n677_), .B1(new_n670_), .B2(new_n668_), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n674_), .A2(new_n677_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n249_), .A2(new_n254_), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n240_), .A2(new_n246_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT12), .B1(new_n250_), .B2(new_n243_), .ZN(new_n868_));
  NOR4_X1   g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n865_), .A4(new_n255_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n234_), .B1(new_n253_), .B2(new_n233_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n866_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n262_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT56), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n872_), .A2(KEYINPUT56), .A3(new_n262_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n265_), .A2(new_n681_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT117), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n864_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n858_), .B1(new_n880_), .B2(new_n688_), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT56), .B1(new_n872_), .B2(new_n262_), .ZN(new_n882_));
  AOI211_X1 g681(.A(new_n874_), .B(new_n264_), .C1(new_n866_), .C2(new_n871_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n878_), .B(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n863_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(KEYINPUT57), .A3(new_n304_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n265_), .A2(new_n890_), .A3(new_n862_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n265_), .B2(new_n862_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n889_), .B1(new_n884_), .B2(new_n893_), .ZN(new_n894_));
  OAI221_X1 g693(.A(KEYINPUT58), .B1(new_n891_), .B2(new_n892_), .C1(new_n882_), .C2(new_n883_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n894_), .A2(new_n309_), .A3(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n881_), .A2(new_n888_), .A3(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n857_), .B1(new_n897_), .B2(new_n336_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n852_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  NOR4_X1   g699(.A1(new_n702_), .A2(new_n715_), .A3(new_n554_), .A4(new_n579_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n898_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n900_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n897_), .A2(new_n336_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n857_), .ZN(new_n906_));
  AOI221_X4 g705(.A(new_n902_), .B1(new_n899_), .B2(new_n852_), .C1(new_n905_), .C2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n681_), .B1(new_n904_), .B2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(G113gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n906_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n910_), .A2(KEYINPUT119), .A3(new_n901_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n898_), .B2(new_n902_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n682_), .A2(G113gat), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n911_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n851_), .B1(new_n909_), .B2(new_n916_), .ZN(new_n917_));
  AOI211_X1 g716(.A(KEYINPUT121), .B(new_n915_), .C1(new_n908_), .C2(G113gat), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1340gat));
  INV_X1    g718(.A(new_n904_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n907_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n273_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT60), .ZN(new_n923_));
  AOI21_X1  g722(.A(G120gat), .B1(new_n272_), .B2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n923_), .B2(G120gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n911_), .A2(new_n913_), .A3(new_n925_), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n926_), .A2(KEYINPUT122), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(KEYINPUT122), .ZN(new_n928_));
  OAI22_X1  g727(.A1(new_n922_), .A2(new_n483_), .B1(new_n927_), .B2(new_n928_), .ZN(G1341gat));
  NAND2_X1  g728(.A1(new_n920_), .A2(new_n921_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n690_), .A2(G127gat), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT123), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n911_), .A2(new_n913_), .A3(new_n690_), .ZN(new_n933_));
  AOI22_X1  g732(.A1(new_n930_), .A2(new_n932_), .B1(new_n480_), .B2(new_n933_), .ZN(G1342gat));
  XOR2_X1   g733(.A(KEYINPUT124), .B(G134gat), .Z(new_n935_));
  NOR2_X1   g734(.A1(new_n308_), .A2(new_n935_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n911_), .A2(new_n913_), .A3(new_n688_), .ZN(new_n937_));
  AOI22_X1  g736(.A1(new_n930_), .A2(new_n936_), .B1(new_n478_), .B2(new_n937_), .ZN(G1343gat));
  NOR2_X1   g737(.A1(new_n898_), .A2(new_n655_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n702_), .A2(new_n554_), .A3(new_n620_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n681_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g743(.A1(new_n942_), .A2(new_n272_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g745(.A1(new_n942_), .A2(new_n690_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(KEYINPUT61), .B(G155gat), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n947_), .B(new_n948_), .ZN(G1346gat));
  OR3_X1    g748(.A1(new_n941_), .A2(G162gat), .A3(new_n304_), .ZN(new_n950_));
  OAI21_X1  g749(.A(G162gat), .B1(new_n941_), .B2(new_n308_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1347gat));
  NOR2_X1   g751(.A1(new_n715_), .A2(new_n555_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n702_), .A2(new_n953_), .A3(new_n655_), .ZN(new_n954_));
  INV_X1    g753(.A(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n910_), .A2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n898_), .A2(new_n954_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(KEYINPUT125), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n958_), .A2(new_n960_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n961_), .A2(new_n353_), .A3(new_n681_), .ZN(new_n962_));
  OAI21_X1  g761(.A(G169gat), .B1(new_n956_), .B2(new_n682_), .ZN(new_n963_));
  AND2_X1   g762(.A1(new_n963_), .A2(KEYINPUT62), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n963_), .A2(KEYINPUT62), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n962_), .B1(new_n964_), .B2(new_n965_), .ZN(G1348gat));
  NAND3_X1  g765(.A1(new_n961_), .A2(new_n354_), .A3(new_n272_), .ZN(new_n967_));
  OAI21_X1  g766(.A(G176gat), .B1(new_n956_), .B2(new_n273_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(new_n968_), .ZN(G1349gat));
  NAND2_X1  g768(.A1(new_n959_), .A2(new_n690_), .ZN(new_n970_));
  OR2_X1    g769(.A1(new_n970_), .A2(KEYINPUT126), .ZN(new_n971_));
  AOI21_X1  g770(.A(G183gat), .B1(new_n970_), .B2(KEYINPUT126), .ZN(new_n972_));
  NOR2_X1   g771(.A1(new_n336_), .A2(new_n365_), .ZN(new_n973_));
  AOI22_X1  g772(.A1(new_n971_), .A2(new_n972_), .B1(new_n961_), .B2(new_n973_), .ZN(G1350gat));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n961_), .A2(new_n366_), .A3(new_n688_), .ZN(new_n976_));
  INV_X1    g775(.A(new_n976_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n308_), .B1(new_n958_), .B2(new_n960_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n978_), .A2(new_n400_), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n975_), .B1(new_n977_), .B2(new_n979_), .ZN(new_n980_));
  OAI211_X1 g779(.A(new_n976_), .B(KEYINPUT127), .C1(new_n400_), .C2(new_n978_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n980_), .A2(new_n981_), .ZN(G1351gat));
  NOR3_X1   g781(.A1(new_n470_), .A2(new_n555_), .A3(new_n620_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n939_), .A2(new_n983_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n984_), .A2(new_n682_), .ZN(new_n985_));
  XNOR2_X1  g784(.A(new_n985_), .B(new_n372_), .ZN(G1352gat));
  NOR2_X1   g785(.A1(new_n984_), .A2(new_n273_), .ZN(new_n987_));
  XNOR2_X1  g786(.A(new_n987_), .B(new_n370_), .ZN(G1353gat));
  INV_X1    g787(.A(new_n984_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n989_), .A2(new_n690_), .ZN(new_n990_));
  NOR2_X1   g789(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n991_));
  AND2_X1   g790(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n992_));
  NOR3_X1   g791(.A1(new_n990_), .A2(new_n991_), .A3(new_n992_), .ZN(new_n993_));
  AOI21_X1  g792(.A(new_n993_), .B1(new_n990_), .B2(new_n991_), .ZN(G1354gat));
  OR3_X1    g793(.A1(new_n984_), .A2(G218gat), .A3(new_n304_), .ZN(new_n995_));
  OAI21_X1  g794(.A(G218gat), .B1(new_n984_), .B2(new_n308_), .ZN(new_n996_));
  NAND2_X1  g795(.A1(new_n995_), .A2(new_n996_), .ZN(G1355gat));
endmodule


