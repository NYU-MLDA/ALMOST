//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_;
  XNOR2_X1  g000(.A(KEYINPUT0), .B(G57gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(G1gat), .B(G29gat), .Z(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(G225gat), .A2(G233gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n206_), .B(KEYINPUT97), .Z(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  AND2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G141gat), .ZN(new_n214_));
  INV_X1    g013(.A(G148gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  AOI22_X1  g015(.A1(new_n209_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT84), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT86), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT85), .ZN(new_n223_));
  OR3_X1    g022(.A1(new_n216_), .A2(new_n223_), .A3(KEYINPUT3), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n223_), .B1(new_n216_), .B2(KEYINPUT3), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G141gat), .A2(G148gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT2), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n222_), .A2(new_n224_), .A3(new_n225_), .A4(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n228_), .A2(KEYINPUT87), .A3(new_n211_), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT87), .B1(new_n228_), .B2(new_n211_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G113gat), .B(G120gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT81), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(G113gat), .A2(G120gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G113gat), .A2(G120gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(KEYINPUT81), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G127gat), .B(G134gat), .Z(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT83), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n238_), .A2(new_n240_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(KEYINPUT82), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n239_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT82), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n246_), .A2(new_n247_), .A3(KEYINPUT83), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n242_), .B1(new_n245_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n244_), .A2(KEYINPUT82), .A3(new_n243_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT83), .B1(new_n246_), .B2(new_n247_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(new_n241_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n220_), .A2(new_n231_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n228_), .A2(new_n211_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT87), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n242_), .A2(new_n244_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n228_), .A2(KEYINPUT87), .A3(new_n211_), .ZN(new_n258_));
  AND4_X1   g057(.A1(new_n220_), .A2(new_n256_), .A3(new_n257_), .A4(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT4), .B1(new_n253_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n249_), .A2(new_n252_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n256_), .A2(new_n220_), .A3(new_n258_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT4), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n208_), .B1(new_n260_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n252_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n241_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n262_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n231_), .A2(new_n220_), .A3(new_n257_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n270_), .A2(new_n207_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n205_), .B1(new_n265_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT100), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n207_), .B1(new_n275_), .B2(new_n263_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n271_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n205_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n272_), .A2(new_n273_), .A3(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n276_), .A2(new_n277_), .A3(KEYINPUT100), .A4(new_n278_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G22gat), .B(G50gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G197gat), .B(G204gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT21), .ZN(new_n286_));
  NOR3_X1   g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT90), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT90), .ZN(new_n289_));
  XOR2_X1   g088(.A(G197gat), .B(G204gat), .Z(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT21), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n291_), .B2(new_n284_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n288_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G204gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(G197gat), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n286_), .B1(new_n295_), .B2(KEYINPUT89), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(new_n285_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n284_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n262_), .B2(KEYINPUT29), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(KEYINPUT29), .B2(new_n262_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n303_));
  OR3_X1    g102(.A1(new_n262_), .A2(KEYINPUT29), .A3(new_n299_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n303_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n283_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n302_), .A2(new_n304_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n303_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n283_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  OAI211_X1 g112(.A(G228gat), .B(G233gat), .C1(new_n300_), .C2(KEYINPUT91), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G78gat), .B(G106gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  AND3_X1   g115(.A1(new_n307_), .A2(new_n313_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n316_), .B1(new_n307_), .B2(new_n313_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT18), .B(G64gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(G92gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G8gat), .B(G36gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325_));
  OR2_X1    g124(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(G176gat), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT94), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n325_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(KEYINPUT94), .A2(G169gat), .A3(G176gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT23), .ZN(new_n333_));
  OR2_X1    g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n333_), .A2(KEYINPUT95), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT95), .B1(new_n333_), .B2(new_n334_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n330_), .B(new_n331_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n332_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT24), .ZN(new_n340_));
  OR3_X1    g139(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n339_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n341_), .A2(KEYINPUT24), .A3(new_n342_), .A4(new_n325_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT25), .B(G183gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT26), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G190gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G190gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT26), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n344_), .B(new_n345_), .C1(new_n349_), .C2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n337_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n299_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT96), .ZN(new_n356_));
  XOR2_X1   g155(.A(KEYINPUT77), .B(G190gat), .Z(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(new_n347_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n344_), .B(new_n345_), .C1(new_n358_), .C2(new_n349_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n333_), .B1(G183gat), .B2(new_n357_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n328_), .A2(KEYINPUT79), .ZN(new_n361_));
  NOR2_X1   g160(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n362_));
  OAI21_X1  g161(.A(G169gat), .B1(new_n362_), .B2(G176gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n359_), .A2(new_n364_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n365_), .A2(new_n299_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT96), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n354_), .A2(new_n367_), .A3(new_n299_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n356_), .A2(KEYINPUT20), .A3(new_n366_), .A4(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(KEYINPUT92), .Z(new_n371_));
  XOR2_X1   g170(.A(new_n371_), .B(KEYINPUT19), .Z(new_n372_));
  XOR2_X1   g171(.A(new_n372_), .B(KEYINPUT93), .Z(new_n373_));
  NAND2_X1  g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n365_), .A2(new_n299_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n372_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT20), .B1(new_n354_), .B2(new_n299_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n324_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n374_), .A2(new_n324_), .A3(new_n379_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT27), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  AOI211_X1 g182(.A(new_n323_), .B(new_n378_), .C1(new_n369_), .C2(new_n373_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT98), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n377_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(KEYINPUT98), .B(KEYINPUT20), .C1(new_n354_), .C2(new_n299_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n375_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n372_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT99), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n369_), .A2(new_n373_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n388_), .A2(KEYINPUT99), .A3(new_n389_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n384_), .B1(new_n395_), .B2(new_n323_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n383_), .B1(new_n396_), .B2(KEYINPUT27), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G71gat), .B(G99gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n365_), .B(KEYINPUT30), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(new_n261_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G15gat), .B(G43gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT80), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT31), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n403_), .A2(new_n406_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n401_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n409_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(new_n407_), .A3(new_n400_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  AND4_X1   g212(.A1(new_n282_), .A2(new_n319_), .A3(new_n397_), .A4(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n324_), .A2(KEYINPUT32), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n395_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n324_), .A2(KEYINPUT32), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n374_), .A2(new_n379_), .A3(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n280_), .A2(new_n417_), .A3(new_n281_), .A4(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n420_), .A2(KEYINPUT101), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(KEYINPUT101), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n279_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n384_), .A2(new_n380_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n208_), .B1(new_n275_), .B2(new_n263_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n426_), .B(new_n205_), .C1(new_n208_), .C2(new_n270_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n276_), .A2(new_n277_), .A3(KEYINPUT33), .A4(new_n278_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n424_), .A2(new_n425_), .A3(new_n427_), .A4(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n307_), .A2(new_n313_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n316_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n307_), .A2(new_n313_), .A3(new_n316_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n429_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n421_), .A2(new_n422_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n395_), .A2(new_n323_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(KEYINPUT27), .A3(new_n382_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n383_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n282_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n432_), .A2(new_n433_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n413_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n415_), .B1(new_n435_), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G71gat), .B(G78gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(G57gat), .A2(G64gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT11), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G57gat), .A2(G64gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n450_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT11), .B1(new_n452_), .B2(new_n447_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n446_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n445_), .B(KEYINPUT11), .C1(new_n447_), .C2(new_n452_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G231gat), .A2(G233gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G1gat), .ZN(new_n459_));
  INV_X1    g258(.A(G8gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT14), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G15gat), .ZN(new_n462_));
  INV_X1    g261(.A(G22gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G15gat), .A2(G22gat), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n461_), .A2(KEYINPUT73), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n466_), .B1(KEYINPUT73), .B2(new_n461_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G1gat), .B(G8gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT74), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n467_), .B(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n458_), .B(new_n470_), .Z(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n472_), .A2(KEYINPUT75), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT16), .B(G183gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(G211gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(G127gat), .B(G155gat), .Z(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT17), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n473_), .B(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n472_), .A2(new_n478_), .A3(new_n477_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n482_), .B(KEYINPUT76), .Z(new_n483_));
  XNOR2_X1  g282(.A(G190gat), .B(G218gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(G134gat), .ZN(new_n485_));
  INV_X1    g284(.A(G162gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n488_), .A2(KEYINPUT36), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G29gat), .B(G36gat), .ZN(new_n490_));
  INV_X1    g289(.A(G43gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G50gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n490_), .B(G43gat), .ZN(new_n494_));
  INV_X1    g293(.A(G50gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT15), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n493_), .A2(new_n496_), .A3(KEYINPUT15), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(G85gat), .A2(G92gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT9), .ZN(new_n506_));
  INV_X1    g305(.A(G106gat), .ZN(new_n507_));
  INV_X1    g306(.A(G99gat), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n508_), .A2(KEYINPUT10), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(KEYINPUT10), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n507_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT6), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n502_), .A2(KEYINPUT9), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n506_), .A2(new_n511_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT7), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(new_n508_), .A3(new_n507_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n520_), .A2(new_n514_), .A3(new_n515_), .A4(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT8), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT64), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n503_), .A2(new_n504_), .A3(new_n524_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n522_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n523_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n518_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT65), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  OAI211_X1 g329(.A(KEYINPUT65), .B(new_n518_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n501_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n497_), .A2(new_n528_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n534_), .A2(KEYINPUT66), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(KEYINPUT66), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n533_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT34), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n539_), .A2(KEYINPUT35), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n537_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n533_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT67), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n542_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n547_), .B2(new_n542_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n489_), .B(new_n546_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT68), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT67), .B1(new_n537_), .B2(new_n543_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n547_), .A2(new_n548_), .A3(new_n542_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n556_), .A2(KEYINPUT68), .A3(new_n489_), .A4(new_n546_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n553_), .A2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n546_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n487_), .B(KEYINPUT36), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT70), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT72), .B1(new_n563_), .B2(KEYINPUT37), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n553_), .A2(new_n557_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT72), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT37), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n558_), .A2(KEYINPUT69), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT69), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n553_), .A2(new_n557_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT71), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n562_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n559_), .A2(KEYINPUT71), .A3(new_n561_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n570_), .A2(new_n572_), .A3(new_n574_), .A4(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT37), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n483_), .B1(new_n569_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n456_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT12), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n522_), .A2(new_n525_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT8), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n522_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT65), .B1(new_n585_), .B2(new_n518_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n531_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n581_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT12), .B1(new_n528_), .B2(new_n579_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n456_), .B(new_n518_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n588_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n593_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n456_), .B1(new_n585_), .B2(new_n518_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n595_), .B1(new_n596_), .B2(new_n591_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(new_n294_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT5), .ZN(new_n601_));
  INV_X1    g400(.A(G176gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n594_), .A2(new_n597_), .A3(new_n603_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n607_), .A2(KEYINPUT13), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(KEYINPUT13), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n470_), .A2(new_n497_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n470_), .B2(new_n501_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n470_), .B(new_n497_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(G229gat), .A3(G233gat), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G113gat), .B(G141gat), .ZN(new_n619_));
  INV_X1    g418(.A(G169gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(G197gat), .Z(new_n622_));
  OR2_X1    g421(.A1(new_n618_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n618_), .A2(new_n622_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n611_), .A2(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n444_), .A2(new_n578_), .A3(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n280_), .A2(new_n281_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n459_), .A3(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n444_), .A2(new_n482_), .A3(new_n627_), .A4(new_n563_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G1gat), .B1(new_n633_), .B2(new_n282_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(G1324gat));
  INV_X1    g434(.A(new_n633_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n397_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(KEYINPUT103), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n633_), .B2(new_n397_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(G8gat), .A3(new_n640_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n641_), .A2(KEYINPUT104), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(KEYINPUT104), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(KEYINPUT39), .A3(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n628_), .A2(new_n460_), .A3(new_n637_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n641_), .A2(KEYINPUT104), .A3(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n644_), .A2(new_n645_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(G1325gat));
  OAI21_X1  g449(.A(G15gat), .B1(new_n633_), .B2(new_n442_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT105), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT41), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n628_), .A2(new_n462_), .A3(new_n413_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1326gat));
  OAI21_X1  g454(.A(G22gat), .B1(new_n633_), .B2(new_n319_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT42), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n628_), .A2(new_n463_), .A3(new_n440_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1327gat));
  INV_X1    g458(.A(G29gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n483_), .A2(new_n627_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n663_));
  AOI22_X1  g462(.A1(new_n564_), .A2(new_n568_), .B1(new_n576_), .B2(KEYINPUT37), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n444_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n629_), .A2(new_n666_), .A3(new_n419_), .A4(new_n417_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n434_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n420_), .A2(KEYINPUT101), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n413_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n414_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n572_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n574_), .A2(new_n575_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n571_), .B1(new_n553_), .B2(new_n557_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n673_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n566_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n678_));
  OAI22_X1  g477(.A1(new_n676_), .A2(new_n567_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT43), .B1(new_n672_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n665_), .A2(new_n680_), .ZN(new_n681_));
  OR2_X1    g480(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT107), .B1(KEYINPUT106), .B2(KEYINPUT44), .ZN(new_n683_));
  AND4_X1   g482(.A1(new_n662_), .A2(new_n681_), .A3(new_n682_), .A4(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n661_), .B1(new_n665_), .B2(new_n680_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n683_), .B1(new_n686_), .B2(new_n682_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n660_), .B(new_n282_), .C1(new_n685_), .C2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n444_), .A2(new_n565_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n661_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n629_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n689_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT108), .ZN(G1328gat));
  INV_X1    g493(.A(KEYINPUT111), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n637_), .B1(new_n684_), .B2(new_n687_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT109), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT109), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n699_), .B(new_n637_), .C1(new_n684_), .C2(new_n687_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(G36gat), .A3(new_n700_), .ZN(new_n701_));
  NOR4_X1   g500(.A1(new_n690_), .A2(G36gat), .A3(new_n397_), .A4(new_n661_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(new_n704_));
  AOI211_X1 g503(.A(new_n695_), .B(new_n696_), .C1(new_n701_), .C2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n695_), .A2(new_n696_), .ZN(new_n707_));
  AND4_X1   g506(.A1(new_n706_), .A2(new_n701_), .A3(new_n707_), .A4(new_n704_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n705_), .A2(new_n708_), .ZN(G1329gat));
  INV_X1    g508(.A(KEYINPUT47), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n413_), .B1(new_n684_), .B2(new_n687_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G43gat), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n691_), .A2(new_n491_), .A3(new_n413_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n712_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n713_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n710_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n717_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(KEYINPUT47), .A3(new_n715_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1330gat));
  AOI21_X1  g520(.A(G50gat), .B1(new_n691_), .B2(new_n440_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n319_), .B1(new_n685_), .B2(new_n688_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(G50gat), .ZN(G1331gat));
  NOR4_X1   g523(.A1(new_n672_), .A2(new_n625_), .A3(new_n610_), .A4(new_n483_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n563_), .ZN(new_n726_));
  INV_X1    g525(.A(G57gat), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n282_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n679_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n629_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n728_), .B1(new_n727_), .B2(new_n731_), .ZN(G1332gat));
  OR3_X1    g531(.A1(new_n729_), .A2(G64gat), .A3(new_n397_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G64gat), .B1(new_n726_), .B2(new_n397_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n734_), .A2(KEYINPUT113), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(KEYINPUT113), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(KEYINPUT48), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT48), .B1(new_n735_), .B2(new_n736_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n733_), .B1(new_n737_), .B2(new_n738_), .ZN(G1333gat));
  OAI21_X1  g538(.A(G71gat), .B1(new_n726_), .B2(new_n442_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT49), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n442_), .A2(G71gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n729_), .B2(new_n742_), .ZN(G1334gat));
  OAI21_X1  g542(.A(G78gat), .B1(new_n726_), .B2(new_n319_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT50), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n319_), .A2(G78gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n729_), .B2(new_n746_), .ZN(G1335gat));
  NAND3_X1  g546(.A1(new_n483_), .A2(new_n626_), .A3(new_n611_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n690_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G85gat), .B1(new_n749_), .B2(new_n629_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(new_n665_), .B2(new_n680_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n629_), .A2(G85gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n750_), .B1(new_n751_), .B2(new_n752_), .ZN(G1336gat));
  AOI21_X1  g552(.A(G92gat), .B1(new_n749_), .B2(new_n637_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n637_), .A2(G92gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n751_), .B2(new_n755_), .ZN(G1337gat));
  AOI21_X1  g555(.A(new_n508_), .B1(new_n751_), .B2(new_n413_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n509_), .A2(new_n510_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n442_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n757_), .B1(new_n749_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT51), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n760_), .B(new_n762_), .ZN(G1338gat));
  NAND3_X1  g562(.A1(new_n749_), .A2(new_n507_), .A3(new_n440_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n751_), .A2(new_n440_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G106gat), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(KEYINPUT52), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(KEYINPUT52), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g569(.A1(new_n610_), .A2(new_n626_), .ZN(new_n771_));
  NOR4_X1   g570(.A1(new_n664_), .A2(KEYINPUT54), .A3(new_n483_), .A4(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773_));
  INV_X1    g572(.A(new_n771_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n578_), .B2(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n772_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n594_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n778_), .B1(new_n594_), .B2(new_n779_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n588_), .A2(new_n592_), .A3(KEYINPUT55), .A4(new_n593_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n590_), .B1(new_n596_), .B2(KEYINPUT12), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n580_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n595_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n782_), .A2(new_n785_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n780_), .A2(new_n781_), .A3(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n777_), .B1(new_n787_), .B2(new_n603_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n594_), .A2(new_n779_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT115), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n594_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n790_), .A2(new_n782_), .A3(new_n785_), .A4(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(KEYINPUT56), .A3(new_n604_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n788_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n616_), .A2(new_n614_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n613_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n622_), .B(new_n795_), .C1(new_n796_), .C2(new_n614_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n623_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n794_), .A2(new_n606_), .A3(new_n798_), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n799_), .B(KEYINPUT58), .Z(new_n800_));
  NOR2_X1   g599(.A1(new_n679_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n788_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT116), .B(new_n777_), .C1(new_n787_), .C2(new_n603_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n793_), .A3(new_n805_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n625_), .A2(new_n606_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT117), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n798_), .A2(new_n607_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n806_), .A2(new_n811_), .A3(new_n807_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n563_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT57), .B1(new_n814_), .B2(KEYINPUT118), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  AOI211_X1 g616(.A(new_n816_), .B(new_n817_), .C1(new_n813_), .C2(new_n563_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n802_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n482_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n776_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n637_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n629_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(G113gat), .B1(new_n824_), .B2(new_n625_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n806_), .A2(new_n811_), .A3(new_n807_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n811_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n810_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT118), .B1(new_n830_), .B2(new_n565_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n817_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n814_), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n801_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n483_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n826_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n776_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n819_), .A2(KEYINPUT120), .A3(new_n483_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  INV_X1    g639(.A(new_n823_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT121), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT59), .B1(new_n821_), .B2(new_n823_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT119), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n846_), .B(KEYINPUT59), .C1(new_n821_), .C2(new_n823_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n839_), .A2(new_n849_), .A3(new_n840_), .A4(new_n841_), .ZN(new_n850_));
  AND4_X1   g649(.A1(new_n625_), .A2(new_n843_), .A3(new_n848_), .A4(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n825_), .B1(new_n851_), .B2(G113gat), .ZN(G1340gat));
  NAND4_X1  g651(.A1(new_n843_), .A2(new_n848_), .A3(new_n611_), .A4(new_n850_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(G120gat), .ZN(new_n854_));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n610_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n824_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n855_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(new_n857_), .ZN(G1341gat));
  AOI21_X1  g657(.A(G127gat), .B1(new_n824_), .B2(new_n835_), .ZN(new_n859_));
  AND4_X1   g658(.A1(new_n482_), .A2(new_n843_), .A3(new_n848_), .A4(new_n850_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g660(.A(G134gat), .B1(new_n824_), .B2(new_n565_), .ZN(new_n862_));
  AND4_X1   g661(.A1(G134gat), .A2(new_n843_), .A3(new_n848_), .A4(new_n850_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n664_), .ZN(G1343gat));
  NOR2_X1   g663(.A1(new_n319_), .A2(new_n413_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n821_), .A2(new_n282_), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n397_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n626_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n214_), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n610_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n215_), .ZN(G1345gat));
  NOR2_X1   g671(.A1(new_n868_), .A2(new_n483_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XOR2_X1   g673(.A(new_n873_), .B(new_n874_), .Z(G1346gat));
  NOR3_X1   g674(.A1(new_n868_), .A2(new_n486_), .A3(new_n679_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n867_), .A2(new_n397_), .A3(new_n565_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n486_), .B2(new_n877_), .ZN(G1347gat));
  NOR2_X1   g677(.A1(new_n397_), .A2(new_n629_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n880_), .A2(new_n442_), .A3(new_n440_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n839_), .A2(new_n625_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(G169gat), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT122), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n882_), .A2(new_n885_), .A3(G169gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n884_), .A2(KEYINPUT62), .A3(new_n886_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n326_), .A2(new_n327_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n882_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n883_), .A2(KEYINPUT122), .A3(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n887_), .A2(new_n889_), .A3(new_n891_), .ZN(G1348gat));
  NAND2_X1  g691(.A1(new_n839_), .A2(new_n881_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n602_), .B1(new_n893_), .B2(new_n610_), .ZN(new_n894_));
  NOR4_X1   g693(.A1(new_n821_), .A2(new_n440_), .A3(new_n442_), .A4(new_n880_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(G176gat), .A3(new_n611_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n894_), .A2(KEYINPUT123), .A3(new_n896_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1349gat));
  NOR3_X1   g700(.A1(new_n893_), .A2(new_n820_), .A3(new_n346_), .ZN(new_n902_));
  AOI21_X1  g701(.A(G183gat), .B1(new_n895_), .B2(new_n835_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n893_), .B2(new_n679_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n565_), .A2(new_n348_), .A3(new_n351_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n893_), .B2(new_n906_), .ZN(G1351gat));
  NOR3_X1   g706(.A1(new_n821_), .A2(new_n866_), .A3(new_n880_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n625_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g709(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n911_));
  INV_X1    g710(.A(new_n908_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n610_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n911_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n915_), .B1(new_n913_), .B2(new_n911_), .ZN(G1353gat));
  INV_X1    g715(.A(KEYINPUT63), .ZN(new_n917_));
  INV_X1    g716(.A(G211gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n482_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n919_), .A2(new_n920_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n908_), .A2(new_n922_), .A3(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT126), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n908_), .A2(new_n926_), .A3(new_n922_), .A4(new_n923_), .ZN(new_n927_));
  AND4_X1   g726(.A1(new_n917_), .A2(new_n925_), .A3(new_n918_), .A4(new_n927_), .ZN(new_n928_));
  AOI22_X1  g727(.A1(new_n925_), .A2(new_n927_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1354gat));
  AOI21_X1  g729(.A(G218gat), .B1(new_n908_), .B2(new_n565_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n908_), .A2(G218gat), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n932_), .B2(new_n664_), .ZN(G1355gat));
endmodule


