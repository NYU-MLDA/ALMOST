//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_;
  XNOR2_X1  g000(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT35), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G29gat), .B(G36gat), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT69), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(KEYINPUT69), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G43gat), .B(G50gat), .Z(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n211_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n208_), .A2(new_n209_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n216_));
  XOR2_X1   g015(.A(new_n215_), .B(new_n216_), .Z(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT6), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  OR3_X1    g020(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G85gat), .B(G92gat), .Z(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT8), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n223_), .A2(new_n228_), .A3(new_n224_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n226_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT10), .B(G99gat), .Z(new_n231_));
  INV_X1    g030(.A(G106gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n224_), .A2(KEYINPUT9), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT9), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G85gat), .A3(G92gat), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n233_), .A2(new_n234_), .A3(new_n220_), .A4(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n230_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n226_), .A2(new_n229_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT64), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n238_), .A2(KEYINPUT65), .A3(new_n240_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n218_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n239_), .A2(new_n237_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(new_n215_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n247_), .B1(new_n205_), .B2(new_n204_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n206_), .B1(new_n245_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n206_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n238_), .A2(KEYINPUT65), .A3(new_n240_), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT65), .B1(new_n238_), .B2(new_n240_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n251_), .B(new_n248_), .C1(new_n254_), .C2(new_n218_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G190gat), .B(G218gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT71), .ZN(new_n257_));
  XOR2_X1   g056(.A(G134gat), .B(G162gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(KEYINPUT36), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n250_), .A2(new_n255_), .A3(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n263_));
  NAND3_X1  g062(.A1(new_n250_), .A2(new_n255_), .A3(KEYINPUT72), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n259_), .B(KEYINPUT36), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT72), .B1(new_n250_), .B2(new_n255_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n262_), .B(new_n263_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n262_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n265_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT37), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G15gat), .B(G22gat), .ZN(new_n275_));
  INV_X1    g074(.A(G1gat), .ZN(new_n276_));
  INV_X1    g075(.A(G8gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT14), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G8gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G231gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G57gat), .B(G64gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT11), .ZN(new_n285_));
  XOR2_X1   g084(.A(G71gat), .B(G78gat), .Z(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n286_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n284_), .A2(KEYINPUT11), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n283_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT17), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G127gat), .B(G155gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT16), .ZN(new_n294_));
  XOR2_X1   g093(.A(G183gat), .B(G211gat), .Z(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n291_), .A2(new_n292_), .A3(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(KEYINPUT17), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n297_), .B1(new_n291_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n274_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G230gat), .A2(G233gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n290_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n246_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n239_), .A2(new_n290_), .A3(new_n237_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n302_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n243_), .A2(new_n244_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(KEYINPUT12), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(KEYINPUT12), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n307_), .A2(new_n309_), .B1(new_n304_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n306_), .B1(new_n311_), .B2(new_n302_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G120gat), .B(G148gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT5), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT67), .ZN(new_n315_));
  XOR2_X1   g114(.A(G176gat), .B(G204gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n317_), .A2(KEYINPUT66), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n312_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT13), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n320_), .A2(new_n321_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n301_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n325_), .B(KEYINPUT74), .Z(new_n326_));
  NAND2_X1  g125(.A1(G226gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT19), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G197gat), .B(G204gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(G211gat), .B(G218gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n330_), .B1(KEYINPUT21), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(KEYINPUT21), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335_));
  INV_X1    g134(.A(G183gat), .ZN(new_n336_));
  INV_X1    g135(.A(G190gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n335_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n338_), .B(new_n339_), .C1(G183gat), .C2(G190gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n340_), .B(KEYINPUT93), .Z(new_n341_));
  NAND2_X1  g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n342_), .B(KEYINPUT77), .Z(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G169gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n344_), .B(KEYINPUT92), .Z(new_n345_));
  INV_X1    g144(.A(G176gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n341_), .A2(new_n343_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n338_), .A2(new_n339_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n342_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT25), .B(G183gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT91), .ZN(new_n356_));
  XOR2_X1   g155(.A(KEYINPUT26), .B(G190gat), .Z(new_n357_));
  OAI211_X1 g156(.A(new_n351_), .B(new_n354_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n334_), .B1(new_n348_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n334_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n343_), .A2(new_n353_), .ZN(new_n361_));
  OR3_X1    g160(.A1(new_n337_), .A2(KEYINPUT76), .A3(KEYINPUT26), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT26), .B1(new_n337_), .B2(KEYINPUT76), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n355_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n364_), .A3(new_n351_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n344_), .A2(new_n346_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n344_), .A2(KEYINPUT78), .A3(new_n346_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n368_), .A2(new_n343_), .A3(new_n340_), .A4(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n365_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT20), .B1(new_n360_), .B2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n329_), .B1(new_n359_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT20), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(new_n360_), .B2(new_n371_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n348_), .A2(new_n358_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(new_n360_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n373_), .B1(new_n329_), .B2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G8gat), .B(G36gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT18), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G64gat), .B(G92gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n380_), .B(new_n381_), .Z(new_n382_));
  NOR2_X1   g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n328_), .B1(new_n359_), .B2(new_n372_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n375_), .B(new_n329_), .C1(new_n376_), .C2(new_n360_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n382_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT27), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT27), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n384_), .A2(new_n385_), .A3(KEYINPUT94), .A4(new_n382_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT94), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n392_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n386_), .A2(new_n387_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n391_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n389_), .B1(new_n390_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G155gat), .A2(G162gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G155gat), .A2(G162gat), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n398_), .B1(KEYINPUT1), .B2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(KEYINPUT1), .B2(new_n399_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G141gat), .A2(G148gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(G141gat), .A2(G148gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n401_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT2), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n402_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n407_), .A2(new_n409_), .A3(new_n410_), .A4(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n417_), .A2(KEYINPUT82), .A3(new_n411_), .A4(new_n407_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n414_), .A2(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(G155gat), .A2(G162gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(new_n399_), .ZN(new_n422_));
  AND2_X1   g221(.A1(G155gat), .A2(G162gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT83), .B1(new_n423_), .B2(new_n398_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT84), .B1(new_n419_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n428_));
  AOI211_X1 g227(.A(new_n428_), .B(new_n425_), .C1(new_n414_), .C2(new_n418_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n405_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G127gat), .B(G134gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G113gat), .B(G120gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT95), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT96), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n405_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n419_), .A2(new_n426_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n428_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n419_), .A2(KEYINPUT84), .A3(new_n426_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n439_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(KEYINPUT96), .A3(new_n433_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT95), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n430_), .A2(new_n445_), .A3(new_n434_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n436_), .A2(new_n438_), .A3(new_n444_), .A4(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G225gat), .A2(G233gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n449_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT97), .B1(new_n435_), .B2(KEYINPUT4), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT97), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n430_), .A2(new_n453_), .A3(new_n454_), .A4(new_n434_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n451_), .B(new_n456_), .C1(new_n447_), .C2(new_n454_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G1gat), .B(G29gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT0), .ZN(new_n459_));
  INV_X1    g258(.A(G57gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G85gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n450_), .A2(new_n457_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n464_), .B1(new_n450_), .B2(new_n457_), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n465_), .A2(new_n466_), .A3(KEYINPUT99), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT99), .B1(new_n465_), .B2(new_n466_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n397_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G78gat), .B(G106gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT29), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n473_), .B(new_n360_), .C1(new_n443_), .C2(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(G228gat), .A2(G233gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n334_), .B1(new_n430_), .B2(KEYINPUT29), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n473_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  AOI211_X1 g280(.A(new_n473_), .B(new_n476_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n472_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT88), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n477_), .A2(new_n480_), .ZN(new_n485_));
  AOI211_X1 g284(.A(KEYINPUT86), .B(new_n334_), .C1(new_n430_), .C2(KEYINPUT29), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n475_), .B(new_n476_), .C1(new_n486_), .C2(new_n473_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n487_), .A3(new_n471_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT89), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n485_), .A2(new_n487_), .A3(new_n490_), .A4(new_n471_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT88), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n492_), .B(new_n472_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n484_), .A2(new_n489_), .A3(new_n491_), .A4(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n443_), .A2(KEYINPUT85), .A3(new_n474_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n496_), .B1(new_n430_), .B2(KEYINPUT29), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n498_), .A2(KEYINPUT28), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(KEYINPUT28), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G22gat), .B(G50gat), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n502_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n494_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT90), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n488_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n488_), .A2(new_n509_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n506_), .A2(new_n510_), .A3(new_n483_), .A4(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n433_), .B(KEYINPUT31), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n371_), .B(KEYINPUT30), .Z(new_n514_));
  XNOR2_X1  g313(.A(G71gat), .B(G99gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT80), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G227gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G15gat), .B(G43gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT79), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n518_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n514_), .B(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n513_), .B1(new_n522_), .B2(KEYINPUT81), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(KEYINPUT81), .B2(new_n522_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n522_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT81), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n513_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n508_), .A2(new_n512_), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n529_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n470_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n508_), .A2(new_n512_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n382_), .A2(KEYINPUT32), .ZN(new_n535_));
  MUX2_X1   g334(.A(new_n378_), .B(new_n386_), .S(new_n535_), .Z(new_n536_));
  OAI21_X1  g335(.A(new_n536_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT98), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n464_), .B1(new_n448_), .B2(new_n451_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n449_), .B(new_n456_), .C1(new_n447_), .C2(new_n454_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n395_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n465_), .A2(KEYINPUT33), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n450_), .A2(new_n457_), .A3(new_n464_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT33), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n542_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n536_), .B(KEYINPUT98), .C1(new_n465_), .C2(new_n466_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n539_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n534_), .A2(new_n549_), .A3(new_n528_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n532_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n217_), .A2(new_n281_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n215_), .A2(new_n281_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT75), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n215_), .B(new_n281_), .Z(new_n558_));
  INV_X1    g357(.A(new_n555_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(new_n557_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G113gat), .B(G141gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G169gat), .B(G197gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n556_), .A2(new_n557_), .A3(new_n566_), .A4(new_n560_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n326_), .A2(new_n551_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n468_), .A2(new_n469_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(new_n276_), .A3(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT38), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n324_), .A2(new_n569_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n532_), .B2(new_n550_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n262_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(new_n300_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(G1gat), .B1(new_n580_), .B2(new_n571_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n574_), .A2(new_n581_), .ZN(G1324gat));
  OAI21_X1  g381(.A(G8gat), .B1(new_n580_), .B2(new_n396_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT100), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT100), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n585_), .B(G8gat), .C1(new_n580_), .C2(new_n396_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT39), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n584_), .A2(KEYINPUT39), .A3(new_n586_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n570_), .A2(new_n277_), .A3(new_n397_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(G1325gat));
  INV_X1    g393(.A(G15gat), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n570_), .A2(new_n595_), .A3(new_n529_), .ZN(new_n596_));
  OAI21_X1  g395(.A(G15gat), .B1(new_n580_), .B2(new_n528_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n597_), .A2(KEYINPUT41), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(KEYINPUT41), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .ZN(G1326gat));
  OAI21_X1  g399(.A(G22gat), .B1(new_n580_), .B2(new_n534_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT42), .ZN(new_n602_));
  INV_X1    g401(.A(G22gat), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n570_), .A2(new_n603_), .A3(new_n533_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(G1327gat));
  NAND2_X1  g404(.A1(new_n578_), .A2(new_n300_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n576_), .A2(new_n607_), .ZN(new_n608_));
  OR3_X1    g407(.A1(new_n608_), .A2(G29gat), .A3(new_n571_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n575_), .A2(new_n299_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT43), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n268_), .A2(KEYINPUT102), .A3(new_n272_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT102), .B1(new_n268_), .B2(new_n272_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n611_), .B1(new_n551_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n274_), .A2(new_n611_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n532_), .B2(new_n550_), .ZN(new_n618_));
  OAI211_X1 g417(.A(KEYINPUT44), .B(new_n610_), .C1(new_n616_), .C2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n551_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n273_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n612_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n532_), .B2(new_n550_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n622_), .B1(new_n626_), .B2(new_n611_), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT44), .B1(new_n627_), .B2(new_n610_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n620_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n572_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n630_), .A2(KEYINPUT103), .A3(G29gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT103), .B1(new_n630_), .B2(G29gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n609_), .B1(new_n631_), .B2(new_n632_), .ZN(G1328gat));
  INV_X1    g432(.A(KEYINPUT107), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT46), .ZN(new_n635_));
  INV_X1    g434(.A(new_n608_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n396_), .B(KEYINPUT105), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(G36gat), .ZN(new_n639_));
  XOR2_X1   g438(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n636_), .A2(new_n639_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n639_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n640_), .B1(new_n608_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n619_), .A2(new_n397_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G36gat), .B1(new_n646_), .B2(new_n628_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n645_), .B1(new_n647_), .B2(KEYINPUT104), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n649_), .B(G36gat), .C1(new_n646_), .C2(new_n628_), .ZN(new_n650_));
  AOI211_X1 g449(.A(new_n634_), .B(new_n635_), .C1(new_n648_), .C2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n647_), .A2(KEYINPUT104), .ZN(new_n652_));
  INV_X1    g451(.A(new_n645_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n650_), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT46), .B1(new_n654_), .B2(KEYINPUT107), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n651_), .A2(new_n655_), .ZN(G1329gat));
  NAND3_X1  g455(.A1(new_n629_), .A2(G43gat), .A3(new_n529_), .ZN(new_n657_));
  INV_X1    g456(.A(G43gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n658_), .B1(new_n608_), .B2(new_n528_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT108), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n657_), .A2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g461(.A(G50gat), .B1(new_n636_), .B2(new_n533_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n619_), .A2(G50gat), .A3(new_n533_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n628_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n663_), .B1(new_n664_), .B2(new_n665_), .ZN(G1331gat));
  NOR2_X1   g465(.A1(new_n324_), .A2(new_n569_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n551_), .A2(new_n667_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n668_), .A2(new_n300_), .A3(new_n274_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n460_), .A3(new_n572_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n551_), .A2(new_n667_), .A3(new_n579_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G57gat), .B1(new_n671_), .B2(new_n571_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1332gat));
  OAI21_X1  g472(.A(G64gat), .B1(new_n671_), .B2(new_n638_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT48), .ZN(new_n675_));
  INV_X1    g474(.A(G64gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n669_), .A2(new_n676_), .A3(new_n637_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT109), .ZN(G1333gat));
  OAI21_X1  g478(.A(G71gat), .B1(new_n671_), .B2(new_n528_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT49), .ZN(new_n681_));
  INV_X1    g480(.A(G71gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n669_), .A2(new_n682_), .A3(new_n529_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1334gat));
  OAI21_X1  g483(.A(G78gat), .B1(new_n671_), .B2(new_n534_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT50), .ZN(new_n686_));
  INV_X1    g485(.A(G78gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n669_), .A2(new_n687_), .A3(new_n533_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1335gat));
  NAND3_X1  g488(.A1(new_n551_), .A2(new_n667_), .A3(new_n607_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(new_n462_), .A3(new_n572_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n469_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n396_), .B1(new_n693_), .B2(new_n467_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n533_), .A2(new_n528_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n508_), .A2(new_n512_), .A3(new_n529_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n508_), .A2(new_n512_), .A3(new_n528_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n539_), .A2(new_n548_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n547_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n615_), .B1(new_n697_), .B2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n618_), .B1(new_n701_), .B2(KEYINPUT43), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n667_), .A2(new_n300_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT110), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705_));
  INV_X1    g504(.A(new_n703_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n627_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n571_), .B1(new_n704_), .B2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n692_), .B1(new_n708_), .B2(new_n462_), .ZN(G1336gat));
  AOI21_X1  g508(.A(G92gat), .B1(new_n691_), .B2(new_n397_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT111), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n704_), .A2(new_n707_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n637_), .A2(G92gat), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT112), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n711_), .B1(new_n712_), .B2(new_n714_), .ZN(G1337gat));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n529_), .A2(new_n231_), .ZN(new_n717_));
  OR3_X1    g516(.A1(new_n690_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n690_), .B2(new_n717_), .ZN(new_n719_));
  AOI22_X1  g518(.A1(new_n718_), .A2(new_n719_), .B1(KEYINPUT114), .B2(KEYINPUT51), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n528_), .B1(new_n704_), .B2(new_n707_), .ZN(new_n721_));
  INV_X1    g520(.A(G99gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT115), .ZN(new_n724_));
  NOR2_X1   g523(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT115), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n726_), .B(new_n720_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n724_), .A2(new_n725_), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n725_), .B1(new_n724_), .B2(new_n727_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1338gat));
  NAND2_X1  g529(.A1(new_n627_), .A2(new_n706_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G106gat), .B1(new_n731_), .B2(new_n534_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT116), .B1(new_n732_), .B2(KEYINPUT52), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n702_), .A2(new_n703_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n232_), .B1(new_n734_), .B2(new_n533_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT116), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n735_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n732_), .A2(KEYINPUT52), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n733_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n691_), .A2(new_n232_), .A3(new_n533_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT53), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT53), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n740_), .A2(new_n744_), .A3(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1339gat));
  NOR2_X1   g545(.A1(new_n571_), .A2(new_n397_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n556_), .A2(new_n566_), .A3(new_n560_), .ZN(new_n748_));
  MUX2_X1   g547(.A(new_n558_), .B(new_n554_), .S(new_n559_), .Z(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(new_n566_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n320_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n317_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT56), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(KEYINPUT118), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n302_), .A2(KEYINPUT117), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n311_), .A2(KEYINPUT55), .A3(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n310_), .A2(new_n304_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n302_), .B(new_n758_), .C1(new_n254_), .C2(new_n308_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n757_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n756_), .B1(new_n311_), .B2(KEYINPUT55), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n752_), .B(new_n754_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n312_), .A2(new_n317_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n569_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n311_), .A2(KEYINPUT55), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n755_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n757_), .A3(new_n761_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n754_), .B1(new_n769_), .B2(new_n752_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n751_), .B1(new_n766_), .B2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n771_), .A2(new_n577_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n771_), .B2(new_n577_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n769_), .A2(new_n752_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT56), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n769_), .A2(new_n753_), .A3(new_n752_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n765_), .A2(new_n750_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n778_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT120), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT58), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n779_), .A2(new_n780_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n753_), .B1(new_n769_), .B2(new_n752_), .ZN(new_n786_));
  OAI211_X1 g585(.A(KEYINPUT120), .B(new_n784_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n783_), .A2(new_n274_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n299_), .B1(new_n776_), .B2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n301_), .A2(new_n324_), .A3(new_n568_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n790_), .B(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n530_), .B(new_n747_), .C1(new_n789_), .C2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(G113gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n795_), .A3(new_n569_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n793_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n775_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n771_), .A2(new_n577_), .A3(new_n773_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n787_), .A2(new_n274_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n784_), .B1(new_n781_), .B2(KEYINPUT120), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n300_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n790_), .B(KEYINPUT54), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n807_), .A2(KEYINPUT59), .A3(new_n530_), .A4(new_n747_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n568_), .B1(new_n798_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n796_), .B1(new_n809_), .B2(new_n795_), .ZN(G1340gat));
  INV_X1    g609(.A(new_n324_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT60), .ZN(new_n812_));
  INV_X1    g611(.A(G120gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n794_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n324_), .B1(new_n798_), .B2(new_n808_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n813_), .ZN(G1341gat));
  INV_X1    g617(.A(G127gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n794_), .A2(new_n819_), .A3(new_n299_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n300_), .B1(new_n798_), .B2(new_n808_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(new_n819_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT121), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n820_), .B(KEYINPUT121), .C1(new_n821_), .C2(new_n819_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1342gat));
  INV_X1    g625(.A(G134gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n794_), .A2(new_n827_), .A3(new_n578_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n273_), .B1(new_n798_), .B2(new_n808_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n827_), .ZN(G1343gat));
  INV_X1    g629(.A(new_n807_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n638_), .A2(new_n572_), .A3(new_n531_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT122), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n569_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n811_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g637(.A1(new_n834_), .A2(new_n299_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT61), .B(G155gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1346gat));
  NAND2_X1  g640(.A1(new_n834_), .A2(new_n578_), .ZN(new_n842_));
  INV_X1    g641(.A(G162gat), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n842_), .A2(KEYINPUT123), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT123), .B1(new_n842_), .B2(new_n843_), .ZN(new_n845_));
  NOR4_X1   g644(.A1(new_n831_), .A2(new_n843_), .A3(new_n625_), .A4(new_n833_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(G1347gat));
  NOR2_X1   g646(.A1(new_n638_), .A2(new_n572_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n807_), .A2(new_n530_), .A3(new_n569_), .A4(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n345_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n849_), .A2(new_n852_), .A3(G169gat), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(G169gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT62), .B1(new_n850_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n853_), .A2(new_n854_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n851_), .B1(new_n858_), .B2(new_n859_), .ZN(G1348gat));
  NAND3_X1  g659(.A1(new_n807_), .A2(new_n530_), .A3(new_n848_), .ZN(new_n861_));
  OR4_X1    g660(.A1(KEYINPUT125), .A2(new_n861_), .A3(G176gat), .A4(new_n324_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT125), .B(G176gat), .Z(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n861_), .B2(new_n324_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1349gat));
  OR2_X1    g664(.A1(new_n861_), .A2(new_n300_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G183gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n866_), .B2(new_n356_), .ZN(G1350gat));
  OAI21_X1  g667(.A(G190gat), .B1(new_n861_), .B2(new_n273_), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n577_), .A2(new_n357_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n861_), .B2(new_n870_), .ZN(G1351gat));
  NAND3_X1  g670(.A1(new_n807_), .A2(new_n531_), .A3(new_n848_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n568_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT126), .B(G197gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1352gat));
  INV_X1    g674(.A(new_n872_), .ZN(new_n876_));
  INV_X1    g675(.A(G204gat), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n876_), .B(new_n811_), .C1(KEYINPUT127), .C2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(KEYINPUT127), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1353gat));
  NOR2_X1   g679(.A1(new_n872_), .A2(new_n300_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  AND2_X1   g681(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n881_), .B2(new_n882_), .ZN(G1354gat));
  OAI21_X1  g684(.A(G218gat), .B1(new_n872_), .B2(new_n273_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n577_), .A2(G218gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n872_), .B2(new_n887_), .ZN(G1355gat));
endmodule


