//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NOR2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n205_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT8), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n208_), .B1(KEYINPUT9), .B2(new_n202_), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT10), .B(G99gat), .Z(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G92gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT9), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(G85gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n211_), .A2(new_n214_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n210_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G57gat), .B(G64gat), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n220_), .A2(KEYINPUT65), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(KEYINPUT65), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT11), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G71gat), .B(G78gat), .Z(new_n224_));
  OR2_X1    g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OR3_X1    g024(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT11), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n219_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n228_), .A2(KEYINPUT12), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n210_), .A2(new_n218_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n225_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(KEYINPUT12), .A3(new_n228_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n229_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G230gat), .A2(G233gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n228_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n235_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G120gat), .B(G148gat), .Z(new_n241_));
  XNOR2_X1  g040(.A(G176gat), .B(G204gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n240_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n236_), .A2(new_n239_), .A3(new_n245_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT13), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n247_), .A2(KEYINPUT13), .A3(new_n248_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G29gat), .B(G36gat), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n253_), .A2(KEYINPUT68), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(KEYINPUT68), .ZN(new_n255_));
  XOR2_X1   g054(.A(G43gat), .B(G50gat), .Z(new_n256_));
  OR3_X1    g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n256_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT15), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G15gat), .B(G22gat), .ZN(new_n261_));
  INV_X1    g060(.A(G1gat), .ZN(new_n262_));
  INV_X1    g061(.A(G8gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT14), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G1gat), .B(G8gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n260_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G229gat), .A2(G233gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n267_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n259_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n268_), .A2(new_n269_), .A3(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n259_), .B(new_n270_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n269_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G113gat), .B(G141gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G169gat), .B(G197gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n276_), .B(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n252_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT77), .ZN(new_n283_));
  INV_X1    g082(.A(G169gat), .ZN(new_n284_));
  INV_X1    g083(.A(G176gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n286_), .A2(KEYINPUT24), .A3(new_n287_), .A4(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT23), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT24), .B1(new_n286_), .B2(new_n287_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT26), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G183gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT25), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT25), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G183gat), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n300_), .A2(KEYINPUT76), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT76), .B1(new_n300_), .B2(new_n305_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n294_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT78), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n310_), .B1(G183gat), .B2(G190gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n290_), .A2(KEYINPUT23), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n309_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n290_), .A2(KEYINPUT23), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT78), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n295_), .A2(new_n296_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n316_), .B1(G183gat), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT22), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n320_));
  OAI21_X1  g119(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n308_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT30), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT80), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G227gat), .A2(G233gat), .ZN(new_n329_));
  INV_X1    g128(.A(G71gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G99gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(G15gat), .B(G43gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT79), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n332_), .B(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n328_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n326_), .A2(new_n327_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n328_), .A2(new_n335_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n336_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340_));
  INV_X1    g139(.A(G134gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G127gat), .ZN(new_n342_));
  INV_X1    g141(.A(G127gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G134gat), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n340_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n342_), .A2(new_n344_), .A3(new_n340_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G113gat), .B(G120gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n348_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n347_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n350_), .B1(new_n351_), .B2(new_n345_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT31), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT81), .B1(new_n354_), .B2(KEYINPUT83), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n339_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT83), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT81), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n339_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n356_), .B1(new_n359_), .B2(new_n354_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G197gat), .A2(G204gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT86), .B(G204gat), .ZN(new_n365_));
  INV_X1    g164(.A(G197gat), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT21), .ZN(new_n368_));
  INV_X1    g167(.A(G218gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(G211gat), .ZN(new_n370_));
  INV_X1    g169(.A(G211gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(G218gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n368_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT88), .B1(new_n367_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G204gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT86), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT86), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G204gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n366_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n373_), .A4(new_n364_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n375_), .A2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n368_), .B1(new_n380_), .B2(new_n363_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n370_), .A2(new_n372_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n377_), .A2(new_n379_), .A3(new_n366_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n368_), .B1(G197gat), .B2(G204gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n386_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n385_), .A2(KEYINPUT87), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT87), .B1(new_n385_), .B2(new_n389_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n384_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT20), .B1(new_n325_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n385_), .A2(new_n389_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n385_), .A2(KEYINPUT87), .A3(new_n389_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n396_), .A2(new_n397_), .B1(new_n375_), .B2(new_n383_), .ZN(new_n398_));
  INV_X1    g197(.A(G190gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n301_), .A2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n322_), .B1(new_n291_), .B2(new_n400_), .ZN(new_n401_));
  AND2_X1   g200(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n302_), .B(new_n304_), .C1(new_n402_), .C2(new_n298_), .ZN(new_n403_));
  OR3_X1    g202(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n289_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n401_), .B1(new_n405_), .B2(new_n316_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n398_), .A2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n362_), .B1(new_n393_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT90), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n396_), .A2(new_n397_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n410_), .A2(new_n384_), .A3(new_n324_), .A4(new_n308_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n406_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n392_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n413_), .A3(KEYINPUT20), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT90), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n362_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n409_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(new_n398_), .B2(new_n406_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n362_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n325_), .A2(new_n392_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(G8gat), .B(G36gat), .Z(new_n424_));
  XNOR2_X1  g223(.A(G64gat), .B(G92gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n426_), .B(new_n427_), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT32), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n417_), .A2(new_n423_), .A3(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(G155gat), .A2(G162gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT84), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G141gat), .A2(G148gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT3), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT3), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(G141gat), .B2(G148gat), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT2), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT85), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n441_), .B(KEYINPUT2), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n437_), .A2(new_n439_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n435_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n436_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n441_), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n434_), .B(KEYINPUT1), .Z(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n452_), .B2(new_n433_), .ZN(new_n453_));
  OAI211_X1 g252(.A(KEYINPUT92), .B(new_n353_), .C1(new_n449_), .C2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n435_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n446_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n455_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n349_), .A2(new_n352_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n453_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n454_), .A2(KEYINPUT4), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n458_), .A2(new_n460_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT4), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n463_), .A2(KEYINPUT92), .A3(new_n464_), .A4(new_n353_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G225gat), .A2(G233gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G29gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(G85gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT0), .B(G57gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n463_), .A2(new_n353_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n468_), .B1(new_n475_), .B2(new_n461_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n469_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n467_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n473_), .B1(new_n479_), .B2(new_n476_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  AND4_X1   g280(.A1(KEYINPUT20), .A2(new_n411_), .A3(new_n420_), .A4(new_n413_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n406_), .B(new_n384_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT20), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT94), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n483_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n421_), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n482_), .B1(new_n488_), .B2(new_n362_), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n431_), .B(new_n481_), .C1(new_n489_), .C2(new_n430_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT33), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n480_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n475_), .A2(new_n468_), .A3(new_n461_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n474_), .B(new_n493_), .C1(new_n466_), .C2(new_n468_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n494_), .A2(KEYINPUT93), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n480_), .A2(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(KEYINPUT93), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n492_), .A2(new_n495_), .A3(new_n496_), .A4(new_n497_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n414_), .A2(new_n415_), .A3(new_n362_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n415_), .B1(new_n414_), .B2(new_n362_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n423_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n428_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n423_), .B(new_n429_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n490_), .B1(new_n498_), .B2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT29), .B1(new_n449_), .B2(new_n453_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n392_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G228gat), .A2(G233gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n506_), .A2(new_n508_), .A3(new_n392_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G78gat), .B(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT89), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n449_), .A2(new_n453_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT29), .ZN(new_n518_));
  XOR2_X1   g317(.A(G22gat), .B(G50gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT28), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n517_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n520_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n506_), .A2(new_n508_), .A3(new_n392_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n508_), .B1(new_n506_), .B2(new_n392_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n512_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n516_), .A2(new_n523_), .B1(new_n514_), .B2(new_n526_), .ZN(new_n527_));
  AND4_X1   g326(.A1(KEYINPUT89), .A2(new_n526_), .A3(new_n514_), .A4(new_n523_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n505_), .A2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT95), .B1(new_n489_), .B2(new_n429_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT95), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n484_), .A2(new_n485_), .B1(new_n392_), .B2(new_n325_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n420_), .B1(new_n533_), .B2(new_n487_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n532_), .B(new_n428_), .C1(new_n534_), .C2(new_n482_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n531_), .A2(KEYINPUT27), .A3(new_n503_), .A4(new_n535_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n527_), .A2(new_n481_), .A3(new_n528_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT27), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n429_), .B1(new_n417_), .B2(new_n423_), .ZN(new_n540_));
  AOI211_X1 g339(.A(new_n428_), .B(new_n422_), .C1(new_n409_), .C2(new_n416_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n539_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT96), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n504_), .A2(KEYINPUT96), .A3(new_n539_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n538_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT97), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n530_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  AOI211_X1 g347(.A(KEYINPUT97), .B(new_n538_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n360_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT96), .B1(new_n504_), .B2(new_n539_), .ZN(new_n551_));
  AOI211_X1 g350(.A(new_n543_), .B(KEYINPUT27), .C1(new_n502_), .C2(new_n503_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n536_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT98), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(KEYINPUT98), .B(new_n536_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n360_), .A2(new_n481_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n555_), .A2(new_n529_), .A3(new_n556_), .A4(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n282_), .B1(new_n550_), .B2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(KEYINPUT67), .B(KEYINPUT34), .Z(new_n560_));
  NAND2_X1  g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n562_), .A2(KEYINPUT35), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n230_), .A2(new_n259_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n562_), .A2(KEYINPUT35), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT69), .Z(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(KEYINPUT70), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n260_), .A2(new_n219_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT70), .B1(new_n564_), .B2(new_n566_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n563_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n563_), .B(KEYINPUT72), .Z(new_n572_));
  NAND4_X1  g371(.A1(new_n568_), .A2(new_n564_), .A3(new_n566_), .A4(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT71), .ZN(new_n575_));
  XOR2_X1   g374(.A(G134gat), .B(G162gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n577_), .A2(KEYINPUT36), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n571_), .A2(new_n573_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n571_), .A2(new_n573_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n577_), .B(KEYINPUT36), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n580_), .B(KEYINPUT37), .C1(new_n581_), .C2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n231_), .B(new_n267_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587_));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT16), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G183gat), .B(G211gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  OR3_X1    g390(.A1(new_n586_), .A2(new_n587_), .A3(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(KEYINPUT17), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n586_), .A2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n571_), .A2(new_n573_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT73), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n582_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n571_), .A2(KEYINPUT73), .A3(new_n573_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n579_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n583_), .B(new_n595_), .C1(new_n600_), .C2(KEYINPUT37), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT74), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n559_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n262_), .A3(new_n481_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT38), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n600_), .B1(new_n550_), .B2(new_n558_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n595_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n282_), .A2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n481_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n605_), .A2(new_n606_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n607_), .A2(new_n614_), .A3(new_n615_), .ZN(G1324gat));
  NAND2_X1  g415(.A1(new_n555_), .A2(new_n556_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n611_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(G8gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT39), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n618_), .A2(new_n621_), .A3(G8gat), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n604_), .A2(new_n263_), .A3(new_n617_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n625_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1325gat));
  INV_X1    g428(.A(G15gat), .ZN(new_n630_));
  INV_X1    g429(.A(new_n360_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n611_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT41), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n630_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n633_), .B1(new_n603_), .B2(new_n634_), .ZN(G1326gat));
  OAI21_X1  g434(.A(G22gat), .B1(new_n612_), .B2(new_n529_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n529_), .A2(G22gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n603_), .B2(new_n639_), .ZN(G1327gat));
  NAND2_X1  g439(.A1(new_n609_), .A2(new_n600_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT102), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n559_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT103), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n559_), .A2(new_n645_), .A3(new_n642_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(G29gat), .B1(new_n647_), .B2(new_n481_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n282_), .A2(new_n595_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n583_), .B1(new_n600_), .B2(KEYINPUT37), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n650_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n550_), .A2(new_n558_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n655_), .B2(new_n651_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n651_), .ZN(new_n657_));
  AOI211_X1 g456(.A(new_n657_), .B(new_n653_), .C1(new_n550_), .C2(new_n558_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n649_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(KEYINPUT44), .B(new_n649_), .C1(new_n656_), .C2(new_n658_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n481_), .A2(G29gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n648_), .B1(new_n663_), .B2(new_n664_), .ZN(G1328gat));
  NAND3_X1  g464(.A1(new_n661_), .A2(new_n617_), .A3(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G36gat), .ZN(new_n667_));
  INV_X1    g466(.A(new_n617_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(G36gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n644_), .A2(new_n646_), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT45), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT45), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n644_), .A2(new_n672_), .A3(new_n646_), .A4(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n667_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n667_), .A2(KEYINPUT46), .A3(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1329gat));
  NAND4_X1  g478(.A1(new_n661_), .A2(G43gat), .A3(new_n631_), .A4(new_n662_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n644_), .A2(new_n631_), .A3(new_n646_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT104), .B(G43gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g484(.A(G50gat), .ZN(new_n686_));
  INV_X1    g485(.A(new_n529_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n647_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n661_), .A2(new_n687_), .A3(new_n662_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n689_), .A2(new_n690_), .A3(G50gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n689_), .B2(G50gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(G1331gat));
  INV_X1    g492(.A(new_n251_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(new_n249_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n280_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n655_), .A2(new_n602_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G57gat), .B1(new_n698_), .B2(new_n481_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n608_), .A2(new_n595_), .A3(new_n697_), .ZN(new_n700_));
  INV_X1    g499(.A(G57gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n481_), .B2(KEYINPUT106), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(KEYINPUT106), .B2(new_n701_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n699_), .B1(new_n700_), .B2(new_n703_), .ZN(G1332gat));
  INV_X1    g503(.A(G64gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n700_), .B2(new_n617_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT48), .Z(new_n707_));
  NAND3_X1  g506(.A1(new_n698_), .A2(new_n705_), .A3(new_n617_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1333gat));
  AOI21_X1  g508(.A(new_n330_), .B1(new_n700_), .B2(new_n631_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT49), .Z(new_n711_));
  NAND3_X1  g510(.A1(new_n698_), .A2(new_n330_), .A3(new_n631_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1334gat));
  INV_X1    g512(.A(G78gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n700_), .B2(new_n687_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT50), .Z(new_n716_));
  NAND3_X1  g515(.A1(new_n698_), .A2(new_n714_), .A3(new_n687_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1335gat));
  NOR3_X1   g517(.A1(new_n695_), .A2(new_n595_), .A3(new_n696_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G85gat), .B1(new_n720_), .B2(new_n613_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n655_), .A2(new_n642_), .A3(new_n697_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT107), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n655_), .A2(new_n642_), .A3(new_n724_), .A4(new_n697_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n613_), .A2(G85gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n721_), .B1(new_n726_), .B2(new_n727_), .ZN(G1336gat));
  NAND2_X1  g527(.A1(new_n723_), .A2(new_n725_), .ZN(new_n729_));
  AOI21_X1  g528(.A(G92gat), .B1(new_n729_), .B2(new_n617_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n720_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n617_), .A2(new_n215_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n730_), .B1(new_n731_), .B2(new_n732_), .ZN(G1337gat));
  NAND2_X1  g532(.A1(new_n631_), .A2(new_n212_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT108), .B1(new_n726_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n631_), .B(new_n719_), .C1(new_n656_), .C2(new_n658_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G99gat), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n729_), .A2(new_n739_), .A3(new_n212_), .A4(new_n631_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n735_), .A2(new_n738_), .A3(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR2_X1   g541(.A1(new_n529_), .A2(G106gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT110), .B1(new_n729_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745_));
  INV_X1    g544(.A(new_n743_), .ZN(new_n746_));
  AOI211_X1 g545(.A(new_n745_), .B(new_n746_), .C1(new_n723_), .C2(new_n725_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n744_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n687_), .B(new_n719_), .C1(new_n656_), .C2(new_n658_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(G106gat), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n749_), .A2(new_n751_), .A3(new_n754_), .A4(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n755_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n751_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(new_n748_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n759_), .ZN(G1339gat));
  NOR2_X1   g559(.A1(new_n252_), .A2(new_n696_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n657_), .A2(new_n761_), .A3(new_n595_), .A4(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n695_), .A2(new_n280_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n762_), .B1(new_n765_), .B2(new_n601_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n247_), .A2(new_n248_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n272_), .A2(new_n275_), .A3(new_n279_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n268_), .A2(new_n271_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n268_), .A2(KEYINPUT114), .A3(new_n271_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n274_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n279_), .B1(new_n273_), .B2(new_n269_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n769_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n768_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n229_), .A2(new_n233_), .A3(new_n238_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n236_), .A2(KEYINPUT55), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n238_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n245_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT113), .B1(new_n779_), .B2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n696_), .B(new_n248_), .C1(new_n783_), .C2(KEYINPUT56), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n783_), .A2(KEYINPUT56), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n777_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n600_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(KEYINPUT57), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT58), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n776_), .A2(new_n793_), .A3(new_n248_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n776_), .B2(new_n248_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n779_), .A2(new_n782_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT56), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n779_), .A2(new_n800_), .A3(new_n782_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n792_), .B1(new_n797_), .B2(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n799_), .A2(new_n801_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n804_), .B(KEYINPUT58), .C1(new_n796_), .C2(new_n795_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n805_), .A3(new_n651_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n790_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n786_), .A2(new_n787_), .A3(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n791_), .A2(new_n806_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n767_), .B1(new_n809_), .B2(new_n609_), .ZN(new_n810_));
  NOR4_X1   g609(.A1(new_n617_), .A2(new_n687_), .A3(new_n613_), .A4(new_n360_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(G113gat), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n696_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n809_), .A2(new_n609_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n767_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT59), .B1(new_n819_), .B2(new_n811_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n810_), .A2(new_n821_), .A3(new_n812_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n816_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n819_), .A2(KEYINPUT59), .A3(new_n811_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n821_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n825_), .A3(KEYINPUT117), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n280_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n815_), .B1(new_n827_), .B2(new_n814_), .ZN(G1340gat));
  INV_X1    g627(.A(G120gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n695_), .B2(KEYINPUT60), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n813_), .B(new_n830_), .C1(KEYINPUT60), .C2(new_n829_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n695_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n829_), .ZN(G1341gat));
  NAND3_X1  g632(.A1(new_n813_), .A2(new_n343_), .A3(new_n595_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n609_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n343_), .ZN(G1342gat));
  NOR2_X1   g635(.A1(new_n657_), .A2(new_n341_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n839_));
  AOI21_X1  g638(.A(G134gat), .B1(new_n813_), .B2(new_n600_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT118), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n824_), .A2(new_n825_), .A3(KEYINPUT117), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT117), .B1(new_n824_), .B2(new_n825_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n837_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845_));
  INV_X1    g644(.A(new_n840_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n841_), .A2(new_n847_), .ZN(G1343gat));
  NOR3_X1   g647(.A1(new_n631_), .A2(new_n529_), .A3(new_n613_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n668_), .A2(new_n849_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT119), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n819_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n819_), .A2(new_n851_), .A3(KEYINPUT120), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n696_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n252_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT121), .B(G148gat), .Z(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1345gat));
  NAND2_X1  g660(.A1(new_n856_), .A2(new_n595_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT61), .B(G155gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  AND2_X1   g663(.A1(new_n854_), .A2(new_n855_), .ZN(new_n865_));
  INV_X1    g664(.A(G162gat), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n657_), .ZN(new_n867_));
  OAI211_X1 g666(.A(KEYINPUT122), .B(new_n866_), .C1(new_n865_), .C2(new_n787_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n787_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(G162gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n867_), .B1(new_n868_), .B2(new_n871_), .ZN(G1347gat));
  XOR2_X1   g671(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n873_));
  NAND3_X1  g672(.A1(new_n617_), .A2(new_n529_), .A3(new_n557_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n810_), .A2(new_n280_), .A3(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n875_), .B2(new_n319_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(G169gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n284_), .B1(new_n875_), .B2(new_n873_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n876_), .B2(new_n878_), .ZN(G1348gat));
  NOR2_X1   g678(.A1(new_n810_), .A2(new_n874_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n252_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n595_), .ZN(new_n883_));
  OR3_X1    g682(.A1(new_n883_), .A2(KEYINPUT124), .A3(new_n305_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT124), .B1(new_n883_), .B2(new_n305_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n301_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(G1350gat));
  OAI211_X1 g686(.A(new_n880_), .B(new_n600_), .C1(new_n298_), .C2(new_n402_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n810_), .A2(new_n657_), .A3(new_n874_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n399_), .ZN(G1351gat));
  NAND3_X1  g689(.A1(new_n617_), .A2(new_n360_), .A3(new_n537_), .ZN(new_n891_));
  NOR4_X1   g690(.A1(new_n810_), .A2(new_n366_), .A3(new_n280_), .A4(new_n891_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n892_), .A2(KEYINPUT125), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(KEYINPUT125), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n810_), .A2(new_n891_), .ZN(new_n895_));
  AOI21_X1  g694(.A(G197gat), .B1(new_n895_), .B2(new_n696_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n893_), .A2(new_n894_), .A3(new_n896_), .ZN(G1352gat));
  NAND3_X1  g696(.A1(new_n895_), .A2(new_n365_), .A3(new_n252_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n898_), .A2(new_n899_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n895_), .A2(new_n252_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G204gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n901_), .B2(new_n903_), .ZN(G1353gat));
  INV_X1    g703(.A(KEYINPUT63), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n595_), .B1(new_n905_), .B2(new_n371_), .ZN(new_n906_));
  XOR2_X1   g705(.A(new_n906_), .B(KEYINPUT127), .Z(new_n907_));
  NAND2_X1  g706(.A1(new_n895_), .A2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n905_), .A2(new_n371_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1354gat));
  NAND3_X1  g709(.A1(new_n895_), .A2(new_n369_), .A3(new_n600_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n810_), .A2(new_n657_), .A3(new_n891_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n369_), .ZN(G1355gat));
endmodule


