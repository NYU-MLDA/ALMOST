//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n952_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT86), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n203_), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT85), .B(G15gat), .Z(new_n208_));
  NAND2_X1  g007(.A1(G227gat), .A2(G233gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT84), .B(G43gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n207_), .B(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT31), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT81), .ZN(new_n217_));
  INV_X1    g016(.A(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n217_), .A2(KEYINPUT24), .A3(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n223_), .A2(KEYINPUT23), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n220_), .A2(KEYINPUT24), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n221_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT26), .B(G190gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT79), .ZN(new_n231_));
  INV_X1    g030(.A(G183gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT25), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n232_), .A2(KEYINPUT25), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n230_), .B(new_n233_), .C1(new_n234_), .C2(new_n231_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT80), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n229_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT22), .B(G169gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n219_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n217_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT23), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n223_), .A2(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(G183gat), .A2(G190gat), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n242_), .B(new_n243_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n240_), .B1(KEYINPUT83), .B2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n245_), .B1(KEYINPUT83), .B2(new_n244_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n237_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT30), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G71gat), .B(G99gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n250_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n215_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n253_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n255_), .A2(KEYINPUT31), .A3(new_n251_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n214_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT31), .B1(new_n255_), .B2(new_n251_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n252_), .A2(new_n253_), .A3(new_n215_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n213_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT102), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G8gat), .B(G36gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT18), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G64gat), .B(G92gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT19), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n216_), .A2(KEYINPUT24), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n270_), .A2(KEYINPUT94), .B1(new_n218_), .B2(new_n219_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n216_), .A2(KEYINPUT24), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT94), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT25), .B(G183gat), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n271_), .A2(new_n274_), .B1(new_n230_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n242_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(new_n228_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT95), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n277_), .A2(KEYINPUT95), .A3(new_n228_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n276_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G197gat), .B(G204gat), .Z(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT21), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G197gat), .B(G204gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT21), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  OR3_X1    g088(.A1(new_n285_), .A2(new_n288_), .A3(new_n286_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT92), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n240_), .A2(KEYINPUT96), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n243_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT96), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n239_), .A2(new_n217_), .A3(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n289_), .A2(new_n290_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT92), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n282_), .A2(new_n293_), .A3(new_n298_), .A4(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT100), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n302_), .A3(KEYINPUT20), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n247_), .A2(new_n299_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n302_), .B1(new_n301_), .B2(KEYINPUT20), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n269_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT20), .B1(new_n247_), .B2(new_n299_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT97), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n298_), .A2(new_n309_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n294_), .A2(new_n295_), .A3(KEYINPUT97), .A4(new_n297_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n291_), .B1(new_n312_), .B2(new_n282_), .ZN(new_n313_));
  OR3_X1    g112(.A1(new_n308_), .A2(new_n313_), .A3(new_n269_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n267_), .B1(new_n307_), .B2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n269_), .B1(new_n308_), .B2(new_n313_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n291_), .A3(new_n282_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n269_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n317_), .A2(new_n304_), .A3(KEYINPUT20), .A4(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n316_), .A2(new_n267_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT27), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n315_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT101), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n316_), .A2(new_n319_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n267_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n320_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT27), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n324_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n316_), .A2(new_n267_), .A3(new_n319_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n267_), .B1(new_n316_), .B2(new_n319_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n324_), .B(new_n329_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n323_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G155gat), .B(G162gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT90), .ZN(new_n337_));
  NOR2_X1   g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n338_), .A2(KEYINPUT3), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(KEYINPUT3), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n339_), .A2(new_n340_), .B1(new_n342_), .B2(KEYINPUT2), .ZN(new_n343_));
  XOR2_X1   g142(.A(KEYINPUT87), .B(KEYINPUT2), .Z(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT88), .B1(new_n344_), .B2(new_n341_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT87), .B(KEYINPUT2), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT88), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n342_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n343_), .B1(new_n345_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n337_), .B1(new_n349_), .B2(KEYINPUT89), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT89), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n344_), .A2(KEYINPUT88), .A3(new_n341_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n347_), .B1(new_n346_), .B2(new_n342_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n351_), .B1(new_n354_), .B2(new_n343_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n350_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT28), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358_));
  NOR2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n359_), .B1(KEYINPUT1), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(KEYINPUT1), .B2(new_n360_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n338_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n341_), .A3(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .A4(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n364_), .B1(new_n350_), .B2(new_n355_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT28), .B1(new_n366_), .B2(KEYINPUT29), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G22gat), .B(G50gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n368_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT93), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT93), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n369_), .ZN(new_n375_));
  INV_X1    g174(.A(G233gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT91), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n377_), .A2(G228gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(G228gat), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n376_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n366_), .A2(KEYINPUT29), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n293_), .A2(new_n300_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n381_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G78gat), .B(G106gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n381_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(new_n299_), .A3(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n387_), .B1(new_n385_), .B2(new_n389_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n372_), .B(new_n375_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n392_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n374_), .B1(new_n373_), .B2(new_n369_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n390_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G1gat), .B(G29gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(G57gat), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(KEYINPUT98), .B(KEYINPUT0), .Z(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT4), .B1(new_n366_), .B2(new_n207_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n366_), .A2(new_n207_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n204_), .A2(new_n206_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n364_), .B(new_n404_), .C1(new_n350_), .C2(new_n355_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n402_), .B1(new_n406_), .B2(KEYINPUT4), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n401_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n411_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n401_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n393_), .A2(new_n396_), .A3(new_n414_), .A4(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n263_), .B1(new_n335_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n329_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT101), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n322_), .B1(new_n420_), .B2(new_n333_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n393_), .A2(new_n396_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n416_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(new_n413_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n421_), .A2(new_n422_), .A3(KEYINPUT102), .A4(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n418_), .A2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT99), .B1(new_n413_), .B2(KEYINPUT33), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n403_), .A2(new_n405_), .A3(new_n409_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n401_), .B(new_n428_), .C1(new_n407_), .C2(new_n409_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n429_), .A2(new_n320_), .A3(new_n327_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT99), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n431_), .B(new_n432_), .C1(new_n415_), .C2(new_n401_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n413_), .A2(KEYINPUT33), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n427_), .A2(new_n430_), .A3(new_n433_), .A4(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n307_), .A2(new_n314_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(KEYINPUT32), .A3(new_n267_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n267_), .A2(KEYINPUT32), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n316_), .A2(new_n319_), .A3(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n437_), .B(new_n439_), .C1(new_n423_), .C2(new_n413_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n422_), .B1(new_n435_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n262_), .B1(new_n426_), .B2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n335_), .A2(new_n422_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n261_), .A2(new_n424_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G229gat), .A2(G233gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G29gat), .B(G36gat), .Z(new_n450_));
  XOR2_X1   g249(.A(G43gat), .B(G50gat), .Z(new_n451_));
  XOR2_X1   g250(.A(new_n450_), .B(new_n451_), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT76), .ZN(new_n453_));
  INV_X1    g252(.A(G1gat), .ZN(new_n454_));
  INV_X1    g253(.A(G8gat), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT14), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT73), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT73), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n458_), .B(KEYINPUT14), .C1(new_n454_), .C2(new_n455_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G15gat), .B(G22gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT74), .ZN(new_n462_));
  XOR2_X1   g261(.A(G1gat), .B(G8gat), .Z(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n462_), .A2(new_n464_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n453_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n453_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n449_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n465_), .A2(new_n466_), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n452_), .B(KEYINPUT15), .Z(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n467_), .A3(new_n448_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G113gat), .B(G141gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT77), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G169gat), .B(G197gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n470_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT78), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n470_), .A2(KEYINPUT78), .A3(new_n474_), .A4(new_n478_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n470_), .A2(new_n474_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n478_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n447_), .A2(KEYINPUT103), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT103), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n435_), .A2(new_n440_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n418_), .B(new_n425_), .C1(new_n490_), .C2(new_n422_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n445_), .B1(new_n491_), .B2(new_n262_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n487_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n489_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n488_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G230gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(KEYINPUT10), .B(G99gat), .Z(new_n498_));
  INV_X1    g297(.A(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G85gat), .B(G92gat), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT9), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT6), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(G99gat), .A3(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(G85gat), .ZN(new_n508_));
  INV_X1    g307(.A(G92gat), .ZN(new_n509_));
  OR3_X1    g308(.A1(new_n508_), .A2(new_n509_), .A3(KEYINPUT9), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n500_), .A2(new_n502_), .A3(new_n507_), .A4(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(G99gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(new_n499_), .A3(KEYINPUT64), .ZN(new_n514_));
  NOR3_X1   g313(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n515_));
  OAI211_X1 g314(.A(KEYINPUT7), .B(new_n514_), .C1(new_n515_), .C2(KEYINPUT64), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT65), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(new_n513_), .A3(new_n499_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT64), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT7), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n507_), .A2(KEYINPUT66), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT66), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n504_), .A2(new_n506_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n501_), .B1(new_n522_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT8), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n514_), .A2(KEYINPUT7), .ZN(new_n529_));
  NOR2_X1   g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT64), .B1(new_n530_), .B2(new_n517_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n521_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n507_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n501_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(KEYINPUT8), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n512_), .B1(new_n528_), .B2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G57gat), .B(G64gat), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n538_), .A2(KEYINPUT11), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(KEYINPUT11), .ZN(new_n540_));
  XOR2_X1   g339(.A(G71gat), .B(G78gat), .Z(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n540_), .A2(new_n541_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n537_), .A2(KEYINPUT67), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT8), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n532_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n547_), .B2(new_n501_), .ZN(new_n548_));
  AOI211_X1 g347(.A(KEYINPUT8), .B(new_n534_), .C1(new_n532_), .C2(new_n507_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n511_), .B(new_n544_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT67), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n545_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n537_), .A2(new_n544_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n497_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n550_), .A2(new_n496_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT12), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n511_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n544_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n504_), .A2(new_n506_), .A3(new_n524_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n524_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n534_), .B1(new_n563_), .B2(new_n532_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n536_), .B1(new_n564_), .B2(new_n546_), .ZN(new_n565_));
  AOI211_X1 g364(.A(KEYINPUT12), .B(new_n544_), .C1(new_n565_), .C2(new_n511_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n556_), .B1(new_n560_), .B2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G120gat), .B(G148gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT5), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G176gat), .B(G204gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n555_), .A2(new_n567_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n572_), .B1(new_n555_), .B2(new_n567_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n576_), .A2(KEYINPUT13), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(KEYINPUT13), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT68), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT37), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n558_), .A2(new_n452_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT70), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT34), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n472_), .B2(new_n558_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT69), .Z(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n584_), .A2(new_n588_), .A3(new_n591_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(KEYINPUT72), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT36), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT71), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n598_), .B(new_n599_), .Z(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n595_), .A2(new_n596_), .A3(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n593_), .A2(new_n600_), .A3(new_n594_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n596_), .B1(new_n595_), .B2(new_n601_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n582_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n595_), .A2(new_n601_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT36), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n608_), .A2(KEYINPUT37), .A3(new_n603_), .A4(new_n602_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n544_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n471_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT17), .ZN(new_n614_));
  XOR2_X1   g413(.A(G127gat), .B(G155gat), .Z(new_n615_));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n613_), .A2(new_n614_), .A3(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(KEYINPUT17), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n620_), .B1(new_n613_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n610_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n581_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n495_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT104), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n424_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n495_), .A2(KEYINPUT104), .A3(new_n624_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n627_), .A2(new_n454_), .A3(new_n628_), .A4(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n604_), .A2(new_n605_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n492_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n579_), .A2(new_n493_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n622_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G1gat), .B1(new_n639_), .B2(new_n424_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n630_), .A2(new_n631_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n632_), .A2(new_n640_), .A3(new_n641_), .ZN(G1324gat));
  XNOR2_X1  g441(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n447_), .A2(new_n335_), .A3(new_n633_), .A4(new_n638_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n644_), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT105), .B1(new_n644_), .B2(G8gat), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT106), .B(KEYINPUT39), .Z(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n645_), .A2(new_n646_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n653_));
  NOR4_X1   g452(.A1(new_n492_), .A2(new_n421_), .A3(new_n634_), .A4(new_n637_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n653_), .B1(new_n654_), .B2(new_n455_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n644_), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n649_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n421_), .A2(G8gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n627_), .A2(new_n629_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n643_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n650_), .B(new_n651_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n655_), .A2(new_n656_), .A3(new_n647_), .ZN(new_n663_));
  AND4_X1   g462(.A1(new_n660_), .A2(new_n662_), .A3(new_n663_), .A4(new_n643_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n661_), .A2(new_n664_), .ZN(G1325gat));
  OAI21_X1  g464(.A(G15gat), .B1(new_n639_), .B2(new_n262_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT41), .Z(new_n667_));
  NOR2_X1   g466(.A1(new_n262_), .A2(G15gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n627_), .A2(new_n629_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1326gat));
  INV_X1    g469(.A(new_n422_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(G22gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n627_), .A2(new_n629_), .A3(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n635_), .A2(new_n422_), .A3(new_n638_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(G22gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT108), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n674_), .A2(new_n677_), .A3(G22gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n676_), .A2(KEYINPUT42), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n673_), .A2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT42), .B1(new_n676_), .B2(new_n678_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1327gat));
  INV_X1    g481(.A(new_n579_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n622_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n634_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n488_), .B2(new_n494_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G29gat), .B1(new_n686_), .B2(new_n628_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT109), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n610_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n606_), .A2(new_n609_), .A3(KEYINPUT109), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT43), .B1(new_n492_), .B2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n610_), .A2(KEYINPUT43), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n447_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n636_), .A2(new_n684_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT44), .B1(new_n695_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  AOI211_X1 g498(.A(new_n699_), .B(new_n696_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n628_), .A2(G29gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n687_), .B1(new_n701_), .B2(new_n702_), .ZN(G1328gat));
  NOR2_X1   g502(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n704_));
  INV_X1    g503(.A(G36gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n701_), .B2(new_n335_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n421_), .A2(G36gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n686_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n707_), .B1(new_n686_), .B2(new_n708_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n704_), .B1(new_n706_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n711_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n709_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n704_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n698_), .A2(new_n700_), .A3(new_n421_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n715_), .B(new_n716_), .C1(new_n717_), .C2(new_n705_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n713_), .A2(new_n718_), .ZN(G1329gat));
  INV_X1    g518(.A(G43gat), .ZN(new_n720_));
  NOR4_X1   g519(.A1(new_n698_), .A2(new_n700_), .A3(new_n720_), .A4(new_n262_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G43gat), .B1(new_n686_), .B2(new_n261_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT47), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n262_), .A2(new_n720_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n701_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n723_), .A2(new_n727_), .ZN(G1330gat));
  NOR3_X1   g527(.A1(new_n698_), .A2(new_n700_), .A3(new_n671_), .ZN(new_n729_));
  INV_X1    g528(.A(G50gat), .ZN(new_n730_));
  INV_X1    g529(.A(new_n686_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n422_), .A2(new_n730_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT111), .ZN(new_n733_));
  OAI22_X1  g532(.A1(new_n729_), .A2(new_n730_), .B1(new_n731_), .B2(new_n733_), .ZN(G1331gat));
  NAND3_X1  g533(.A1(new_n447_), .A2(KEYINPUT112), .A3(new_n493_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(new_n492_), .B2(new_n487_), .ZN(new_n737_));
  AOI211_X1 g536(.A(new_n683_), .B(new_n623_), .C1(new_n735_), .C2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G57gat), .B1(new_n738_), .B2(new_n628_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n580_), .A2(new_n487_), .A3(new_n684_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n635_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n424_), .A2(KEYINPUT113), .ZN(new_n743_));
  MUX2_X1   g542(.A(KEYINPUT113), .B(new_n743_), .S(G57gat), .Z(new_n744_));
  AOI21_X1  g543(.A(new_n739_), .B1(new_n742_), .B2(new_n744_), .ZN(G1332gat));
  OAI21_X1  g544(.A(G64gat), .B1(new_n741_), .B2(new_n421_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT48), .ZN(new_n747_));
  INV_X1    g546(.A(G64gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n738_), .A2(new_n748_), .A3(new_n335_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1333gat));
  OAI21_X1  g549(.A(G71gat), .B1(new_n741_), .B2(new_n262_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT49), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n262_), .A2(G71gat), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT114), .Z(new_n754_));
  NAND2_X1  g553(.A1(new_n738_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(G1334gat));
  INV_X1    g555(.A(G78gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n738_), .A2(new_n757_), .A3(new_n422_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G78gat), .B1(new_n741_), .B2(new_n671_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(KEYINPUT50), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(KEYINPUT50), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n758_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT115), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n487_), .A2(new_n622_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n692_), .A2(KEYINPUT116), .A3(new_n694_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT116), .B1(new_n692_), .B2(new_n694_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n579_), .B(new_n764_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768_), .B2(new_n424_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n581_), .A2(new_n684_), .A3(new_n634_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(new_n508_), .A3(new_n628_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n769_), .A2(new_n772_), .ZN(G1336gat));
  OAI21_X1  g572(.A(G92gat), .B1(new_n768_), .B2(new_n421_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n509_), .A3(new_n335_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1337gat));
  AND2_X1   g575(.A1(new_n261_), .A2(new_n498_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n771_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n778_), .B(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n579_), .A2(new_n764_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n695_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n781_), .B1(new_n783_), .B2(new_n765_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n513_), .B1(new_n784_), .B2(new_n261_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT51), .B1(new_n780_), .B2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G99gat), .B1(new_n768_), .B2(new_n262_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n778_), .B(KEYINPUT117), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n787_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n786_), .A2(new_n790_), .ZN(G1338gat));
  NAND3_X1  g590(.A1(new_n771_), .A2(new_n499_), .A3(new_n422_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n781_), .A2(new_n671_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n499_), .B1(new_n695_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n794_), .A2(new_n795_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n792_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT53), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n800_), .B(new_n792_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1339gat));
  NAND4_X1  g601(.A1(new_n610_), .A2(new_n493_), .A3(new_n683_), .A4(new_n622_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n610_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n448_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n485_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n468_), .A2(new_n448_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n809_), .A2(new_n810_), .B1(new_n473_), .B2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n808_), .A2(KEYINPUT119), .A3(new_n485_), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n812_), .A2(new_n813_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n807_), .B1(new_n814_), .B2(new_n573_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n809_), .A2(new_n810_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n811_), .A2(new_n473_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n813_), .A3(new_n817_), .ZN(new_n818_));
  AND4_X1   g617(.A1(new_n807_), .A2(new_n483_), .A3(new_n818_), .A4(new_n573_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n815_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n552_), .B(new_n545_), .C1(new_n560_), .C2(new_n566_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n497_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT12), .B1(new_n537_), .B2(new_n544_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n558_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n824_), .B1(new_n827_), .B2(new_n556_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n556_), .B(new_n824_), .C1(new_n560_), .C2(new_n566_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n823_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT118), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n567_), .A2(KEYINPUT55), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n829_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(new_n823_), .ZN(new_n836_));
  AOI211_X1 g635(.A(new_n821_), .B(new_n572_), .C1(new_n832_), .C2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n838_));
  AOI221_X4 g637(.A(KEYINPUT118), .B1(new_n822_), .B2(new_n497_), .C1(new_n833_), .C2(new_n829_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n835_), .B1(new_n834_), .B2(new_n823_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n571_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n821_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n837_), .B1(new_n838_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n841_), .A2(KEYINPUT121), .A3(new_n821_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n820_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT122), .B(new_n806_), .C1(new_n845_), .C2(KEYINPUT58), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n572_), .B1(new_n832_), .B2(new_n836_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n838_), .B1(new_n848_), .B2(KEYINPUT56), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(KEYINPUT56), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n844_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n818_), .A2(new_n483_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT120), .B1(new_n852_), .B2(new_n574_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n814_), .A2(new_n807_), .A3(new_n573_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT58), .B1(new_n851_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n847_), .B1(new_n856_), .B2(new_n610_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n845_), .A2(KEYINPUT58), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n846_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n487_), .A2(new_n573_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n850_), .B2(new_n842_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n852_), .A2(new_n576_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n633_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT57), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n859_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n805_), .B1(new_n865_), .B2(new_n684_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NOR4_X1   g666(.A1(new_n262_), .A2(new_n335_), .A3(new_n422_), .A4(new_n424_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(KEYINPUT123), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n622_), .B1(new_n859_), .B2(new_n864_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n870_), .B2(new_n805_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n869_), .A2(new_n487_), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(G113gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n867_), .A2(KEYINPUT59), .A3(new_n868_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n871_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n875_), .B1(new_n487_), .B2(KEYINPUT124), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(KEYINPUT124), .B2(new_n875_), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n874_), .A2(new_n875_), .B1(new_n879_), .B2(new_n881_), .ZN(G1340gat));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n883_), .A2(KEYINPUT60), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n683_), .B2(KEYINPUT60), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n869_), .A2(new_n873_), .A3(new_n884_), .A4(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n580_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n883_), .ZN(G1341gat));
  INV_X1    g687(.A(G127gat), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n869_), .A2(new_n889_), .A3(new_n622_), .A4(new_n873_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n684_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n889_), .ZN(G1342gat));
  INV_X1    g691(.A(G134gat), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n869_), .A2(new_n893_), .A3(new_n634_), .A4(new_n873_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n610_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n893_), .ZN(G1343gat));
  NOR4_X1   g695(.A1(new_n671_), .A2(new_n335_), .A3(new_n261_), .A4(new_n424_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n867_), .A2(new_n487_), .A3(new_n897_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT125), .B(G141gat), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1344gat));
  NAND3_X1  g699(.A1(new_n867_), .A2(new_n581_), .A3(new_n897_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g701(.A1(new_n867_), .A2(new_n622_), .A3(new_n897_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G155gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  AND2_X1   g704(.A1(new_n867_), .A2(new_n897_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n634_), .ZN(new_n907_));
  INV_X1    g706(.A(G162gat), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n691_), .A2(new_n908_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n907_), .A2(new_n908_), .B1(new_n906_), .B2(new_n909_), .ZN(G1347gat));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n262_), .A2(new_n421_), .A3(new_n628_), .A4(new_n422_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n487_), .ZN(new_n913_));
  OAI211_X1 g712(.A(KEYINPUT62), .B(G169gat), .C1(new_n866_), .C2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n913_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n238_), .B(new_n915_), .C1(new_n870_), .C2(new_n805_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n870_), .B2(new_n805_), .ZN(new_n918_));
  AOI21_X1  g717(.A(KEYINPUT62), .B1(new_n918_), .B2(G169gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n911_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(G169gat), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n923_), .A2(KEYINPUT126), .A3(new_n916_), .A4(new_n914_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n920_), .A2(new_n924_), .ZN(G1348gat));
  NAND2_X1  g724(.A1(new_n867_), .A2(new_n912_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G176gat), .B1(new_n926_), .B2(new_n580_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n579_), .A2(new_n219_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(G1349gat));
  NOR3_X1   g728(.A1(new_n926_), .A2(new_n275_), .A3(new_n684_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n926_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n622_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n930_), .B1(new_n232_), .B2(new_n932_), .ZN(G1350gat));
  OAI21_X1  g732(.A(G190gat), .B1(new_n926_), .B2(new_n610_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n634_), .A2(new_n230_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n926_), .B2(new_n935_), .ZN(G1351gat));
  NOR3_X1   g735(.A1(new_n421_), .A2(new_n261_), .A3(new_n417_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n867_), .A2(new_n487_), .A3(new_n937_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g738(.A1(new_n867_), .A2(new_n581_), .A3(new_n937_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g740(.A1(new_n867_), .A2(new_n937_), .ZN(new_n942_));
  XOR2_X1   g741(.A(KEYINPUT63), .B(G211gat), .Z(new_n943_));
  NAND3_X1  g742(.A1(new_n942_), .A2(new_n622_), .A3(new_n943_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n867_), .A2(new_n937_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n946_), .B2(new_n684_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n944_), .A2(new_n947_), .ZN(G1354gat));
  NAND2_X1  g747(.A1(new_n942_), .A2(new_n634_), .ZN(new_n949_));
  INV_X1    g748(.A(G218gat), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n806_), .A2(G218gat), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(KEYINPUT127), .ZN(new_n952_));
  AOI22_X1  g751(.A1(new_n949_), .A2(new_n950_), .B1(new_n942_), .B2(new_n952_), .ZN(G1355gat));
endmodule


