//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_;
  AND2_X1   g000(.A1(G71gat), .A2(G78gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G57gat), .B(G64gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n204_), .B1(new_n205_), .B2(KEYINPUT11), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(new_n205_), .B2(KEYINPUT11), .ZN(new_n208_));
  INV_X1    g007(.A(G64gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G57gat), .ZN(new_n210_));
  INV_X1    g009(.A(G57gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G64gat), .ZN(new_n212_));
  AND4_X1   g011(.A1(new_n207_), .A2(new_n210_), .A3(new_n212_), .A4(KEYINPUT11), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n206_), .B1(new_n208_), .B2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(new_n212_), .A3(KEYINPUT11), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT67), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n210_), .A2(new_n212_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n210_), .A2(new_n212_), .A3(new_n207_), .A4(KEYINPUT11), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n216_), .A2(new_n219_), .A3(new_n204_), .A4(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n214_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT69), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G99gat), .A2(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT6), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT6), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  OR3_X1    g028(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G85gat), .ZN(new_n232_));
  INV_X1    g031(.A(G92gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G85gat), .A2(G92gat), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT8), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT8), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n231_), .A2(new_n239_), .A3(new_n236_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT66), .B(G106gat), .ZN(new_n241_));
  OR2_X1    g040(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n242_), .A2(KEYINPUT65), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT65), .B1(new_n242_), .B2(new_n243_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n241_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n234_), .A2(KEYINPUT9), .A3(new_n235_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n235_), .A2(KEYINPUT9), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n228_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n238_), .A2(new_n240_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT12), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n223_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G230gat), .A2(G233gat), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n254_), .B(KEYINPUT64), .Z(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(new_n250_), .B2(new_n222_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n246_), .A2(new_n249_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n231_), .A2(new_n239_), .A3(new_n236_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n239_), .B1(new_n231_), .B2(new_n236_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n214_), .A2(new_n221_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n258_), .B1(new_n264_), .B2(new_n251_), .ZN(new_n265_));
  AOI211_X1 g064(.A(KEYINPUT70), .B(KEYINPUT12), .C1(new_n262_), .C2(new_n263_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n253_), .B(new_n257_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT68), .B1(new_n262_), .B2(new_n263_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n238_), .A2(new_n240_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(new_n222_), .A4(new_n259_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n222_), .B1(new_n269_), .B2(new_n259_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n256_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G120gat), .B(G148gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G176gat), .B(G204gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n267_), .A2(new_n274_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n280_), .B1(new_n267_), .B2(new_n274_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n284_), .B1(new_n287_), .B2(new_n285_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G29gat), .B(G36gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT73), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G43gat), .B(G50gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n291_), .B(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n250_), .A2(new_n294_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G232gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT34), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT35), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n294_), .A2(new_n298_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT15), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n299_), .B(new_n304_), .C1(new_n306_), .C2(new_n250_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT15), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n305_), .B(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n308_), .B1(new_n310_), .B2(new_n262_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n302_), .A2(new_n303_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n307_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n262_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n315_), .A2(new_n308_), .A3(new_n312_), .A4(new_n299_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G190gat), .B(G218gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G134gat), .B(G162gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n319_), .B(KEYINPUT36), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT75), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n314_), .A2(new_n316_), .A3(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n319_), .A2(KEYINPUT36), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT37), .B1(new_n322_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n314_), .A2(new_n316_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n323_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT37), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n314_), .A2(new_n316_), .A3(new_n320_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n326_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n332_), .B1(new_n326_), .B2(new_n331_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G15gat), .B(G22gat), .ZN(new_n336_));
  INV_X1    g135(.A(G1gat), .ZN(new_n337_));
  INV_X1    g136(.A(G8gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT14), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n336_), .B1(new_n339_), .B2(KEYINPUT77), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n339_), .A2(KEYINPUT77), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G1gat), .B(G8gat), .ZN(new_n342_));
  OR3_X1    g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n342_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT78), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G231gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n348_), .A2(new_n222_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n222_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G127gat), .B(G155gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT16), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G183gat), .B(G211gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT17), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n349_), .A2(new_n350_), .A3(new_n355_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n356_), .A2(KEYINPUT80), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(KEYINPUT80), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n359_));
  AOI211_X1 g158(.A(new_n354_), .B(new_n359_), .C1(new_n348_), .C2(new_n223_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(new_n223_), .B2(new_n348_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n357_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n335_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT81), .ZN(new_n365_));
  NAND2_X1  g164(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(G169gat), .ZN(new_n367_));
  INV_X1    g166(.A(G169gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n369_));
  INV_X1    g168(.A(G176gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n367_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT85), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n367_), .A2(new_n369_), .A3(KEYINPUT85), .A4(new_n370_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT23), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(G183gat), .A3(G190gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT86), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT23), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n382_), .A2(new_n377_), .A3(G183gat), .A4(G190gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n379_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT82), .B(G183gat), .ZN(new_n385_));
  INV_X1    g184(.A(G190gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n387_), .ZN(new_n388_));
  OR3_X1    g187(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n374_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n389_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n393_));
  INV_X1    g192(.A(G183gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n385_), .B2(new_n393_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT26), .B(G190gat), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n392_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n381_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n380_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n378_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n376_), .A2(new_n388_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G227gat), .A2(G233gat), .ZN(new_n404_));
  INV_X1    g203(.A(G71gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(G99gat), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n403_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n403_), .A2(new_n407_), .ZN(new_n409_));
  INV_X1    g208(.A(G134gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(G127gat), .ZN(new_n411_));
  INV_X1    g210(.A(G127gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(G134gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(G120gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G113gat), .ZN(new_n416_));
  INV_X1    g215(.A(G113gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(G120gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n414_), .A2(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n411_), .A2(new_n413_), .A3(new_n416_), .A4(new_n418_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OR3_X1    g222(.A1(new_n408_), .A2(new_n409_), .A3(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n423_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G15gat), .B(G43gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT87), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT30), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT31), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n426_), .B(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G228gat), .A2(G233gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(G78gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(G106gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G22gat), .B(G50gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(G141gat), .A2(G148gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT3), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT2), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n440_), .A2(new_n443_), .A3(new_n444_), .A4(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(G155gat), .A2(G162gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G155gat), .A2(G162gat), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(KEYINPUT1), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT1), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(G155gat), .A3(G162gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n452_), .A3(new_n447_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G141gat), .B(G148gat), .Z(new_n454_));
  AOI22_X1  g253(.A1(new_n446_), .A2(new_n449_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT29), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n457_), .B(KEYINPUT28), .Z(new_n458_));
  OR2_X1    g257(.A1(G197gat), .A2(G204gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G197gat), .A2(G204gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(KEYINPUT21), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT21), .ZN(new_n462_));
  AND2_X1   g261(.A1(G197gat), .A2(G204gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(G197gat), .A2(G204gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n462_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G211gat), .B(G218gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n463_), .A2(new_n464_), .A3(new_n462_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G211gat), .B(G218gat), .Z(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n458_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n458_), .A2(new_n473_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n437_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n476_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n474_), .A3(new_n436_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G29gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(G85gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT0), .B(G57gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT91), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n485_), .B1(new_n455_), .B2(new_n422_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n446_), .A2(new_n449_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n453_), .A2(new_n454_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n423_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n486_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n423_), .A3(new_n485_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G225gat), .A2(G233gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT92), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT92), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n497_), .A3(new_n494_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n490_), .A2(KEYINPUT4), .ZN(new_n500_));
  AOI211_X1 g299(.A(new_n494_), .B(new_n500_), .C1(new_n493_), .C2(KEYINPUT4), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n484_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n493_), .A2(KEYINPUT4), .ZN(new_n503_));
  INV_X1    g302(.A(new_n494_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n500_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n484_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n506_), .A2(new_n496_), .A3(new_n507_), .A4(new_n498_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n502_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n384_), .A2(new_n389_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n378_), .A2(KEYINPUT86), .B1(KEYINPUT23), .B2(new_n380_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n513_), .B1(new_n514_), .B2(new_n383_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT89), .ZN(new_n516_));
  NAND2_X1  g315(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT88), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT88), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n395_), .A2(new_n521_), .A3(new_n517_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n391_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n523_), .A2(new_n397_), .B1(new_n374_), .B2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n512_), .A2(new_n516_), .A3(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n402_), .B1(G183gat), .B2(G190gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT22), .B(G169gat), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n390_), .B1(new_n528_), .B2(new_n370_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n471_), .B1(new_n526_), .B2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n390_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n388_), .A2(new_n375_), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n513_), .B1(new_n524_), .B2(new_n374_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n394_), .A2(KEYINPUT82), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT82), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(G183gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n519_), .B1(new_n538_), .B2(KEYINPUT25), .ZN(new_n539_));
  INV_X1    g338(.A(new_n397_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n402_), .B(new_n534_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n533_), .A2(new_n471_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT20), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G226gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT19), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n531_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT90), .B1(new_n403_), .B2(new_n471_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT20), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n471_), .B1(new_n533_), .B2(new_n541_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT94), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n524_), .A2(new_n374_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n518_), .A2(new_n519_), .A3(KEYINPUT88), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n521_), .B1(new_n395_), .B2(new_n517_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n397_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n553_), .B(new_n556_), .C1(new_n515_), .C2(KEYINPUT89), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n510_), .A2(new_n511_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n552_), .B(new_n530_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n471_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n552_), .B1(new_n526_), .B2(new_n530_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n547_), .B(new_n551_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n546_), .B1(new_n562_), .B2(new_n545_), .ZN(new_n563_));
  XOR2_X1   g362(.A(G8gat), .B(G36gat), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT18), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G64gat), .B(G92gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT32), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT95), .B1(new_n563_), .B2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n545_), .B1(new_n531_), .B2(new_n543_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n551_), .A2(new_n547_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n526_), .A2(new_n471_), .A3(new_n530_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n545_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n568_), .B(new_n570_), .C1(new_n571_), .C2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT93), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n551_), .A2(new_n547_), .A3(new_n573_), .A4(new_n572_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n578_), .A2(KEYINPUT93), .A3(new_n568_), .A4(new_n570_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT95), .ZN(new_n581_));
  INV_X1    g380(.A(new_n568_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n384_), .A2(new_n387_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n541_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n550_), .A3(new_n472_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT20), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n549_), .A2(new_n550_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n530_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT94), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n471_), .A3(new_n559_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n573_), .B1(new_n589_), .B2(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n581_), .B(new_n582_), .C1(new_n593_), .C2(new_n546_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n509_), .A2(new_n569_), .A3(new_n580_), .A4(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT33), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n503_), .A2(new_n494_), .A3(new_n505_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n507_), .B1(new_n493_), .B2(new_n504_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n508_), .A2(new_n596_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n499_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n600_), .A2(KEYINPUT33), .A3(new_n507_), .A4(new_n506_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n578_), .A2(new_n567_), .A3(new_n570_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n567_), .B1(new_n578_), .B2(new_n570_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n599_), .A2(new_n601_), .A3(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n480_), .B1(new_n595_), .B2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n578_), .A2(new_n567_), .A3(new_n570_), .ZN(new_n607_));
  OAI211_X1 g406(.A(KEYINPUT27), .B(new_n607_), .C1(new_n563_), .C2(new_n567_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT27), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n609_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n480_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n509_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n431_), .B1(new_n606_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT96), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT96), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n616_), .B(new_n431_), .C1(new_n606_), .C2(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n431_), .A2(new_n509_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n611_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n619_), .A2(new_n620_), .A3(KEYINPUT97), .A4(new_n612_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n622_));
  INV_X1    g421(.A(new_n509_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n430_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n426_), .B(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n612_), .A2(new_n608_), .A3(new_n610_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n622_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n621_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n618_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n310_), .A2(new_n345_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n345_), .A2(new_n305_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G229gat), .A2(G233gat), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n345_), .B(new_n305_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n634_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n632_), .A2(new_n635_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(G113gat), .B(G141gat), .Z(new_n639_));
  XNOR2_X1  g438(.A(G169gat), .B(G197gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n638_), .B(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n630_), .A2(new_n631_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n629_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n642_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT98), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n290_), .B(new_n365_), .C1(new_n643_), .C2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n337_), .A3(new_n509_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n650_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n328_), .A2(new_n330_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n645_), .A2(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n290_), .A2(new_n646_), .A3(new_n362_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT100), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n658_), .A2(new_n509_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n651_), .B(new_n652_), .C1(new_n337_), .C2(new_n659_), .ZN(G1324gat));
  NAND2_X1  g459(.A1(new_n657_), .A2(new_n611_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G8gat), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT39), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n648_), .A2(new_n338_), .A3(new_n611_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n665_), .B(new_n667_), .ZN(G1325gat));
  INV_X1    g467(.A(G15gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n648_), .A2(new_n669_), .A3(new_n625_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n658_), .A2(new_n625_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n671_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT41), .B1(new_n671_), .B2(G15gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n672_), .B2(new_n673_), .ZN(G1326gat));
  INV_X1    g473(.A(G22gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n648_), .A2(new_n675_), .A3(new_n480_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n658_), .A2(new_n480_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G22gat), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n678_), .A2(KEYINPUT42), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(KEYINPUT42), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(G1327gat));
  NOR2_X1   g480(.A1(new_n363_), .A2(new_n653_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n289_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n643_), .B2(new_n647_), .ZN(new_n684_));
  INV_X1    g483(.A(G29gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n509_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n362_), .A2(new_n289_), .A3(new_n642_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n333_), .A2(new_n334_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n630_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT43), .B1(new_n645_), .B2(new_n335_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n687_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT102), .B(new_n688_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT103), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n688_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n689_), .B1(new_n630_), .B2(new_n690_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n645_), .A2(KEYINPUT43), .A3(new_n335_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT102), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n691_), .A2(new_n692_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(new_n694_), .A3(new_n698_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n702_), .A2(new_n703_), .A3(new_n687_), .A4(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n697_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n693_), .A2(KEYINPUT44), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n709_), .A2(new_n623_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n707_), .A2(KEYINPUT104), .A3(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G29gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT104), .B1(new_n707_), .B2(new_n710_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n686_), .B1(new_n712_), .B2(new_n713_), .ZN(G1328gat));
  INV_X1    g513(.A(G36gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n684_), .A2(new_n715_), .A3(new_n611_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT45), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n708_), .A2(new_n611_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n697_), .B2(new_n706_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n717_), .B(KEYINPUT46), .C1(new_n719_), .C2(new_n715_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n717_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n718_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT44), .B1(new_n701_), .B2(KEYINPUT102), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n703_), .B1(new_n723_), .B2(new_n705_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n695_), .A2(KEYINPUT103), .A3(new_n696_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n722_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n721_), .B1(new_n726_), .B2(G36gat), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n720_), .B1(new_n727_), .B2(new_n728_), .ZN(G1329gat));
  NAND2_X1  g528(.A1(new_n625_), .A2(G43gat), .ZN(new_n730_));
  AOI211_X1 g529(.A(new_n709_), .B(new_n730_), .C1(new_n697_), .C2(new_n706_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G43gat), .B1(new_n684_), .B2(new_n625_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT106), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT47), .B1(new_n731_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n707_), .A2(new_n708_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n736_), .B(new_n733_), .C1(new_n737_), .C2(new_n730_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n735_), .A2(new_n738_), .ZN(G1330gat));
  AOI21_X1  g538(.A(G50gat), .B1(new_n684_), .B2(new_n480_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n737_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n480_), .A2(G50gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(new_n741_), .B2(new_n742_), .ZN(G1331gat));
  NOR4_X1   g542(.A1(new_n365_), .A2(new_n645_), .A3(new_n642_), .A4(new_n289_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(new_n211_), .A3(new_n509_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n655_), .A2(new_n646_), .A3(new_n290_), .A4(new_n363_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G57gat), .B1(new_n746_), .B2(new_n623_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT107), .Z(G1332gat));
  OAI21_X1  g548(.A(G64gat), .B1(new_n746_), .B2(new_n620_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT48), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n744_), .A2(new_n209_), .A3(new_n611_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1333gat));
  OAI21_X1  g552(.A(G71gat), .B1(new_n746_), .B2(new_n431_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT49), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n744_), .A2(new_n405_), .A3(new_n625_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1334gat));
  OAI21_X1  g556(.A(G78gat), .B1(new_n746_), .B2(new_n612_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT50), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n612_), .A2(G78gat), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT108), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n744_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n762_), .ZN(G1335gat));
  NAND4_X1  g562(.A1(new_n630_), .A2(new_n646_), .A3(new_n290_), .A4(new_n682_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT109), .Z(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(new_n232_), .A3(new_n509_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n363_), .A2(new_n642_), .A3(new_n289_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n699_), .A2(new_n700_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n704_), .A2(KEYINPUT110), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n773_), .A2(new_n509_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n766_), .B1(new_n774_), .B2(new_n232_), .ZN(G1336gat));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n611_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n620_), .A2(G92gat), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n776_), .A2(G92gat), .B1(new_n765_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n778_), .B(new_n779_), .ZN(G1337gat));
  NAND2_X1  g579(.A1(new_n773_), .A2(new_n625_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(G99gat), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n244_), .A2(new_n245_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n431_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT112), .B1(new_n765_), .B2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n782_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1338gat));
  NAND2_X1  g588(.A1(new_n767_), .A2(new_n480_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G106gat), .B1(new_n769_), .B2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT52), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n765_), .A2(new_n480_), .A3(new_n241_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g594(.A1(new_n289_), .A2(new_n646_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n364_), .A2(KEYINPUT54), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n690_), .A2(new_n362_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n796_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n797_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n642_), .A2(new_n281_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n268_), .A2(new_n271_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n805_), .B(new_n253_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n256_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n267_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT70), .B1(new_n273_), .B2(KEYINPUT12), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n264_), .A2(new_n258_), .A3(new_n251_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n814_), .A2(KEYINPUT55), .A3(new_n253_), .A4(new_n257_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n811_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n807_), .B1(new_n806_), .B2(new_n256_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n809_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n804_), .B1(new_n818_), .B2(new_n280_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n253_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n256_), .B1(new_n820_), .B2(new_n272_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT114), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n822_), .A2(new_n808_), .A3(new_n811_), .A4(new_n815_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(KEYINPUT56), .A3(new_n279_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n803_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n632_), .A2(new_n633_), .A3(new_n637_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n641_), .B1(new_n636_), .B2(new_n634_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n638_), .A2(new_n641_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n653_), .B1(new_n825_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT57), .B(new_n653_), .C1(new_n825_), .C2(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n828_), .A2(new_n281_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT116), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n828_), .A2(new_n838_), .A3(new_n281_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n823_), .A2(KEYINPUT56), .A3(new_n279_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT56), .B1(new_n823_), .B2(new_n279_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n840_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT58), .B(new_n840_), .C1(new_n841_), .C2(new_n842_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n690_), .A3(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n834_), .A2(new_n835_), .A3(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n363_), .B1(new_n848_), .B2(KEYINPUT117), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n834_), .A2(new_n847_), .A3(new_n850_), .A4(new_n835_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n802_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n627_), .A2(new_n623_), .A3(new_n431_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n417_), .A3(new_n642_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT59), .B1(new_n852_), .B2(new_n854_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n854_), .A2(KEYINPUT59), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT118), .B1(new_n834_), .B2(new_n847_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n835_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n834_), .A2(KEYINPUT118), .A3(new_n847_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n363_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n858_), .B1(new_n863_), .B2(new_n802_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n857_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n857_), .B2(new_n864_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n646_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n856_), .B1(new_n868_), .B2(new_n417_), .ZN(G1340gat));
  OAI21_X1  g668(.A(new_n415_), .B1(new_n289_), .B2(KEYINPUT60), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n855_), .B(new_n870_), .C1(KEYINPUT60), .C2(new_n415_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n857_), .A2(new_n864_), .A3(new_n290_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n415_), .ZN(G1341gat));
  NAND3_X1  g672(.A1(new_n855_), .A2(new_n412_), .A3(new_n363_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n866_), .A2(new_n867_), .A3(new_n362_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n412_), .ZN(G1342gat));
  NAND3_X1  g675(.A1(new_n855_), .A2(new_n410_), .A3(new_n654_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n866_), .A2(new_n867_), .A3(new_n335_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n410_), .ZN(G1343gat));
  NAND2_X1  g678(.A1(new_n848_), .A2(KEYINPUT117), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(new_n362_), .A3(new_n851_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n802_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884_));
  NOR4_X1   g683(.A1(new_n611_), .A2(new_n623_), .A3(new_n625_), .A4(new_n612_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n885_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT120), .B1(new_n852_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n642_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT121), .B(G141gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1344gat));
  NAND2_X1  g691(.A1(new_n889_), .A2(new_n290_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n889_), .B2(new_n363_), .ZN(new_n898_));
  AOI211_X1 g697(.A(KEYINPUT122), .B(new_n362_), .C1(new_n886_), .C2(new_n888_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n896_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n884_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n852_), .A2(KEYINPUT120), .A3(new_n887_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n363_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT122), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n889_), .A2(new_n897_), .A3(new_n363_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n904_), .A2(new_n905_), .A3(new_n895_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n900_), .A2(new_n906_), .ZN(G1346gat));
  INV_X1    g706(.A(new_n889_), .ZN(new_n908_));
  OR3_X1    g707(.A1(new_n908_), .A2(G162gat), .A3(new_n653_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G162gat), .B1(new_n908_), .B2(new_n335_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1347gat));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n863_), .A2(new_n802_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n620_), .A2(new_n626_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n480_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n913_), .A2(new_n528_), .A3(new_n642_), .A4(new_n916_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n642_), .B(new_n916_), .C1(new_n863_), .C2(new_n802_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n918_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(KEYINPUT62), .B1(new_n918_), .B2(G169gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n912_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n921_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n923_), .A2(KEYINPUT123), .A3(new_n917_), .A4(new_n919_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1348gat));
  NOR2_X1   g724(.A1(new_n852_), .A2(new_n480_), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n926_), .A2(G176gat), .A3(new_n290_), .A4(new_n914_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n863_), .A2(new_n802_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n916_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n928_), .A2(new_n289_), .A3(new_n929_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n927_), .B1(new_n930_), .B2(G176gat), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(KEYINPUT124), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933_));
  OAI211_X1 g732(.A(new_n933_), .B(new_n927_), .C1(new_n930_), .C2(G176gat), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n934_), .ZN(G1349gat));
  NAND3_X1  g734(.A1(new_n926_), .A2(new_n363_), .A3(new_n914_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(KEYINPUT125), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n928_), .A2(new_n929_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n362_), .A2(new_n523_), .ZN(new_n939_));
  AOI22_X1  g738(.A1(new_n937_), .A2(new_n385_), .B1(new_n938_), .B2(new_n939_), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n938_), .A2(new_n397_), .A3(new_n654_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n928_), .A2(new_n335_), .A3(new_n929_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n386_), .B2(new_n942_), .ZN(G1351gat));
  NOR3_X1   g742(.A1(new_n625_), .A2(new_n612_), .A3(new_n509_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(KEYINPUT126), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n944_), .A2(KEYINPUT126), .ZN(new_n946_));
  NOR4_X1   g745(.A1(new_n852_), .A2(new_n620_), .A3(new_n945_), .A4(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n642_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n290_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g750(.A1(new_n947_), .A2(new_n363_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  AND2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n952_), .A2(new_n953_), .A3(new_n954_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n955_), .B1(new_n952_), .B2(new_n953_), .ZN(G1354gat));
  NAND2_X1  g755(.A1(new_n947_), .A2(new_n654_), .ZN(new_n957_));
  XOR2_X1   g756(.A(KEYINPUT127), .B(G218gat), .Z(new_n958_));
  NOR2_X1   g757(.A1(new_n335_), .A2(new_n958_), .ZN(new_n959_));
  AOI22_X1  g758(.A1(new_n957_), .A2(new_n958_), .B1(new_n947_), .B2(new_n959_), .ZN(G1355gat));
endmodule


