//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_;
  INV_X1    g000(.A(KEYINPUT107), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n203_), .B(KEYINPUT101), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT4), .ZN(new_n206_));
  INV_X1    g005(.A(G120gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G113gat), .ZN(new_n208_));
  INV_X1    g007(.A(G113gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G120gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G127gat), .B(G134gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(G127gat), .A2(G134gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G127gat), .A2(G134gat), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n214_), .A2(new_n208_), .A3(new_n210_), .A4(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G141gat), .A2(G148gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n221_), .B1(new_n222_), .B2(KEYINPUT87), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT87), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n224_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(KEYINPUT87), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n223_), .A2(new_n225_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(G141gat), .A2(G148gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(KEYINPUT3), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n220_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n218_), .A2(new_n232_), .A3(new_n219_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n233_), .A2(new_n229_), .A3(new_n221_), .A4(new_n234_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n231_), .A2(KEYINPUT88), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT88), .B1(new_n231_), .B2(new_n235_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n217_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n217_), .A2(KEYINPUT100), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT100), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n213_), .A2(new_n240_), .A3(new_n216_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n239_), .A2(new_n231_), .A3(new_n235_), .A4(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n206_), .B1(new_n238_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n231_), .A2(new_n235_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT88), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n231_), .A2(KEYINPUT88), .A3(new_n235_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT4), .B1(new_n248_), .B2(new_n217_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n205_), .B1(new_n243_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT102), .ZN(new_n251_));
  INV_X1    g050(.A(new_n242_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n252_), .B1(new_n248_), .B2(new_n217_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(new_n203_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT102), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n255_), .B(new_n205_), .C1(new_n243_), .C2(new_n249_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n251_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G1gat), .B(G29gat), .ZN(new_n258_));
  INV_X1    g057(.A(G85gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G57gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(new_n261_), .Z(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n262_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n251_), .A2(new_n254_), .A3(new_n256_), .A4(new_n264_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT95), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT89), .B(G204gat), .ZN(new_n268_));
  INV_X1    g067(.A(G197gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT91), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G204gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT89), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT89), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(G204gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT91), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(G197gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n269_), .A2(G204gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n270_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G211gat), .B(G218gat), .Z(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(KEYINPUT21), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT21), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n270_), .A2(new_n277_), .A3(new_n283_), .A4(new_n278_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT92), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT90), .B1(new_n275_), .B2(G197gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n271_), .A2(G197gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT90), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n268_), .A2(new_n289_), .A3(new_n269_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n280_), .B1(new_n291_), .B2(KEYINPUT21), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n282_), .B1(new_n286_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT29), .B1(new_n236_), .B2(new_n237_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G228gat), .A2(G233gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n276_), .B1(new_n275_), .B2(G197gat), .ZN(new_n298_));
  AOI211_X1 g097(.A(KEYINPUT91), .B(new_n269_), .C1(new_n272_), .C2(new_n274_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n300_), .A2(new_n285_), .A3(new_n283_), .A4(new_n278_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n284_), .A2(KEYINPUT92), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n292_), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n281_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n244_), .A2(KEYINPUT29), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n295_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n267_), .B1(new_n297_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G78gat), .B(G106gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT93), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n304_), .A2(new_n295_), .A3(new_n294_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n303_), .A2(new_n281_), .B1(KEYINPUT29), .B2(new_n244_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n310_), .B(KEYINPUT95), .C1(new_n295_), .C2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n307_), .A2(new_n309_), .A3(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n297_), .A2(new_n306_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n309_), .B(KEYINPUT94), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  OR3_X1    g115(.A1(new_n248_), .A2(KEYINPUT29), .A3(G50gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT28), .B(G22gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(G50gat), .B1(new_n248_), .B2(KEYINPUT29), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n318_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n313_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT96), .ZN(new_n324_));
  INV_X1    g123(.A(new_n316_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n314_), .A2(new_n315_), .ZN(new_n326_));
  OAI22_X1  g125(.A1(new_n325_), .A2(new_n326_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT96), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n313_), .A2(new_n328_), .A3(new_n322_), .A4(new_n316_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n324_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT20), .ZN(new_n331_));
  INV_X1    g130(.A(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT26), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT26), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(G190gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT97), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n341_));
  INV_X1    g140(.A(G183gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT97), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(new_n337_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n336_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT98), .ZN(new_n348_));
  INV_X1    g147(.A(G169gat), .ZN(new_n349_));
  INV_X1    g148(.A(G176gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT24), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(G169gat), .B2(G176gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n347_), .A2(new_n348_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT98), .B1(new_n346_), .B2(new_n353_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT23), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n351_), .A2(KEYINPUT24), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n355_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n358_), .B1(G183gat), .B2(G190gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT83), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT22), .B(G169gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n363_), .B(new_n365_), .C1(G176gat), .C2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n362_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n331_), .B1(new_n304_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n352_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n365_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT84), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT81), .B(G183gat), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n339_), .B1(new_n374_), .B2(KEYINPUT25), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(KEYINPUT26), .B2(new_n332_), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n335_), .B(KEYINPUT82), .Z(new_n377_));
  AOI21_X1  g176(.A(new_n360_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(G176gat), .B1(new_n367_), .B2(KEYINPUT85), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT85), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n380_), .B1(new_n349_), .B2(KEYINPUT22), .ZN(new_n381_));
  INV_X1    g180(.A(new_n374_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n332_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n379_), .A2(new_n381_), .B1(new_n383_), .B2(new_n358_), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n373_), .A2(new_n378_), .B1(new_n365_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n293_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n370_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT19), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394_));
  XOR2_X1   g193(.A(new_n393_), .B(new_n394_), .Z(new_n395_));
  NAND4_X1  g194(.A1(new_n303_), .A2(new_n281_), .A3(new_n368_), .A4(new_n362_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT20), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n293_), .A2(new_n385_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n389_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n390_), .B(new_n395_), .C1(new_n397_), .C2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT27), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n396_), .A2(KEYINPUT104), .A3(KEYINPUT20), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT104), .B1(new_n396_), .B2(KEYINPUT20), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n293_), .A2(new_n385_), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT105), .B1(new_n406_), .B2(new_n399_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n387_), .A2(new_n389_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT104), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n397_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n396_), .A2(KEYINPUT104), .A3(KEYINPUT20), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n398_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT105), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(new_n389_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n407_), .A2(new_n409_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n395_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n402_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT106), .B(KEYINPUT27), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n405_), .A2(new_n397_), .A3(new_n389_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n399_), .B1(new_n370_), .B2(new_n386_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n417_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n420_), .B1(new_n401_), .B2(new_n423_), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n330_), .A2(new_n418_), .A3(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n421_), .A2(new_n422_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n395_), .A2(KEYINPUT32), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n263_), .A2(new_n265_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n413_), .A2(new_n414_), .A3(new_n389_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n414_), .B1(new_n413_), .B2(new_n389_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n408_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n428_), .B1(new_n431_), .B2(new_n427_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT103), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n238_), .A2(new_n206_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(new_n253_), .B2(new_n206_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n255_), .B1(new_n435_), .B2(new_n205_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n256_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n438_), .A2(KEYINPUT33), .A3(new_n254_), .A4(new_n264_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n265_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n435_), .A2(new_n203_), .B1(new_n253_), .B2(new_n205_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n262_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n401_), .A2(new_n423_), .A3(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n433_), .B1(new_n442_), .B2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n401_), .A2(new_n423_), .A3(new_n444_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n447_), .A2(KEYINPUT103), .A3(new_n441_), .A4(new_n439_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n432_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n266_), .A2(new_n425_), .B1(new_n449_), .B2(new_n330_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n385_), .B(KEYINPUT30), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G43gat), .ZN(new_n452_));
  XOR2_X1   g251(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n454_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G227gat), .A2(G233gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(G15gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G71gat), .B(G99gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(new_n217_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n455_), .A2(new_n456_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n461_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n202_), .B1(new_n450_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n330_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n418_), .A2(new_n424_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n266_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n449_), .A2(new_n330_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n468_), .A3(new_n266_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(KEYINPUT107), .A3(new_n467_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n466_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G29gat), .B(G36gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G50gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(KEYINPUT73), .B(G43gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT15), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT68), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT65), .B1(KEYINPUT66), .B2(KEYINPUT7), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G99gat), .A2(G106gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n488_), .B(new_n489_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G85gat), .B(G92gat), .Z(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n482_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  OAI211_X1 g293(.A(KEYINPUT68), .B(new_n492_), .C1(new_n485_), .C2(new_n490_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(KEYINPUT8), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT67), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT8), .B1(new_n491_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT67), .B1(new_n485_), .B2(new_n490_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n492_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT9), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n503_), .B1(new_n492_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT64), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n488_), .A2(new_n489_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT10), .B(G99gat), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n509_), .A2(G106gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n506_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n507_), .A2(new_n508_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n501_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n481_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n501_), .A2(new_n512_), .A3(new_n480_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G232gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT34), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n514_), .B(new_n515_), .C1(KEYINPUT35), .C2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(KEYINPUT35), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT72), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n518_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G190gat), .B(G218gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G134gat), .B(G162gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OR3_X1    g324(.A1(new_n521_), .A2(KEYINPUT36), .A3(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n524_), .B(KEYINPUT36), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n521_), .A2(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT37), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n528_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT37), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G57gat), .B(G64gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT69), .B(G71gat), .ZN(new_n536_));
  INV_X1    g335(.A(G78gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT11), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n536_), .A2(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n537_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(KEYINPUT11), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n535_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n543_), .A2(new_n535_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(G1gat), .ZN(new_n549_));
  INV_X1    g348(.A(G8gat), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT14), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n551_), .A2(KEYINPUT74), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G15gat), .B(G22gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(KEYINPUT74), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT75), .ZN(new_n556_));
  XOR2_X1   g355(.A(G1gat), .B(G8gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n548_), .B(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT77), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G183gat), .B(G211gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(G127gat), .B(G155gat), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT17), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n560_), .B(new_n566_), .ZN(new_n567_));
  OR3_X1    g366(.A1(new_n559_), .A2(KEYINPUT17), .A3(new_n565_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n530_), .A2(new_n533_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n501_), .A2(new_n512_), .A3(new_n546_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n546_), .B1(new_n501_), .B2(new_n512_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n574_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(G230gat), .ZN(new_n578_));
  INV_X1    g377(.A(G233gat), .ZN(new_n579_));
  OAI22_X1  g378(.A1(new_n575_), .A2(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n578_), .A2(new_n579_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G120gat), .B(G148gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT71), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G176gat), .B(G204gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n587_), .B(new_n588_), .Z(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n589_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n580_), .A2(new_n582_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT13), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n590_), .A2(KEYINPUT13), .A3(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n558_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n481_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n480_), .B(KEYINPUT78), .Z(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n558_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n600_), .B(new_n558_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n603_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G113gat), .B(G141gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G169gat), .B(G197gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(KEYINPUT79), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT80), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n608_), .B(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n597_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n476_), .A2(new_n571_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT108), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n266_), .B(KEYINPUT109), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n549_), .A3(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(KEYINPUT110), .B(KEYINPUT38), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n616_), .B(KEYINPUT111), .Z(new_n625_));
  NAND4_X1  g424(.A1(new_n476_), .A2(new_n531_), .A3(new_n569_), .A4(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n266_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT112), .Z(new_n628_));
  NAND2_X1  g427(.A1(new_n624_), .A2(new_n628_), .ZN(G1324gat));
  INV_X1    g428(.A(new_n470_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n619_), .A2(new_n550_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  INV_X1    g431(.A(new_n626_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n630_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n632_), .B1(new_n634_), .B2(G8gat), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n632_), .B(G8gat), .C1(new_n626_), .C2(new_n470_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n631_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n631_), .B(KEYINPUT40), .C1(new_n635_), .C2(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1325gat));
  NAND2_X1  g441(.A1(new_n633_), .A2(new_n465_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT41), .B1(new_n643_), .B2(G15gat), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n467_), .A2(G15gat), .ZN(new_n647_));
  OAI22_X1  g446(.A1(new_n645_), .A2(new_n646_), .B1(new_n617_), .B2(new_n647_), .ZN(G1326gat));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n633_), .A2(new_n468_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(G22gat), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n649_), .B(G22gat), .C1(new_n626_), .C2(new_n330_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n330_), .A2(G22gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT113), .ZN(new_n655_));
  OAI22_X1  g454(.A1(new_n651_), .A2(new_n653_), .B1(new_n617_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT114), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(G1327gat));
  INV_X1    g457(.A(new_n569_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n529_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT115), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n476_), .A2(new_n616_), .A3(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n266_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(G29gat), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n625_), .A2(new_n659_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n530_), .A2(new_n533_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n476_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n667_), .B1(new_n476_), .B2(new_n668_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n673_), .A2(G29gat), .A3(new_n621_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n666_), .B(KEYINPUT44), .C1(new_n669_), .C2(new_n670_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n664_), .B1(new_n674_), .B2(new_n675_), .ZN(G1328gat));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  INV_X1    g476(.A(G36gat), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n476_), .A2(new_n668_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT43), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n476_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n665_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n470_), .B1(new_n682_), .B2(KEYINPUT44), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n678_), .B1(new_n683_), .B2(new_n673_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n662_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n678_), .A3(new_n630_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT45), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n687_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n677_), .B1(new_n684_), .B2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n682_), .A2(KEYINPUT44), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n675_), .A2(new_n630_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G36gat), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n694_), .A2(KEYINPUT46), .A3(new_n689_), .A4(new_n688_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n691_), .A2(new_n695_), .ZN(G1329gat));
  NAND4_X1  g495(.A1(new_n673_), .A2(G43gat), .A3(new_n465_), .A4(new_n675_), .ZN(new_n697_));
  INV_X1    g496(.A(G43gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n698_), .B1(new_n662_), .B2(new_n467_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT47), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n697_), .A2(new_n702_), .A3(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1330gat));
  AOI21_X1  g503(.A(G50gat), .B1(new_n685_), .B2(new_n468_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n675_), .A2(G50gat), .A3(new_n468_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(new_n673_), .ZN(G1331gat));
  AND3_X1   g506(.A1(new_n476_), .A2(new_n531_), .A3(new_n569_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n597_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n615_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n708_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(G57gat), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n712_), .A2(new_n713_), .A3(new_n266_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n476_), .A2(new_n615_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT116), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n717_), .A2(new_n597_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n621_), .A3(new_n571_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n714_), .B1(new_n719_), .B2(new_n713_), .ZN(G1332gat));
  INV_X1    g519(.A(new_n712_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n630_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n723_), .A3(G64gat), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n723_), .B1(new_n722_), .B2(G64gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n718_), .A2(new_n571_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n470_), .A2(G64gat), .ZN(new_n728_));
  OAI22_X1  g527(.A1(new_n725_), .A2(new_n726_), .B1(new_n727_), .B2(new_n728_), .ZN(G1333gat));
  NAND2_X1  g528(.A1(new_n721_), .A2(new_n465_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT49), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(G71gat), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n730_), .B2(G71gat), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n467_), .A2(G71gat), .ZN(new_n735_));
  OAI22_X1  g534(.A1(new_n733_), .A2(new_n734_), .B1(new_n727_), .B2(new_n735_), .ZN(G1334gat));
  NAND2_X1  g535(.A1(new_n721_), .A2(new_n468_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n738_), .A3(G78gat), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n737_), .B2(G78gat), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n468_), .A2(new_n537_), .ZN(new_n742_));
  OAI22_X1  g541(.A1(new_n740_), .A2(new_n741_), .B1(new_n727_), .B2(new_n742_), .ZN(G1335gat));
  NAND3_X1  g542(.A1(new_n718_), .A2(new_n621_), .A3(new_n661_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n711_), .A2(new_n659_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n266_), .A2(new_n259_), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n744_), .A2(new_n259_), .B1(new_n746_), .B2(new_n747_), .ZN(G1336gat));
  NAND3_X1  g547(.A1(new_n718_), .A2(new_n630_), .A3(new_n661_), .ZN(new_n749_));
  INV_X1    g548(.A(G92gat), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n470_), .A2(new_n750_), .ZN(new_n751_));
  AOI22_X1  g550(.A1(new_n749_), .A2(new_n750_), .B1(new_n746_), .B2(new_n751_), .ZN(G1337gat));
  NAND2_X1  g551(.A1(new_n746_), .A2(new_n465_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G99gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n717_), .A2(new_n597_), .A3(new_n661_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n467_), .A2(new_n509_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n754_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT51), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n754_), .B(new_n760_), .C1(new_n755_), .C2(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1338gat));
  NOR2_X1   g561(.A1(new_n330_), .A2(G106gat), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n717_), .A2(new_n597_), .A3(new_n661_), .A4(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n745_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n468_), .B(new_n765_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G106gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n772_), .B(new_n764_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1339gat));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n570_), .A2(new_n597_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n615_), .ZN(new_n777_));
  NOR4_X1   g576(.A1(new_n570_), .A2(new_n597_), .A3(KEYINPUT54), .A4(new_n710_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n580_), .A2(KEYINPUT117), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n546_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n513_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n501_), .A2(new_n512_), .A3(new_n546_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(KEYINPUT12), .A3(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(KEYINPUT118), .A3(new_n576_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n783_), .A2(new_n581_), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n581_), .B1(new_n787_), .B2(new_n576_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT55), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n781_), .A2(new_n789_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n589_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n589_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(KEYINPUT119), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n793_), .A2(new_n799_), .A3(KEYINPUT56), .A4(new_n589_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n798_), .A2(new_n592_), .A3(new_n710_), .A4(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n602_), .A2(new_n603_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n605_), .A2(new_n606_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n611_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n604_), .A2(new_n607_), .A3(new_n612_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n593_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n806_), .B2(new_n593_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n801_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n531_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n796_), .A2(new_n797_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(new_n592_), .A3(new_n806_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT58), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(new_n817_), .A3(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n668_), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n811_), .A2(KEYINPUT57), .A3(new_n531_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n814_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n779_), .B1(new_n824_), .B2(new_n659_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n469_), .A2(new_n470_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n825_), .A2(new_n620_), .A3(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n710_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT122), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n825_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n827_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n826_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT57), .B1(new_n811_), .B2(new_n531_), .ZN(new_n834_));
  AOI211_X1 g633(.A(new_n813_), .B(new_n529_), .C1(new_n801_), .C2(new_n810_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n569_), .B1(new_n836_), .B2(new_n822_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n621_), .B(new_n833_), .C1(new_n837_), .C2(new_n779_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT122), .B1(new_n837_), .B2(new_n779_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n829_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n832_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n710_), .A2(G113gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT123), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n828_), .B1(new_n841_), .B2(new_n843_), .ZN(G1340gat));
  INV_X1    g643(.A(KEYINPUT60), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n709_), .B2(G120gat), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n827_), .B(new_n846_), .C1(new_n845_), .C2(G120gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n709_), .B1(new_n832_), .B2(new_n840_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(new_n207_), .ZN(G1341gat));
  AOI21_X1  g648(.A(G127gat), .B1(new_n827_), .B2(new_n569_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n659_), .B1(new_n832_), .B2(new_n840_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g651(.A(G134gat), .B1(new_n827_), .B2(new_n529_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n668_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n832_), .B2(new_n840_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n855_), .B2(G134gat), .ZN(G1343gat));
  INV_X1    g655(.A(new_n425_), .ZN(new_n857_));
  NOR4_X1   g656(.A1(new_n825_), .A2(new_n620_), .A3(new_n465_), .A4(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n710_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n597_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g661(.A1(new_n858_), .A2(new_n569_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1346gat));
  AOI21_X1  g664(.A(G162gat), .B1(new_n858_), .B2(new_n529_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n668_), .A2(G162gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n858_), .B2(new_n867_), .ZN(G1347gat));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n824_), .A2(new_n659_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n779_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n621_), .A2(new_n470_), .ZN(new_n873_));
  AND4_X1   g672(.A1(new_n710_), .A2(new_n872_), .A3(new_n469_), .A4(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n869_), .B1(new_n874_), .B2(new_n349_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n825_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n710_), .A3(new_n873_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n874_), .A2(new_n366_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n875_), .A2(new_n878_), .A3(new_n879_), .ZN(G1348gat));
  NAND3_X1  g679(.A1(new_n876_), .A2(new_n597_), .A3(new_n873_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G176gat), .ZN(G1349gat));
  NAND4_X1  g681(.A1(new_n872_), .A2(new_n569_), .A3(new_n469_), .A4(new_n873_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n340_), .A2(new_n345_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n382_), .B2(new_n883_), .ZN(G1350gat));
  NAND2_X1  g685(.A1(new_n876_), .A2(new_n873_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G190gat), .B1(new_n887_), .B2(new_n854_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n531_), .A2(new_n336_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n887_), .B2(new_n889_), .ZN(G1351gat));
  INV_X1    g689(.A(KEYINPUT125), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n467_), .A2(new_n266_), .A3(new_n468_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT124), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n872_), .A2(new_n710_), .A3(new_n630_), .A4(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n891_), .B1(new_n895_), .B2(new_n269_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n269_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n825_), .A2(new_n470_), .A3(new_n893_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n898_), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n710_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n896_), .A2(new_n897_), .A3(new_n899_), .ZN(G1352gat));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n597_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G204gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n268_), .B2(new_n901_), .ZN(G1353gat));
  XOR2_X1   g702(.A(KEYINPUT63), .B(G211gat), .Z(new_n904_));
  AND3_X1   g703(.A1(new_n898_), .A2(new_n569_), .A3(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n898_), .A2(new_n569_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(G1354gat));
  NAND2_X1  g707(.A1(new_n668_), .A2(G218gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(KEYINPUT126), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n872_), .A2(new_n630_), .A3(new_n894_), .A4(new_n910_), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n825_), .A2(new_n531_), .A3(new_n470_), .A4(new_n893_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(G218gat), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT127), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  OAI211_X1 g714(.A(KEYINPUT127), .B(new_n911_), .C1(new_n912_), .C2(G218gat), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1355gat));
endmodule


