//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_;
  XNOR2_X1  g000(.A(KEYINPUT80), .B(G8gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT81), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n207_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G29gat), .B(G36gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT85), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n214_), .A2(KEYINPUT84), .A3(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n215_), .B1(new_n214_), .B2(KEYINPUT84), .ZN(new_n217_));
  OAI22_X1  g016(.A1(new_n216_), .A2(new_n217_), .B1(new_n210_), .B2(new_n213_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(KEYINPUT84), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT85), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n210_), .A2(new_n213_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n214_), .A2(KEYINPUT84), .A3(new_n215_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n218_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n207_), .B(new_n208_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n213_), .B(KEYINPUT15), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n214_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n224_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n226_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G141gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G169gat), .B(G197gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n226_), .A2(new_n231_), .A3(new_n235_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT86), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G120gat), .B(G148gat), .Z(new_n242_));
  XNOR2_X1  g041(.A(G176gat), .B(G204gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n244_), .B(new_n245_), .Z(new_n246_));
  XOR2_X1   g045(.A(G85gat), .B(G92gat), .Z(new_n247_));
  NOR2_X1   g046(.A1(KEYINPUT9), .A2(G92gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n249_));
  OR3_X1    g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G99gat), .A2(G106gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT6), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n249_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT10), .B(G99gat), .Z(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT64), .B(G106gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n250_), .A2(new_n252_), .A3(new_n253_), .A4(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n257_), .A2(KEYINPUT68), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n259_));
  OR3_X1    g058(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n252_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT8), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G85gat), .B(G92gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n261_), .A2(new_n247_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n265_), .B1(new_n261_), .B2(new_n247_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT67), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n261_), .A2(new_n247_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n265_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n266_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n257_), .A2(KEYINPUT68), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n258_), .A2(new_n269_), .A3(new_n274_), .A4(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G57gat), .B(G64gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT11), .ZN(new_n278_));
  XOR2_X1   g077(.A(G71gat), .B(G78gat), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n277_), .A2(KEYINPUT11), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n278_), .A2(new_n279_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n276_), .A2(KEYINPUT12), .A3(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n267_), .A2(new_n268_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n257_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n284_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT12), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n284_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n286_), .A2(new_n292_), .A3(new_n257_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G230gat), .A2(G233gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(KEYINPUT69), .A3(new_n294_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n291_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n288_), .A2(new_n293_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(G230gat), .A3(G233gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n246_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n302_), .A3(new_n246_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n300_), .A2(KEYINPUT71), .A3(new_n302_), .A4(new_n246_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n303_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n308_), .A2(new_n312_), .ZN(new_n313_));
  AOI211_X1 g112(.A(new_n303_), .B(new_n310_), .C1(new_n306_), .C2(new_n307_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n308_), .A2(new_n312_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT73), .B1(new_n318_), .B2(new_n314_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n241_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n210_), .B(new_n292_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G231gat), .A2(G233gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n323_), .B(KEYINPUT82), .Z(new_n324_));
  XNOR2_X1  g123(.A(new_n322_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT83), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G127gat), .B(G155gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT16), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G183gat), .B(G211gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT17), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n327_), .B(new_n332_), .ZN(new_n333_));
  OR3_X1    g132(.A1(new_n325_), .A2(KEYINPUT17), .A3(new_n331_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G134gat), .B(G162gat), .Z(new_n337_));
  XNOR2_X1  g136(.A(G190gat), .B(G218gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT36), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n341_), .B(KEYINPUT77), .Z(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G232gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT35), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n346_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n349_), .A2(KEYINPUT76), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n345_), .A2(KEYINPUT35), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n286_), .A2(KEYINPUT75), .A3(new_n213_), .A4(new_n257_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n257_), .A2(new_n272_), .A3(new_n213_), .A4(new_n266_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n351_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n276_), .A2(new_n228_), .ZN(new_n357_));
  AOI211_X1 g156(.A(new_n348_), .B(new_n350_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(KEYINPUT76), .A4(new_n349_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n342_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT78), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n363_), .B(new_n342_), .C1(new_n358_), .C2(new_n360_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n350_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(new_n347_), .B2(new_n346_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n339_), .A2(new_n340_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n366_), .A2(new_n359_), .A3(new_n341_), .A4(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n362_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n368_), .A2(new_n361_), .ZN(new_n370_));
  XOR2_X1   g169(.A(KEYINPUT79), .B(KEYINPUT37), .Z(new_n371_));
  AOI22_X1  g170(.A1(new_n369_), .A2(KEYINPUT37), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n336_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G113gat), .B(G120gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G134gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(G127gat), .ZN(new_n377_));
  INV_X1    g176(.A(G127gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G134gat), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n377_), .A2(new_n379_), .A3(KEYINPUT90), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT90), .B1(new_n377_), .B2(new_n379_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n375_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n377_), .A2(new_n379_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT90), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n377_), .A2(new_n379_), .A3(KEYINPUT90), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n374_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT31), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT25), .B(G183gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT26), .B(G190gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G183gat), .A2(G190gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT23), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT23), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(G183gat), .A3(G190gat), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n391_), .A2(new_n392_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT24), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT87), .B1(G169gat), .B2(G176gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(KEYINPUT87), .A2(G169gat), .A3(G176gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n398_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT87), .ZN(new_n403_));
  INV_X1    g202(.A(G169gat), .ZN(new_n404_));
  INV_X1    g203(.A(G176gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(KEYINPUT24), .A3(new_n399_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G169gat), .A2(G176gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT88), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n397_), .B(new_n402_), .C1(new_n407_), .C2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n394_), .A2(new_n396_), .ZN(new_n411_));
  INV_X1    g210(.A(G183gat), .ZN(new_n412_));
  INV_X1    g211(.A(G190gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(KEYINPUT89), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n393_), .A2(new_n395_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(new_n414_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT88), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n408_), .B(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n404_), .A2(KEYINPUT22), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n404_), .A2(KEYINPUT22), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n405_), .A3(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n415_), .A2(new_n420_), .A3(new_n422_), .A4(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n410_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G71gat), .B(G99gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(G43gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n427_), .B(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G227gat), .A2(G233gat), .ZN(new_n431_));
  INV_X1    g230(.A(G15gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT30), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n430_), .B(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT91), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n390_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(new_n436_), .B2(new_n435_), .ZN(new_n438_));
  OR3_X1    g237(.A1(new_n435_), .A2(new_n436_), .A3(new_n389_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT21), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G197gat), .A2(G204gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(G197gat), .A2(G204gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n441_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G197gat), .ZN(new_n446_));
  INV_X1    g245(.A(G204gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(KEYINPUT21), .A3(new_n442_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G211gat), .B(G218gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n445_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n443_), .A2(new_n444_), .A3(new_n441_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G211gat), .B(G218gat), .Z(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n410_), .A2(new_n455_), .A3(new_n426_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n406_), .A2(KEYINPUT24), .A3(new_n399_), .A4(new_n408_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n412_), .A2(KEYINPUT25), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT25), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G183gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n413_), .A2(KEYINPUT26), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT26), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G190gat), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n458_), .A2(new_n460_), .A3(new_n461_), .A4(new_n463_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n402_), .A2(new_n457_), .A3(new_n411_), .A4(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n425_), .A2(new_n422_), .A3(new_n418_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n451_), .A2(new_n454_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n456_), .A2(new_n469_), .A3(KEYINPUT20), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G226gat), .A2(G233gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT19), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n427_), .A2(new_n468_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n472_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n455_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n474_), .A2(KEYINPUT20), .A3(new_n475_), .A4(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G8gat), .B(G36gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT18), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G64gat), .B(G92gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n473_), .A2(new_n477_), .A3(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n470_), .A2(new_n472_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n474_), .A2(KEYINPUT20), .A3(new_n476_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n472_), .B2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(KEYINPUT27), .B(new_n482_), .C1(new_n485_), .C2(new_n481_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n473_), .A2(new_n477_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n481_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT97), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n482_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT27), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n487_), .A2(KEYINPUT97), .A3(new_n488_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n495_));
  INV_X1    g294(.A(KEYINPUT92), .ZN(new_n496_));
  INV_X1    g295(.A(G155gat), .ZN(new_n497_));
  INV_X1    g296(.A(G162gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT92), .B1(G155gat), .B2(G162gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G155gat), .A2(G162gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G141gat), .ZN(new_n504_));
  INV_X1    g303(.A(G148gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(KEYINPUT3), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT3), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(G141gat), .B2(G148gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n509_), .A2(new_n512_), .A3(KEYINPUT94), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT94), .B1(new_n509_), .B2(new_n512_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n503_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G141gat), .A2(G148gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(G141gat), .A2(G148gat), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n501_), .A2(KEYINPUT1), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n499_), .A2(new_n520_), .A3(new_n500_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT93), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n499_), .A2(new_n520_), .A3(KEYINPUT93), .A4(new_n500_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n501_), .A2(KEYINPUT1), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n519_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n515_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n495_), .B1(new_n528_), .B2(KEYINPUT29), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT29), .ZN(new_n530_));
  INV_X1    g329(.A(new_n495_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n515_), .A2(new_n527_), .A3(new_n530_), .A4(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G22gat), .B(G50gat), .Z(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G78gat), .B(G106gat), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n534_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n529_), .A2(new_n538_), .A3(new_n532_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT96), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n536_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n535_), .B2(new_n539_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n528_), .A2(KEYINPUT29), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n468_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G228gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n541_), .A2(new_n544_), .A3(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n546_), .B(new_n547_), .Z(new_n550_));
  INV_X1    g349(.A(new_n539_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n538_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n542_), .B(new_n536_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n550_), .B1(new_n553_), .B2(new_n540_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n486_), .B(new_n494_), .C1(new_n549_), .C2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G1gat), .B(G29gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G57gat), .B(G85gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n519_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n524_), .A2(new_n525_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n521_), .A2(new_n522_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT94), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n506_), .A2(new_n508_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT2), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n516_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n565_), .B1(new_n566_), .B2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n509_), .A2(new_n512_), .A3(KEYINPUT94), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n502_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n388_), .B1(new_n564_), .B2(new_n573_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n382_), .A2(new_n387_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(new_n515_), .A3(new_n527_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(KEYINPUT4), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT98), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT98), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n574_), .A2(new_n579_), .A3(KEYINPUT4), .A4(new_n576_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT4), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n528_), .A2(new_n582_), .A3(new_n388_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G225gat), .A2(G233gat), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n581_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n574_), .A2(new_n576_), .A3(new_n584_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT100), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT100), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n574_), .A2(new_n591_), .A3(new_n576_), .A4(new_n584_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n560_), .B1(new_n588_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n560_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n586_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n555_), .A2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n548_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n553_), .A2(new_n550_), .A3(new_n540_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n604_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n491_), .A2(new_n493_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n560_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n604_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n588_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n581_), .A2(new_n584_), .A3(new_n583_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n574_), .A2(new_n576_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n560_), .B1(new_n612_), .B2(new_n585_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n605_), .A2(new_n606_), .A3(new_n610_), .A4(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n481_), .A2(KEYINPUT32), .ZN(new_n616_));
  MUX2_X1   g415(.A(new_n485_), .B(new_n487_), .S(new_n616_), .Z(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n603_), .B1(new_n615_), .B2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n440_), .B1(new_n600_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n494_), .A2(new_n486_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n549_), .A2(new_n554_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n598_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n620_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n321_), .A2(new_n373_), .A3(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT102), .Z(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(new_n203_), .A3(new_n599_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n615_), .A2(new_n618_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n623_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n622_), .A2(new_n598_), .A3(new_n603_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n626_), .B1(new_n637_), .B2(new_n440_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n370_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT103), .ZN(new_n640_));
  INV_X1    g439(.A(new_n320_), .ZN(new_n641_));
  AND4_X1   g440(.A1(new_n335_), .A2(new_n640_), .A3(new_n641_), .A4(new_n239_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n203_), .B1(new_n642_), .B2(new_n599_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n633_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n644_), .B1(new_n632_), .B2(new_n631_), .ZN(G1324gat));
  NAND3_X1  g444(.A1(new_n630_), .A2(new_n202_), .A3(new_n621_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n642_), .A2(new_n621_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  AND4_X1   g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .A4(G8gat), .ZN(new_n650_));
  INV_X1    g449(.A(G8gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(KEYINPUT104), .B2(KEYINPUT39), .ZN(new_n652_));
  AOI22_X1  g451(.A1(new_n648_), .A2(new_n652_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n646_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(G1325gat));
  INV_X1    g455(.A(new_n440_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n432_), .B1(new_n642_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT41), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n630_), .A2(new_n432_), .A3(new_n657_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1326gat));
  INV_X1    g460(.A(G22gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n642_), .B2(new_n603_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT42), .Z(new_n664_));
  NAND3_X1  g463(.A1(new_n630_), .A2(new_n662_), .A3(new_n603_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1327gat));
  INV_X1    g465(.A(new_n370_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n335_), .A2(new_n667_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n321_), .A2(new_n628_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G29gat), .B1(new_n669_), .B2(new_n599_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n657_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n671_), .B(new_n372_), .C1(new_n672_), .C2(new_n626_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n628_), .A2(KEYINPUT105), .A3(new_n671_), .A4(new_n372_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n372_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n638_), .B2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(new_n676_), .A3(new_n678_), .ZN(new_n679_));
  AND4_X1   g478(.A1(new_n336_), .A2(new_n317_), .A3(new_n319_), .A4(new_n239_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(KEYINPUT44), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT44), .B1(new_n679_), .B2(new_n680_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n599_), .A2(G29gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n670_), .B1(new_n683_), .B2(new_n684_), .ZN(G1328gat));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n622_), .A2(G36gat), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n321_), .A2(new_n628_), .A3(new_n668_), .A4(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT45), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n681_), .A2(new_n682_), .A3(new_n622_), .ZN(new_n692_));
  INV_X1    g491(.A(G36gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT106), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n682_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n679_), .A2(KEYINPUT44), .A3(new_n680_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n621_), .A3(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(G36gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n691_), .B1(new_n694_), .B2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n686_), .B(new_n687_), .C1(new_n700_), .C2(KEYINPUT107), .ZN(new_n701_));
  INV_X1    g500(.A(new_n691_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n692_), .A2(KEYINPUT106), .A3(new_n693_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n698_), .B1(new_n697_), .B2(G36gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT108), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT46), .B1(new_n700_), .B2(new_n686_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n701_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(G1329gat));
  NAND3_X1  g509(.A1(new_n683_), .A2(G43gat), .A3(new_n657_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n669_), .A2(new_n657_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(G43gat), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g513(.A(G50gat), .B1(new_n669_), .B2(new_n603_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n603_), .A2(G50gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n683_), .B2(new_n716_), .ZN(G1331gat));
  NOR2_X1   g516(.A1(new_n638_), .A2(new_n239_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n373_), .A2(new_n320_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(G57gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n599_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n240_), .A2(new_n336_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n640_), .A2(new_n320_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n599_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n725_), .B2(new_n720_), .ZN(G1332gat));
  INV_X1    g525(.A(G64gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n723_), .B2(new_n621_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT48), .Z(new_n729_));
  NAND3_X1  g528(.A1(new_n719_), .A2(new_n727_), .A3(new_n621_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1333gat));
  INV_X1    g530(.A(G71gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n723_), .B2(new_n657_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT49), .Z(new_n734_));
  NAND3_X1  g533(.A1(new_n719_), .A2(new_n732_), .A3(new_n657_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1334gat));
  INV_X1    g535(.A(G78gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n723_), .B2(new_n603_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT50), .Z(new_n739_));
  NAND2_X1  g538(.A1(new_n603_), .A2(new_n737_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT109), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n719_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(G1335gat));
  INV_X1    g542(.A(new_n239_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n320_), .A2(new_n336_), .A3(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT110), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n679_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n598_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n320_), .A2(new_n668_), .A3(new_n718_), .ZN(new_n749_));
  INV_X1    g548(.A(G85gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n599_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1336gat));
  OAI21_X1  g551(.A(G92gat), .B1(new_n747_), .B2(new_n622_), .ZN(new_n753_));
  INV_X1    g552(.A(G92gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n749_), .A2(new_n754_), .A3(new_n621_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1337gat));
  OAI21_X1  g555(.A(G99gat), .B1(new_n747_), .B2(new_n440_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n749_), .A2(new_n254_), .A3(new_n657_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g559(.A1(new_n749_), .A2(new_n255_), .A3(new_n603_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n746_), .A2(new_n603_), .A3(new_n679_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G106gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G106gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g566(.A1(new_n624_), .A2(new_n598_), .A3(new_n440_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT115), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n291_), .A2(new_n770_), .A3(new_n293_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n285_), .A2(new_n290_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n293_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT112), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n294_), .B1(new_n771_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n776_), .A2(KEYINPUT55), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(KEYINPUT55), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n300_), .B2(new_n778_), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n776_), .B(KEYINPUT55), .C1(new_n291_), .C2(new_n299_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n775_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT56), .B1(new_n781_), .B2(new_n246_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n218_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n224_), .B1(new_n230_), .B2(KEYINPUT113), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n214_), .A2(new_n229_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n235_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n783_), .A2(new_n788_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n238_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  INV_X1    g590(.A(new_n246_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n300_), .A2(new_n778_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n777_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n300_), .A2(new_n778_), .A3(new_n777_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n791_), .B(new_n792_), .C1(new_n797_), .C2(new_n775_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n306_), .A2(new_n307_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n782_), .A2(new_n790_), .A3(new_n798_), .A4(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n769_), .B1(new_n802_), .B2(new_n677_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n800_), .A2(new_n801_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n677_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(KEYINPUT115), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT116), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n239_), .A2(new_n782_), .A3(new_n799_), .A4(new_n798_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n238_), .A2(new_n789_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n812_), .A2(new_n308_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n810_), .B1(new_n814_), .B2(new_n667_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n810_), .B1(KEYINPUT116), .B2(new_n809_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n370_), .B(new_n816_), .C1(new_n811_), .C2(new_n813_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n335_), .B1(new_n807_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n372_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n722_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n820_), .B1(new_n722_), .B2(new_n821_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n768_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n819_), .A2(new_n824_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n825_), .B(new_n826_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n829_));
  OAI221_X1 g628(.A(new_n768_), .B1(KEYINPUT118), .B2(KEYINPUT59), .C1(new_n819_), .C2(new_n824_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G113gat), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n241_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n239_), .B(new_n768_), .C1(new_n819_), .C2(new_n824_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n832_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n835_), .A3(new_n832_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n834_), .A2(new_n840_), .A3(KEYINPUT119), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n836_), .A2(new_n835_), .A3(new_n832_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n837_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n833_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n842_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n841_), .A2(new_n847_), .ZN(G1340gat));
  OR2_X1    g647(.A1(new_n819_), .A2(new_n824_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT60), .ZN(new_n850_));
  AOI21_X1  g649(.A(G120gat), .B1(new_n320_), .B2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n850_), .B2(G120gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n849_), .A2(new_n768_), .A3(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT120), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n641_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n855_));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n855_), .B2(new_n856_), .ZN(G1341gat));
  INV_X1    g656(.A(new_n825_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n378_), .A3(new_n335_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n336_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n378_), .ZN(G1342gat));
  NAND3_X1  g660(.A1(new_n858_), .A2(new_n376_), .A3(new_n370_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n677_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n376_), .ZN(G1343gat));
  NOR4_X1   g663(.A1(new_n827_), .A2(new_n598_), .A3(new_n555_), .A4(new_n657_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n239_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n320_), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT121), .B(G148gat), .Z(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1345gat));
  NAND2_X1  g669(.A1(new_n865_), .A2(new_n335_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  NAND3_X1  g672(.A1(new_n865_), .A2(new_n498_), .A3(new_n370_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n865_), .A2(new_n372_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n874_), .B1(new_n876_), .B2(new_n498_), .ZN(G1347gat));
  NOR3_X1   g676(.A1(new_n625_), .A2(new_n603_), .A3(new_n622_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n849_), .A2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G169gat), .B1(new_n879_), .B2(new_n744_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n880_), .A2(KEYINPUT62), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n880_), .A2(KEYINPUT62), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n239_), .A2(new_n424_), .A3(new_n423_), .ZN(new_n883_));
  XOR2_X1   g682(.A(new_n883_), .B(KEYINPUT122), .Z(new_n884_));
  OAI22_X1  g683(.A1(new_n881_), .A2(new_n882_), .B1(new_n879_), .B2(new_n884_), .ZN(G1348gat));
  INV_X1    g684(.A(new_n879_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n320_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n335_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n391_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n412_), .B2(new_n889_), .ZN(G1350gat));
  NAND3_X1  g690(.A1(new_n886_), .A2(new_n370_), .A3(new_n392_), .ZN(new_n892_));
  OAI21_X1  g691(.A(G190gat), .B1(new_n879_), .B2(new_n677_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n893_), .A2(new_n894_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n892_), .B1(new_n895_), .B2(new_n896_), .ZN(G1351gat));
  NOR3_X1   g696(.A1(new_n657_), .A2(new_n623_), .A3(new_n599_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n899_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n900_), .A2(new_n901_), .A3(new_n622_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n849_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT125), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n849_), .A2(new_n905_), .A3(new_n902_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(G197gat), .B1(new_n907_), .B2(new_n239_), .ZN(new_n908_));
  AOI211_X1 g707(.A(new_n446_), .B(new_n744_), .C1(new_n904_), .C2(new_n906_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1352gat));
  INV_X1    g709(.A(new_n906_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n905_), .B1(new_n849_), .B2(new_n902_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n320_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G204gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n907_), .A2(new_n447_), .A3(new_n320_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1353gat));
  NOR2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n335_), .A2(new_n919_), .ZN(new_n920_));
  XOR2_X1   g719(.A(new_n920_), .B(KEYINPUT126), .Z(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n918_), .B1(new_n907_), .B2(new_n922_), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n917_), .B(new_n921_), .C1(new_n904_), .C2(new_n906_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1354gat));
  INV_X1    g724(.A(G218gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n907_), .A2(new_n926_), .A3(new_n370_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n677_), .B1(new_n904_), .B2(new_n906_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(G1355gat));
endmodule


