//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n933_, new_n934_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n963_, new_n964_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n980_,
    new_n981_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n989_, new_n990_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT36), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT77), .ZN(new_n206_));
  AND3_X1   g005(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G99gat), .ZN(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT65), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT7), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT7), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n214_), .A2(new_n210_), .A3(new_n211_), .A4(KEYINPUT65), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n209_), .A2(new_n213_), .A3(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G85gat), .B(G92gat), .Z(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(KEYINPUT66), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n216_), .A2(new_n217_), .A3(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n220_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT69), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n216_), .A2(new_n217_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n219_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT69), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n216_), .A2(new_n217_), .A3(new_n220_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(KEYINPUT10), .B(G99gat), .Z(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT64), .B(G106gat), .Z(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n217_), .A2(KEYINPUT9), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT9), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(G85gat), .A3(G92gat), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n232_), .A2(new_n233_), .A3(new_n235_), .A4(new_n209_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n229_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT15), .ZN(new_n238_));
  XOR2_X1   g037(.A(G29gat), .B(G36gat), .Z(new_n239_));
  XOR2_X1   g038(.A(G43gat), .B(G50gat), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT74), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G29gat), .B(G36gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G43gat), .B(G50gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(new_n242_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n242_), .B1(new_n241_), .B2(new_n245_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n238_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n248_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(KEYINPUT15), .A3(new_n246_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n237_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT75), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n241_), .A2(new_n245_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n236_), .B(new_n255_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(KEYINPUT34), .Z(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n253_), .A2(new_n254_), .A3(new_n256_), .A4(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n236_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(new_n223_), .B2(new_n228_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n249_), .A2(new_n251_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n254_), .B(new_n256_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n258_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n260_), .A2(KEYINPUT35), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n256_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(new_n237_), .B2(new_n252_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT35), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n265_), .B2(new_n260_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n206_), .B1(new_n266_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT76), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n266_), .A2(new_n271_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n260_), .A2(new_n265_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n270_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n260_), .A2(new_n265_), .A3(KEYINPUT35), .ZN(new_n280_));
  AND4_X1   g079(.A1(new_n273_), .A2(new_n279_), .A3(new_n280_), .A4(new_n275_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n272_), .B1(new_n276_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT78), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(KEYINPUT37), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(KEYINPUT37), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n274_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n279_), .A2(new_n280_), .A3(new_n275_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT76), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n291_), .A2(new_n283_), .A3(KEYINPUT37), .A4(new_n272_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G15gat), .B(G22gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G1gat), .A2(G8gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT14), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G1gat), .B(G8gat), .Z(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G231gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G57gat), .B(G64gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT11), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT67), .B(G71gat), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n302_), .A2(new_n303_), .B1(new_n304_), .B2(G78gat), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n304_), .A2(G78gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT68), .B1(new_n302_), .B2(new_n303_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n301_), .A2(new_n309_), .A3(KEYINPUT11), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n305_), .A2(new_n308_), .A3(new_n306_), .A4(new_n310_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n300_), .B(new_n314_), .Z(new_n315_));
  XNOR2_X1  g114(.A(G127gat), .B(G155gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT16), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G183gat), .ZN(new_n318_));
  INV_X1    g117(.A(G211gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT17), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n320_), .A2(new_n321_), .ZN(new_n323_));
  OR3_X1    g122(.A1(new_n315_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n315_), .A2(new_n323_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n287_), .A2(new_n292_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(G169gat), .ZN(new_n331_));
  INV_X1    g130(.A(G176gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT22), .B(G169gat), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n334_), .B2(new_n332_), .ZN(new_n335_));
  INV_X1    g134(.A(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT81), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(G190gat), .ZN(new_n339_));
  INV_X1    g138(.A(G183gat), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n337_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n342_), .B1(new_n340_), .B2(new_n336_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n335_), .B1(new_n341_), .B2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n337_), .A2(new_n339_), .A3(KEYINPUT26), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n336_), .A2(KEYINPUT26), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT25), .B(G183gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT82), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT82), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n347_), .A2(new_n352_), .A3(new_n348_), .A4(new_n349_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT83), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT83), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n356_), .B1(G169gat), .B2(G176gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT24), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(G169gat), .B2(G176gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n351_), .A2(new_n353_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n358_), .A2(new_n360_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n343_), .A2(new_n344_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(KEYINPUT84), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT84), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT24), .B1(new_n355_), .B2(new_n357_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n368_), .B2(new_n345_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n346_), .B1(new_n363_), .B2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT30), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT86), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G127gat), .B(G134gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G113gat), .B(G120gat), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n376_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT31), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT85), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n380_), .B2(new_n379_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G227gat), .A2(G233gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n382_), .B(new_n383_), .Z(new_n384_));
  XNOR2_X1  g183(.A(G71gat), .B(G99gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n382_), .B(new_n383_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n385_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G15gat), .B(G43gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n386_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n374_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n389_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n387_), .A2(new_n388_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n390_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n373_), .A3(new_n392_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G155gat), .A2(G162gat), .ZN(new_n401_));
  NOR2_X1   g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(KEYINPUT1), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT88), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT1), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n406_), .B1(G155gat), .B2(G162gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(KEYINPUT88), .A3(new_n401_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n401_), .A2(KEYINPUT1), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n405_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412_));
  INV_X1    g211(.A(G141gat), .ZN(new_n413_));
  INV_X1    g212(.A(G148gat), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n413_), .A2(new_n414_), .A3(KEYINPUT87), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT87), .B1(new_n413_), .B2(new_n414_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n412_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n411_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n377_), .A2(KEYINPUT92), .A3(new_n378_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT92), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n375_), .A2(new_n376_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n375_), .A2(new_n376_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  OR2_X1    g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n401_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n413_), .A2(new_n414_), .A3(KEYINPUT3), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT3), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(G141gat), .B2(G148gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n426_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n419_), .A2(new_n420_), .A3(new_n424_), .A4(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n409_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n417_), .B1(new_n437_), .B2(new_n408_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n421_), .B(new_n379_), .C1(new_n438_), .C2(new_n434_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G225gat), .A2(G233gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G1gat), .B(G29gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G57gat), .B(G85gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n440_), .A2(KEYINPUT4), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n441_), .B(KEYINPUT93), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n434_), .B1(new_n411_), .B2(new_n418_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n377_), .A2(new_n454_), .A3(new_n378_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT94), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n422_), .A2(new_n423_), .A3(KEYINPUT4), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT94), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n457_), .B(new_n458_), .C1(new_n438_), .C2(new_n434_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n452_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n450_), .A2(new_n460_), .A3(KEYINPUT95), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT95), .B1(new_n450_), .B2(new_n460_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n449_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT95), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n407_), .A2(KEYINPUT88), .A3(new_n401_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT88), .B1(new_n407_), .B2(new_n401_), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n409_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n435_), .B1(new_n467_), .B2(new_n417_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n458_), .B1(new_n468_), .B2(new_n457_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n453_), .A2(KEYINPUT94), .A3(new_n455_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n451_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n454_), .B1(new_n436_), .B2(new_n439_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n464_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n450_), .A2(new_n460_), .A3(KEYINPUT95), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n473_), .A2(new_n474_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n463_), .B1(new_n475_), .B2(new_n447_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n400_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT18), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(G64gat), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n481_), .A2(G92gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(G92gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G226gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT19), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n350_), .A2(KEYINPUT82), .B1(new_n359_), .B2(new_n361_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n488_), .A2(new_n353_), .A3(new_n369_), .A4(new_n366_), .ZN(new_n489_));
  INV_X1    g288(.A(G218gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G211gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n319_), .A2(G218gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT21), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G197gat), .B(G204gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n491_), .A2(new_n492_), .A3(KEYINPUT21), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n495_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n496_), .A2(KEYINPUT21), .A3(new_n491_), .A4(new_n492_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT89), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n499_), .A2(KEYINPUT89), .A3(new_n500_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n489_), .B(new_n346_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT20), .ZN(new_n504_));
  NOR2_X1   g303(.A1(G183gat), .A2(G190gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n335_), .B1(new_n345_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT26), .B(G190gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n349_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n354_), .A2(new_n360_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n365_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT91), .B1(new_n333_), .B2(new_n360_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n361_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n358_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n506_), .B1(new_n510_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n499_), .A2(new_n500_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n504_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n487_), .B1(new_n503_), .B2(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(KEYINPUT20), .B(new_n487_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n502_), .A2(new_n501_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n371_), .B2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n484_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n517_), .B1(new_n371_), .B2(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n486_), .ZN(new_n524_));
  INV_X1    g323(.A(G92gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n481_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n519_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n371_), .A2(new_n520_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n526_), .A3(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n522_), .A2(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n531_), .A2(KEYINPUT27), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT20), .B1(new_n515_), .B2(new_n516_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT98), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(KEYINPUT98), .B(KEYINPUT20), .C1(new_n515_), .C2(new_n516_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n528_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(new_n486_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n486_), .B2(new_n523_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n484_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(KEYINPUT27), .A3(new_n530_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n532_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G78gat), .B(G106gat), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n468_), .A2(KEYINPUT29), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n516_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(G228gat), .A3(G233gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G228gat), .A2(G233gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n545_), .A2(new_n520_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n544_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT28), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n468_), .B2(KEYINPUT29), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT29), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n453_), .A2(KEYINPUT28), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G22gat), .B(G50gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT90), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n560_), .B1(new_n550_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n553_), .A2(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n551_), .A2(new_n561_), .A3(new_n552_), .A4(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n542_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n478_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n448_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n569_), .B1(new_n570_), .B2(KEYINPUT33), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT33), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n463_), .A2(KEYINPUT97), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(KEYINPUT33), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n447_), .B1(new_n440_), .B2(new_n451_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n441_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n575_), .B1(new_n576_), .B2(new_n472_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n522_), .A2(new_n530_), .A3(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n571_), .A2(new_n573_), .A3(new_n574_), .A4(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n524_), .A2(new_n529_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n482_), .A2(KEYINPUT32), .A3(new_n483_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n539_), .B2(new_n581_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n476_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n579_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n566_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT99), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n565_), .B1(new_n579_), .B2(new_n584_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT99), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n532_), .A2(new_n565_), .A3(new_n477_), .A4(new_n541_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n588_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n400_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n568_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n237_), .A2(KEYINPUT12), .A3(new_n314_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n236_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n314_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT12), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n314_), .A2(new_n596_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n597_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n595_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n599_), .ZN(new_n603_));
  OAI211_X1 g402(.A(G230gat), .B(G233gat), .C1(new_n603_), .C2(new_n597_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT71), .ZN(new_n606_));
  XOR2_X1   g405(.A(G120gat), .B(G148gat), .Z(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  XNOR2_X1  g407(.A(G176gat), .B(G204gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n602_), .A2(new_n604_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT72), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT72), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n602_), .A2(new_n613_), .A3(new_n604_), .A4(new_n610_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n602_), .A2(new_n604_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n610_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(KEYINPUT13), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(KEYINPUT13), .B1(new_n615_), .B2(new_n618_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n620_), .A2(KEYINPUT73), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT73), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n615_), .A2(new_n618_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT13), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n623_), .B1(new_n626_), .B2(new_n619_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n622_), .A2(new_n627_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n263_), .A2(new_n298_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n298_), .A2(new_n255_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G229gat), .A2(G233gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n629_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n298_), .B(new_n255_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n631_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G113gat), .B(G141gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(G169gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(G197gat), .Z(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n640_), .A2(KEYINPUT80), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n636_), .B(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n628_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n594_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n330_), .A2(new_n644_), .ZN(new_n645_));
  OR3_X1    g444(.A1(new_n645_), .A2(G1gat), .A3(new_n477_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT38), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n591_), .B1(new_n589_), .B2(KEYINPUT99), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n587_), .B(new_n565_), .C1(new_n579_), .C2(new_n584_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n593_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n478_), .A2(new_n567_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT100), .B1(new_n652_), .B2(new_n282_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654_));
  INV_X1    g453(.A(new_n274_), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n288_), .A2(new_n290_), .B1(new_n655_), .B2(new_n206_), .ZN(new_n656_));
  AOI211_X1 g455(.A(new_n654_), .B(new_n656_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n653_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n643_), .A2(new_n326_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n476_), .A3(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(KEYINPUT101), .A3(G1gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT101), .B1(new_n660_), .B2(G1gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n647_), .B1(new_n661_), .B2(new_n662_), .ZN(G1324gat));
  OR3_X1    g462(.A1(new_n645_), .A2(G8gat), .A3(new_n542_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n542_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n665_), .B(new_n659_), .C1(new_n653_), .C2(new_n657_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n666_), .A2(new_n667_), .A3(G8gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n666_), .B2(G8gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n664_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(G1325gat));
  OR3_X1    g471(.A1(new_n645_), .A2(G15gat), .A3(new_n593_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n658_), .A2(new_n400_), .A3(new_n659_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n674_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT41), .B1(new_n674_), .B2(G15gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n675_), .B2(new_n676_), .ZN(G1326gat));
  OR3_X1    g476(.A1(new_n645_), .A2(G22gat), .A3(new_n566_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n658_), .A2(new_n565_), .A3(new_n659_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G22gat), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(KEYINPUT42), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(KEYINPUT42), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(G1327gat));
  INV_X1    g482(.A(new_n642_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n622_), .A2(new_n627_), .A3(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n282_), .A2(new_n327_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n652_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT102), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n652_), .A2(new_n685_), .A3(new_n689_), .A4(new_n686_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n476_), .ZN(new_n692_));
  INV_X1    g491(.A(G29gat), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n685_), .A2(new_n326_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n287_), .A2(new_n292_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT43), .B1(new_n594_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n652_), .A2(new_n699_), .A3(new_n696_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n695_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT44), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(G29gat), .A3(new_n476_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n701_), .A2(KEYINPUT44), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n694_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n694_), .B(KEYINPUT103), .C1(new_n703_), .C2(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1328gat));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710_));
  INV_X1    g509(.A(G36gat), .ZN(new_n711_));
  INV_X1    g510(.A(new_n704_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n542_), .B1(new_n701_), .B2(KEYINPUT44), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n711_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n688_), .A2(new_n711_), .A3(new_n665_), .A4(new_n690_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT105), .Z(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n715_), .B(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n710_), .B1(new_n714_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n702_), .A2(new_n665_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G36gat), .B1(new_n721_), .B2(new_n704_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n715_), .B(new_n717_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(KEYINPUT46), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n720_), .A2(new_n724_), .ZN(G1329gat));
  NAND2_X1  g524(.A1(new_n691_), .A2(new_n400_), .ZN(new_n726_));
  INV_X1    g525(.A(G43gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n702_), .A2(G43gat), .A3(new_n400_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n704_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n728_), .B(new_n731_), .C1(new_n729_), .C2(new_n704_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1330gat));
  AOI21_X1  g534(.A(G50gat), .B1(new_n691_), .B2(new_n565_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n702_), .A2(G50gat), .A3(new_n565_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n712_), .ZN(G1331gat));
  NAND2_X1  g537(.A1(new_n652_), .A2(new_n684_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n628_), .B1(new_n739_), .B2(KEYINPUT107), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n652_), .A2(new_n741_), .A3(new_n684_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n740_), .A2(new_n330_), .A3(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT108), .ZN(new_n744_));
  INV_X1    g543(.A(new_n742_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n628_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n642_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(new_n741_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n745_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n330_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n477_), .A2(G57gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n744_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n684_), .A2(new_n327_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n628_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n658_), .A2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G57gat), .B1(new_n756_), .B2(new_n477_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n753_), .A2(new_n757_), .ZN(G1332gat));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n542_), .A2(G64gat), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n744_), .A2(new_n751_), .A3(new_n760_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n665_), .B(new_n755_), .C1(new_n653_), .C2(new_n657_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G64gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G64gat), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n759_), .B1(new_n761_), .B2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n744_), .A2(new_n751_), .A3(new_n760_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(KEYINPUT109), .C1(new_n765_), .C2(new_n764_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1333gat));
  NOR2_X1   g569(.A1(new_n593_), .A2(G71gat), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT110), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n744_), .A2(new_n751_), .A3(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G71gat), .B1(new_n756_), .B2(new_n593_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(KEYINPUT49), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(KEYINPUT49), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n773_), .B1(new_n775_), .B2(new_n776_), .ZN(G1334gat));
  NOR2_X1   g576(.A1(new_n566_), .A2(G78gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n744_), .A2(new_n751_), .A3(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G78gat), .B1(new_n756_), .B2(new_n566_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(KEYINPUT50), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(KEYINPUT50), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n779_), .B1(new_n781_), .B2(new_n782_), .ZN(G1335gat));
  OAI21_X1  g582(.A(KEYINPUT107), .B1(new_n594_), .B2(new_n642_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n784_), .A2(new_n746_), .A3(new_n686_), .A4(new_n742_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G85gat), .B1(new_n786_), .B2(new_n476_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n327_), .A2(new_n642_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n622_), .B2(new_n627_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT111), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n788_), .C1(new_n622_), .C2(new_n627_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n698_), .A2(new_n700_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n476_), .A2(G85gat), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT112), .Z(new_n795_));
  AOI21_X1  g594(.A(new_n787_), .B1(new_n793_), .B2(new_n795_), .ZN(G1336gat));
  NAND3_X1  g595(.A1(new_n793_), .A2(G92gat), .A3(new_n665_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n798_), .B(new_n525_), .C1(new_n785_), .C2(new_n542_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n740_), .A2(new_n665_), .A3(new_n686_), .A4(new_n742_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n798_), .B1(new_n801_), .B2(new_n525_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n797_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT114), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n797_), .B(new_n805_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1337gat));
  NAND2_X1  g606(.A1(new_n790_), .A2(new_n792_), .ZN(new_n808_));
  AOI221_X4 g607(.A(KEYINPUT43), .B1(new_n287_), .B2(new_n292_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n699_), .B1(new_n652_), .B2(new_n696_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n400_), .B(new_n808_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n811_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT115), .B1(new_n811_), .B2(G99gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT117), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n400_), .A2(new_n230_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n749_), .A2(KEYINPUT116), .A3(new_n686_), .A4(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n785_), .B2(new_n815_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT51), .B1(new_n814_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n811_), .A2(G99gat), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n811_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n817_), .A2(new_n819_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n826_), .A2(KEYINPUT117), .A3(new_n827_), .A4(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n821_), .A2(new_n829_), .ZN(G1338gat));
  NAND3_X1  g629(.A1(new_n786_), .A2(new_n565_), .A3(new_n231_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n565_), .B(new_n808_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n832_), .A2(new_n833_), .A3(G106gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(G106gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT53), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n831_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1339gat));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n593_), .A2(new_n567_), .A3(new_n477_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(KEYINPUT122), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(KEYINPUT122), .B2(new_n842_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n601_), .B1(new_n595_), .B2(new_n600_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n602_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n595_), .A2(new_n600_), .A3(KEYINPUT55), .A4(new_n601_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT56), .B1(new_n849_), .B2(new_n617_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n851_), .B(new_n610_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n615_), .B(new_n642_), .C1(new_n850_), .C2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n629_), .A2(new_n630_), .A3(new_n634_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n639_), .B1(new_n633_), .B2(new_n631_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n854_), .A2(KEYINPUT118), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT118), .B1(new_n854_), .B2(new_n855_), .ZN(new_n857_));
  OAI22_X1  g656(.A1(new_n856_), .A2(new_n857_), .B1(new_n640_), .B2(new_n636_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n624_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n656_), .B1(new_n853_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT57), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT121), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(new_n864_), .A3(KEYINPUT57), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n858_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n866_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n850_), .A2(new_n852_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n871_), .A2(KEYINPUT120), .A3(KEYINPUT58), .A4(new_n867_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n868_), .A2(new_n869_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n870_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n863_), .A2(new_n865_), .B1(new_n874_), .B2(new_n696_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n853_), .A2(new_n860_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n656_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n327_), .B1(new_n875_), .B2(new_n878_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n620_), .A2(new_n754_), .A3(new_n621_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n697_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT54), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n697_), .A2(new_n883_), .A3(new_n880_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n844_), .B1(new_n879_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n842_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n865_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n864_), .B1(new_n861_), .B2(KEYINPUT57), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n870_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n890_));
  OAI22_X1  g689(.A1(new_n888_), .A2(new_n889_), .B1(new_n890_), .B2(new_n697_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n892_), .B(new_n876_), .C1(new_n877_), .C2(new_n656_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT119), .B1(new_n861_), .B2(KEYINPUT57), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n326_), .B1(new_n891_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n882_), .A2(new_n884_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n887_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n886_), .B(new_n642_), .C1(new_n898_), .C2(new_n841_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G113gat), .ZN(new_n900_));
  INV_X1    g699(.A(G113gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n898_), .A2(new_n901_), .A3(new_n642_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1340gat));
  OAI211_X1 g702(.A(new_n886_), .B(new_n746_), .C1(new_n898_), .C2(new_n841_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(G120gat), .ZN(new_n905_));
  INV_X1    g704(.A(G120gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(KEYINPUT60), .B1(new_n746_), .B2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(KEYINPUT60), .B2(new_n906_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n895_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n327_), .B1(new_n875_), .B2(new_n909_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n842_), .B(new_n908_), .C1(new_n910_), .C2(new_n885_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n898_), .A2(KEYINPUT123), .A3(new_n908_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n905_), .A2(new_n915_), .ZN(G1341gat));
  OAI211_X1 g715(.A(new_n886_), .B(new_n327_), .C1(new_n898_), .C2(new_n841_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(G127gat), .ZN(new_n918_));
  INV_X1    g717(.A(G127gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n898_), .A2(new_n919_), .A3(new_n327_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(G1342gat));
  OAI211_X1 g720(.A(new_n886_), .B(new_n696_), .C1(new_n898_), .C2(new_n841_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(G134gat), .ZN(new_n923_));
  INV_X1    g722(.A(G134gat), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n898_), .A2(new_n924_), .A3(new_n656_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1343gat));
  NAND2_X1  g725(.A1(new_n896_), .A2(new_n897_), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n665_), .A2(new_n400_), .A3(new_n477_), .A4(new_n566_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n927_), .A2(new_n642_), .A3(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g729(.A1(new_n927_), .A2(new_n746_), .A3(new_n928_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g731(.A1(new_n927_), .A2(new_n327_), .A3(new_n928_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(KEYINPUT61), .B(G155gat), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(G1346gat));
  AND4_X1   g734(.A1(G162gat), .A2(new_n927_), .A3(new_n696_), .A4(new_n928_), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n656_), .B(new_n928_), .C1(new_n910_), .C2(new_n885_), .ZN(new_n937_));
  INV_X1    g736(.A(G162gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n937_), .A2(KEYINPUT124), .A3(new_n938_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n936_), .B1(new_n941_), .B2(new_n942_), .ZN(G1347gat));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n944_));
  OAI221_X1 g743(.A(new_n878_), .B1(new_n697_), .B2(new_n890_), .C1(new_n888_), .C2(new_n889_), .ZN(new_n945_));
  AOI22_X1  g744(.A1(new_n945_), .A2(new_n326_), .B1(new_n882_), .B2(new_n884_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n478_), .A2(new_n542_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n947_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(new_n565_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n949_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n946_), .A2(new_n684_), .A3(new_n950_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n944_), .B1(new_n951_), .B2(new_n331_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n949_), .B1(new_n879_), .B2(new_n885_), .ZN(new_n953_));
  OAI211_X1 g752(.A(KEYINPUT62), .B(G169gat), .C1(new_n953_), .C2(new_n684_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n951_), .A2(new_n334_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n952_), .A2(new_n954_), .A3(new_n955_), .ZN(G1348gat));
  NOR2_X1   g755(.A1(new_n910_), .A2(new_n885_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n957_), .A2(new_n565_), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n628_), .A2(new_n948_), .A3(new_n332_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n332_), .B1(new_n953_), .B2(new_n628_), .ZN(new_n961_));
  AND2_X1   g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1349gat));
  NOR3_X1   g761(.A1(new_n953_), .A2(new_n349_), .A3(new_n326_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n958_), .A2(new_n327_), .A3(new_n947_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n963_), .B1(new_n964_), .B2(new_n340_), .ZN(G1350gat));
  OAI211_X1 g764(.A(new_n696_), .B(new_n949_), .C1(new_n879_), .C2(new_n885_), .ZN(new_n966_));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n967_));
  AND3_X1   g766(.A1(new_n966_), .A2(new_n967_), .A3(G190gat), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n967_), .B1(new_n966_), .B2(G190gat), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n656_), .A2(new_n507_), .ZN(new_n970_));
  OAI22_X1  g769(.A1(new_n968_), .A2(new_n969_), .B1(new_n953_), .B2(new_n970_), .ZN(G1351gat));
  NOR3_X1   g770(.A1(new_n400_), .A2(new_n476_), .A3(new_n566_), .ZN(new_n972_));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973_));
  OR2_X1    g772(.A1(new_n972_), .A2(new_n973_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n972_), .A2(new_n973_), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n974_), .A2(new_n665_), .A3(new_n975_), .ZN(new_n976_));
  INV_X1    g775(.A(new_n976_), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n927_), .A2(new_n642_), .A3(new_n977_), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n978_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g778(.A1(new_n927_), .A2(new_n746_), .A3(new_n977_), .ZN(new_n980_));
  XNOR2_X1  g779(.A(KEYINPUT127), .B(G204gat), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n980_), .B(new_n981_), .ZN(G1353gat));
  XNOR2_X1  g781(.A(KEYINPUT63), .B(G211gat), .ZN(new_n983_));
  NOR4_X1   g782(.A1(new_n957_), .A2(new_n326_), .A3(new_n976_), .A4(new_n983_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n957_), .A2(new_n976_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n985_), .A2(new_n327_), .ZN(new_n986_));
  NOR2_X1   g785(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n987_));
  AOI21_X1  g786(.A(new_n984_), .B1(new_n986_), .B2(new_n987_), .ZN(G1354gat));
  NAND3_X1  g787(.A1(new_n985_), .A2(new_n490_), .A3(new_n656_), .ZN(new_n989_));
  NOR3_X1   g788(.A1(new_n957_), .A2(new_n697_), .A3(new_n976_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n989_), .B1(new_n490_), .B2(new_n990_), .ZN(G1355gat));
endmodule


