//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n971_, new_n972_,
    new_n974_, new_n975_, new_n976_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n984_, new_n985_, new_n986_, new_n988_,
    new_n989_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT7), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT67), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT67), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n214_), .A2(new_n203_), .A3(new_n204_), .A4(new_n205_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n207_), .A2(new_n212_), .A3(new_n213_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n217_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT69), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n216_), .A2(new_n218_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT8), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT69), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n219_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT10), .B(G99gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n212_), .B1(new_n227_), .B2(G106gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT66), .B(G92gat), .ZN(new_n230_));
  INV_X1    g029(.A(G85gat), .ZN(new_n231_));
  AND2_X1   g030(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n232_));
  OAI22_X1  g031(.A1(KEYINPUT65), .A2(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n233_));
  OAI22_X1  g032(.A1(new_n230_), .A2(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n228_), .B1(new_n229_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n222_), .A2(new_n226_), .A3(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G57gat), .B(G64gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G71gat), .B(G78gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(KEYINPUT11), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n241_));
  INV_X1    g040(.A(new_n239_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n240_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n237_), .A2(KEYINPUT12), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G230gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT64), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n235_), .B1(new_n224_), .B2(new_n219_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n250_), .B1(new_n251_), .B2(new_n245_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n236_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(new_n246_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT12), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT70), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n257_));
  AOI211_X1 g056(.A(new_n257_), .B(KEYINPUT12), .C1(new_n253_), .C2(new_n246_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n247_), .B(new_n252_), .C1(new_n256_), .C2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n251_), .A2(new_n245_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n254_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT68), .B1(new_n251_), .B2(new_n245_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n250_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G120gat), .B(G148gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT5), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G176gat), .B(G204gat), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n266_), .B(new_n267_), .Z(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n259_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT71), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n259_), .B2(new_n264_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n259_), .A2(new_n264_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n268_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(KEYINPUT71), .A3(new_n270_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n273_), .A2(new_n276_), .A3(KEYINPUT13), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT13), .B1(new_n273_), .B2(new_n276_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n202_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n273_), .A2(new_n276_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT13), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(KEYINPUT72), .A3(new_n277_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G29gat), .B(G36gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT73), .ZN(new_n287_));
  XOR2_X1   g086(.A(G43gat), .B(G50gat), .Z(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT15), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT79), .B(G8gat), .ZN(new_n291_));
  INV_X1    g090(.A(G1gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT80), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT80), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n297_), .A3(new_n294_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G8gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n296_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n290_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n302_), .A2(new_n303_), .A3(new_n289_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G229gat), .A2(G233gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n306_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n289_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G113gat), .B(G141gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G169gat), .B(G197gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n308_), .A2(new_n312_), .A3(new_n316_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n285_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n290_), .A2(new_n237_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n251_), .A2(new_n289_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G232gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT34), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT35), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n326_), .A2(new_n327_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n322_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT77), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n322_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n323_), .A2(KEYINPUT74), .A3(new_n328_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n322_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n333_), .A2(new_n335_), .B1(new_n339_), .B2(new_n330_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G190gat), .B(G218gat), .Z(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT75), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G134gat), .B(G162gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n340_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n344_), .B(KEYINPUT36), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n347_), .B(KEYINPUT37), .C1(new_n340_), .C2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(new_n340_), .B2(new_n348_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n348_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n335_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n334_), .B1(new_n322_), .B2(new_n331_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n339_), .A2(new_n330_), .ZN(new_n357_));
  OAI211_X1 g156(.A(KEYINPUT78), .B(new_n353_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n352_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n347_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT37), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n350_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G231gat), .A2(G233gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n245_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(new_n303_), .A3(new_n302_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n304_), .A2(new_n364_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G127gat), .B(G155gat), .Z(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G183gat), .B(G211gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT17), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n369_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n369_), .A2(new_n375_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AOI211_X1 g177(.A(KEYINPUT17), .B(new_n374_), .C1(new_n366_), .C2(new_n368_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT83), .B1(new_n378_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n382_));
  AOI211_X1 g181(.A(new_n382_), .B(new_n379_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n362_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT93), .ZN(new_n386_));
  INV_X1    g185(.A(G204gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT89), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT89), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G204gat), .ZN(new_n390_));
  INV_X1    g189(.A(G197gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT21), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n393_), .B1(G197gat), .B2(G204gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(G218gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(G211gat), .ZN(new_n397_));
  INV_X1    g196(.A(G211gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G218gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n399_), .A3(KEYINPUT90), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT90), .B1(new_n397_), .B2(new_n399_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n395_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n389_), .A2(G204gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n387_), .A2(KEYINPUT89), .ZN(new_n405_));
  OAI21_X1  g204(.A(G197gat), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G197gat), .A2(G204gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT21), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n406_), .A2(KEYINPUT21), .A3(new_n408_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n397_), .A2(new_n399_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT90), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n400_), .ZN(new_n414_));
  OAI22_X1  g213(.A1(new_n403_), .A2(new_n409_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT91), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n391_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n393_), .B1(new_n418_), .B2(new_n407_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(new_n414_), .A3(new_n395_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n418_), .A2(new_n407_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n421_), .A2(KEYINPUT21), .A3(new_n400_), .A4(new_n413_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n422_), .A3(KEYINPUT91), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G228gat), .A2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  OR2_X1    g224(.A1(G155gat), .A2(G162gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G141gat), .A2(G148gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT2), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(KEYINPUT88), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n432_));
  INV_X1    g231(.A(G141gat), .ZN(new_n433_));
  INV_X1    g232(.A(G148gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n431_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n430_), .B1(new_n429_), .B2(KEYINPUT88), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n428_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n433_), .A2(new_n434_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n440_), .A2(new_n429_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT1), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n426_), .A2(new_n443_), .A3(new_n427_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n439_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n425_), .B1(new_n446_), .B2(KEYINPUT29), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n417_), .A2(new_n423_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(KEYINPUT29), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n415_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n425_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G78gat), .B(G106gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n448_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n448_), .B2(new_n451_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT92), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n448_), .A2(new_n451_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(new_n456_), .A3(new_n452_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT28), .B1(new_n446_), .B2(KEYINPUT29), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n429_), .A2(KEYINPUT88), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT2), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n462_), .A2(new_n431_), .A3(new_n435_), .A4(new_n436_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n463_), .A2(new_n428_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT28), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT29), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G22gat), .B(G50gat), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n460_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n468_), .B1(new_n460_), .B2(new_n467_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n459_), .A2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n386_), .B1(new_n457_), .B2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n471_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n458_), .A2(new_n452_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT92), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n475_), .B(KEYINPUT93), .C1(new_n477_), .C2(new_n454_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n453_), .A2(KEYINPUT94), .ZN(new_n480_));
  OAI221_X1 g279(.A(new_n471_), .B1(new_n458_), .B2(new_n480_), .C1(new_n476_), .C2(KEYINPUT94), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT27), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT100), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G226gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT19), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT99), .ZN(new_n487_));
  INV_X1    g286(.A(G190gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT26), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT26), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G190gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT25), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G183gat), .ZN(new_n493_));
  INV_X1    g292(.A(G183gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT25), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n489_), .A2(new_n491_), .A3(new_n493_), .A4(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(G169gat), .A2(G176gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G169gat), .A2(G176gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(KEYINPUT24), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT95), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G183gat), .A2(G190gat), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT23), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n504_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT96), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n504_), .A2(KEYINPUT96), .A3(new_n507_), .A4(new_n508_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT95), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n496_), .A2(new_n500_), .A3(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n502_), .A2(new_n511_), .A3(new_n512_), .A4(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT22), .B(G169gat), .ZN(new_n516_));
  INV_X1    g315(.A(G176gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT97), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n499_), .B(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n494_), .A2(new_n488_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n507_), .A2(new_n521_), .A3(KEYINPUT98), .A4(new_n508_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n518_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n507_), .A2(new_n508_), .A3(new_n521_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT98), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  AOI221_X4 g326(.A(new_n487_), .B1(new_n420_), .B2(new_n422_), .C1(new_n515_), .C2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n515_), .A2(new_n527_), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT99), .B1(new_n529_), .B2(new_n415_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT26), .B(G190gat), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT84), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT25), .B1(new_n533_), .B2(new_n494_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n492_), .A2(KEYINPUT84), .A3(G183gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n532_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT85), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT85), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n532_), .A2(new_n538_), .A3(new_n534_), .A4(new_n535_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  AND4_X1   g339(.A1(new_n507_), .A2(new_n500_), .A3(new_n508_), .A4(new_n504_), .ZN(new_n541_));
  INV_X1    g340(.A(G169gat), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT86), .B1(new_n542_), .B2(KEYINPUT22), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n517_), .B(new_n543_), .C1(new_n516_), .C2(KEYINPUT86), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n524_), .A2(new_n499_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n540_), .A2(new_n541_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n420_), .A2(new_n422_), .A3(KEYINPUT91), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT91), .B1(new_n420_), .B2(new_n422_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT20), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n484_), .B(new_n486_), .C1(new_n531_), .C2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT20), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n523_), .A2(new_n526_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n496_), .A2(new_n500_), .A3(new_n513_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n513_), .B1(new_n496_), .B2(new_n500_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n511_), .A2(new_n512_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n553_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n415_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n552_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n540_), .A2(new_n541_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n545_), .A2(new_n544_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n417_), .A2(new_n563_), .A3(new_n423_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(new_n486_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n551_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n487_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n529_), .A2(KEYINPUT99), .A3(new_n415_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n417_), .A2(new_n423_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n552_), .B1(new_n572_), .B2(new_n546_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n484_), .B1(new_n574_), .B2(new_n486_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G64gat), .B(G92gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT102), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G8gat), .B(G36gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n568_), .A2(new_n575_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n486_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n566_), .B1(new_n585_), .B2(new_n484_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n486_), .B1(new_n531_), .B2(new_n550_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT100), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n581_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n483_), .B1(new_n583_), .B2(new_n589_), .ZN(new_n590_));
  AOI211_X1 g389(.A(KEYINPUT104), .B(new_n584_), .C1(new_n560_), .C2(new_n564_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n571_), .A2(new_n573_), .A3(new_n584_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT104), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n565_), .B2(new_n486_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n591_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n483_), .B1(new_n595_), .B2(new_n582_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n586_), .A2(new_n581_), .A3(new_n588_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G71gat), .B(G99gat), .ZN(new_n599_));
  INV_X1    g398(.A(G43gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n546_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G127gat), .B(G134gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G113gat), .B(G120gat), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n604_), .A2(new_n605_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n603_), .B(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G227gat), .A2(G233gat), .ZN(new_n610_));
  INV_X1    g409(.A(G15gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT30), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT31), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n609_), .B(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n464_), .A2(new_n608_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n606_), .A2(new_n607_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n446_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(new_n618_), .A3(KEYINPUT4), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT4), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n446_), .A2(new_n620_), .A3(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G225gat), .A2(G233gat), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G1gat), .B(G29gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(G85gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT0), .B(G57gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n627_), .B(new_n628_), .Z(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n616_), .A2(new_n618_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n623_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n625_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n623_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n629_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n633_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(KEYINPUT105), .B(new_n629_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n615_), .A2(new_n640_), .ZN(new_n641_));
  AND4_X1   g440(.A1(new_n482_), .A2(new_n590_), .A3(new_n598_), .A4(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n582_), .B1(new_n568_), .B2(new_n575_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n636_), .A2(KEYINPUT33), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n645_), .B(new_n629_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n616_), .A2(new_n618_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n629_), .B1(new_n647_), .B2(new_n624_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n648_), .B1(new_n624_), .B2(new_n622_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT103), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n648_), .B(new_n651_), .C1(new_n624_), .C2(new_n622_), .ZN(new_n652_));
  AOI22_X1  g451(.A1(new_n644_), .A2(new_n646_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n643_), .A2(new_n597_), .A3(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n581_), .A2(KEYINPUT32), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n586_), .A2(new_n588_), .A3(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n581_), .A2(KEYINPUT32), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n595_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(new_n658_), .A3(new_n640_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n654_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n482_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n640_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n590_), .A2(new_n662_), .A3(new_n598_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n615_), .B(KEYINPUT87), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n642_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n321_), .A2(new_n385_), .A3(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(new_n292_), .A3(new_n640_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT38), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  AOI22_X1  g470(.A1(new_n352_), .A2(new_n358_), .B1(new_n340_), .B2(new_n346_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n667_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n320_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n280_), .B2(new_n284_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n673_), .A2(new_n384_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n640_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G1gat), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n669_), .A2(new_n670_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n671_), .A2(new_n678_), .A3(new_n679_), .ZN(G1324gat));
  NAND2_X1  g479(.A1(new_n643_), .A2(new_n597_), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n681_), .A2(new_n483_), .B1(new_n597_), .B2(new_n596_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n668_), .A2(new_n291_), .A3(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT106), .ZN(new_n685_));
  OAI21_X1  g484(.A(G8gat), .B1(new_n676_), .B2(new_n682_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT39), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n687_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n685_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n685_), .A2(KEYINPUT40), .A3(new_n688_), .A4(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1325gat));
  OAI21_X1  g493(.A(G15gat), .B1(new_n676_), .B2(new_n666_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT41), .Z(new_n696_));
  NAND3_X1  g495(.A1(new_n668_), .A2(new_n611_), .A3(new_n665_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1326gat));
  OAI21_X1  g497(.A(G22gat), .B1(new_n676_), .B2(new_n482_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT42), .ZN(new_n700_));
  INV_X1    g499(.A(G22gat), .ZN(new_n701_));
  INV_X1    g500(.A(new_n482_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n668_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(new_n703_), .ZN(G1327gat));
  NOR2_X1   g503(.A1(new_n321_), .A2(new_n667_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n360_), .A2(new_n384_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G29gat), .B1(new_n708_), .B2(new_n640_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n384_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n675_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n682_), .A2(new_n482_), .A3(new_n641_), .ZN(new_n714_));
  AOI22_X1  g513(.A1(new_n682_), .A2(new_n662_), .B1(new_n660_), .B2(new_n482_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(new_n665_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n349_), .B1(new_n672_), .B2(KEYINPUT37), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n665_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n713_), .B(new_n717_), .C1(new_n719_), .C2(new_n642_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n712_), .B1(new_n718_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n722_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT43), .B1(new_n667_), .B2(new_n362_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n711_), .B1(new_n726_), .B2(new_n720_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT107), .B1(new_n727_), .B2(KEYINPUT44), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(KEYINPUT44), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n640_), .A2(G29gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n709_), .B1(new_n731_), .B2(new_n732_), .ZN(G1328gat));
  INV_X1    g532(.A(KEYINPUT46), .ZN(new_n734_));
  INV_X1    g533(.A(G36gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n682_), .B1(new_n727_), .B2(KEYINPUT44), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n729_), .B2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n682_), .A2(G36gat), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n675_), .A2(new_n716_), .A3(new_n706_), .A4(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT108), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n739_), .A2(KEYINPUT108), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n739_), .A2(KEYINPUT108), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT45), .B1(new_n745_), .B2(new_n740_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n734_), .B1(new_n737_), .B2(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n744_), .A2(new_n746_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n730_), .A2(new_n683_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n728_), .B2(new_n725_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT46), .B(new_n749_), .C1(new_n751_), .C2(new_n735_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n748_), .A2(new_n752_), .ZN(G1329gat));
  NOR2_X1   g552(.A1(new_n615_), .A2(new_n600_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n723_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n727_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n730_), .B(new_n754_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n600_), .B1(new_n707_), .B2(new_n666_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1330gat));
  AOI21_X1  g561(.A(G50gat), .B1(new_n708_), .B2(new_n702_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n702_), .A2(G50gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n731_), .B2(new_n764_), .ZN(G1331gat));
  NAND2_X1  g564(.A1(new_n378_), .A2(new_n380_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n382_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n378_), .A2(new_n380_), .A3(KEYINPUT83), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n674_), .ZN(new_n769_));
  NOR4_X1   g568(.A1(new_n667_), .A2(new_n285_), .A3(new_n672_), .A4(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n640_), .ZN(new_n771_));
  NOR4_X1   g570(.A1(new_n385_), .A2(new_n667_), .A3(new_n285_), .A4(new_n320_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n677_), .A2(G57gat), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n771_), .A2(G57gat), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n774_), .B(KEYINPUT110), .Z(G1332gat));
  INV_X1    g574(.A(G64gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n770_), .B2(new_n683_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT48), .Z(new_n778_));
  NAND3_X1  g577(.A1(new_n772_), .A2(new_n776_), .A3(new_n683_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1333gat));
  INV_X1    g579(.A(G71gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n770_), .B2(new_n665_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n772_), .A2(new_n781_), .A3(new_n665_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(G1334gat));
  INV_X1    g585(.A(G78gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n770_), .B2(new_n702_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT50), .Z(new_n789_));
  NAND3_X1  g588(.A1(new_n772_), .A2(new_n787_), .A3(new_n702_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1335gat));
  INV_X1    g590(.A(new_n285_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(new_n710_), .A3(new_n674_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n726_), .A2(new_n720_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT112), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n726_), .A2(new_n796_), .A3(new_n720_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n793_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n231_), .B1(new_n798_), .B2(new_n640_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n667_), .A2(new_n285_), .A3(new_n320_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n706_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n802_), .A2(G85gat), .A3(new_n677_), .ZN(new_n803_));
  OR3_X1    g602(.A1(new_n799_), .A2(new_n800_), .A3(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n799_), .B2(new_n803_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1336gat));
  INV_X1    g605(.A(new_n802_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G92gat), .B1(new_n807_), .B2(new_n683_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n682_), .A2(new_n230_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n798_), .B2(new_n809_), .ZN(G1337gat));
  AOI21_X1  g609(.A(new_n204_), .B1(new_n798_), .B2(new_n665_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n802_), .A2(new_n227_), .A3(new_n615_), .ZN(new_n812_));
  OR3_X1    g611(.A1(new_n811_), .A2(KEYINPUT51), .A3(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT51), .B1(new_n811_), .B2(new_n812_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1338gat));
  NOR2_X1   g614(.A1(new_n793_), .A2(new_n482_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n205_), .B1(new_n816_), .B2(new_n794_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n817_), .A2(KEYINPUT52), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n702_), .A2(new_n205_), .ZN(new_n819_));
  OR3_X1    g618(.A1(new_n802_), .A2(KEYINPUT114), .A3(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT114), .B1(new_n802_), .B2(new_n819_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n817_), .A2(KEYINPUT52), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n818_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT53), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n818_), .A2(new_n822_), .A3(new_n826_), .A4(new_n823_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1339gat));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n769_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n384_), .A2(KEYINPUT115), .A3(new_n674_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n283_), .A2(new_n277_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n832_), .A2(new_n362_), .A3(new_n833_), .A4(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n834_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n830_), .A2(new_n833_), .A3(new_n831_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n717_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n835_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(KEYINPUT58), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n247_), .B(new_n260_), .C1(new_n256_), .C2(new_n258_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n250_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n259_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n255_), .B1(new_n251_), .B2(new_n245_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n257_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n254_), .A2(KEYINPUT70), .A3(new_n255_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n849_), .A2(KEYINPUT55), .A3(new_n247_), .A4(new_n252_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n843_), .A2(new_n845_), .A3(new_n850_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n851_), .A2(KEYINPUT56), .A3(new_n268_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT56), .B1(new_n851_), .B2(new_n268_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n852_), .A2(new_n853_), .A3(KEYINPUT118), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n268_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(KEYINPUT118), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n311_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n309_), .B1(new_n858_), .B2(new_n306_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(KEYINPUT117), .A3(new_n317_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n859_), .B2(new_n316_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n305_), .A2(new_n306_), .A3(new_n309_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n865_), .A2(new_n319_), .A3(new_n270_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n857_), .A2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n841_), .B1(new_n854_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n855_), .A2(new_n856_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n851_), .A2(KEYINPUT56), .A3(new_n268_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n841_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n872_), .A2(new_n873_), .A3(new_n857_), .A4(new_n866_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n868_), .A2(new_n717_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n320_), .A2(new_n270_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n877_));
  AND4_X1   g676(.A1(new_n319_), .A2(new_n273_), .A3(new_n276_), .A4(new_n865_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n360_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n360_), .B(KEYINPUT57), .C1(new_n877_), .C2(new_n878_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n875_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n710_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n839_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n683_), .A2(new_n702_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n677_), .A2(new_n615_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n885_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT59), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n883_), .A2(KEYINPUT121), .A3(new_n710_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT121), .B1(new_n883_), .B2(new_n710_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n839_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n888_), .A2(KEYINPUT59), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n320_), .B(new_n891_), .C1(new_n895_), .C2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G113gat), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n890_), .A2(KEYINPUT120), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n890_), .A2(KEYINPUT120), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n674_), .A2(G113gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n899_), .A2(new_n903_), .ZN(G1340gat));
  OAI211_X1 g703(.A(new_n792_), .B(new_n891_), .C1(new_n895_), .C2(new_n897_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(G120gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n285_), .A2(KEYINPUT60), .ZN(new_n907_));
  MUX2_X1   g706(.A(new_n907_), .B(KEYINPUT60), .S(G120gat), .Z(new_n908_));
  NAND3_X1  g707(.A1(new_n900_), .A2(new_n901_), .A3(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n906_), .A2(new_n909_), .ZN(G1341gat));
  NAND3_X1  g709(.A1(new_n900_), .A2(new_n901_), .A3(new_n384_), .ZN(new_n911_));
  INV_X1    g710(.A(G127gat), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n894_), .A2(new_n896_), .B1(new_n890_), .B2(KEYINPUT59), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n384_), .A2(G127gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT122), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n911_), .A2(new_n912_), .B1(new_n913_), .B2(new_n915_), .ZN(G1342gat));
  OAI211_X1 g715(.A(new_n717_), .B(new_n891_), .C1(new_n895_), .C2(new_n897_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(G134gat), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n360_), .A2(G134gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n900_), .A2(new_n901_), .A3(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(G1343gat));
  NAND2_X1  g720(.A1(new_n835_), .A2(new_n838_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n710_), .B2(new_n883_), .ZN(new_n923_));
  NOR4_X1   g722(.A1(new_n683_), .A2(new_n665_), .A3(new_n677_), .A4(new_n482_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(KEYINPUT123), .B1(new_n923_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n885_), .A2(new_n927_), .A3(new_n924_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT124), .B(G141gat), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n929_), .A2(new_n320_), .A3(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n929_), .B2(new_n320_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1344gat));
  XNOR2_X1  g732(.A(KEYINPUT125), .B(G148gat), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n929_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n936_), .B2(new_n285_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n929_), .A2(new_n792_), .A3(new_n934_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1345gat));
  XNOR2_X1  g738(.A(KEYINPUT61), .B(G155gat), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n940_), .B1(new_n936_), .B2(new_n710_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n940_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n929_), .A2(new_n384_), .A3(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1346gat));
  OAI21_X1  g743(.A(G162gat), .B1(new_n936_), .B2(new_n362_), .ZN(new_n945_));
  INV_X1    g744(.A(G162gat), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n929_), .A2(new_n946_), .A3(new_n672_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n947_), .ZN(G1347gat));
  NOR3_X1   g747(.A1(new_n666_), .A2(new_n640_), .A3(new_n682_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n894_), .A2(new_n482_), .A3(new_n320_), .A4(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(G169gat), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  AND2_X1   g752(.A1(new_n894_), .A2(new_n482_), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n954_), .A2(new_n516_), .A3(new_n320_), .A4(new_n949_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n950_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n953_), .A2(new_n955_), .A3(new_n956_), .ZN(G1348gat));
  NAND2_X1  g756(.A1(new_n885_), .A2(new_n482_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n949_), .ZN(new_n959_));
  NOR4_X1   g758(.A1(new_n958_), .A2(new_n517_), .A3(new_n285_), .A4(new_n959_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n954_), .A2(new_n792_), .A3(new_n949_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n960_), .B1(new_n961_), .B2(new_n517_), .ZN(G1349gat));
  NAND2_X1  g761(.A1(new_n949_), .A2(new_n384_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n963_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n954_), .A2(KEYINPUT126), .A3(new_n964_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n494_), .B1(new_n958_), .B2(new_n963_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n894_), .A2(new_n482_), .A3(new_n964_), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(new_n968_), .ZN(new_n969_));
  AND3_X1   g768(.A1(new_n965_), .A2(new_n966_), .A3(new_n969_), .ZN(G1350gat));
  NAND4_X1  g769(.A1(new_n954_), .A2(new_n672_), .A3(new_n532_), .A4(new_n949_), .ZN(new_n971_));
  NOR4_X1   g770(.A1(new_n895_), .A2(new_n362_), .A3(new_n702_), .A4(new_n959_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n972_), .B2(new_n488_), .ZN(G1351gat));
  NOR3_X1   g772(.A1(new_n665_), .A2(new_n640_), .A3(new_n482_), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n885_), .A2(new_n683_), .A3(new_n974_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n975_), .A2(new_n674_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(new_n391_), .ZN(G1352gat));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n975_), .A2(new_n285_), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n978_), .B1(new_n979_), .B2(new_n387_), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n979_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n981_));
  OAI211_X1 g780(.A(KEYINPUT127), .B(G204gat), .C1(new_n975_), .C2(new_n285_), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n980_), .A2(new_n981_), .A3(new_n982_), .ZN(G1353gat));
  NOR2_X1   g782(.A1(new_n975_), .A2(new_n710_), .ZN(new_n984_));
  NOR3_X1   g783(.A1(new_n984_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n985_));
  XOR2_X1   g784(.A(KEYINPUT63), .B(G211gat), .Z(new_n986_));
  AOI21_X1  g785(.A(new_n985_), .B1(new_n984_), .B2(new_n986_), .ZN(G1354gat));
  OAI21_X1  g786(.A(G218gat), .B1(new_n975_), .B2(new_n362_), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n672_), .A2(new_n396_), .ZN(new_n989_));
  OAI21_X1  g788(.A(new_n988_), .B1(new_n975_), .B2(new_n989_), .ZN(G1355gat));
endmodule


