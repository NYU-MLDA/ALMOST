//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n931_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n953_;
  NOR2_X1   g000(.A1(G197gat), .A2(G204gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT94), .B(G197gat), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n202_), .B1(new_n203_), .B2(G204gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G211gat), .B(G218gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(KEYINPUT21), .A3(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n204_), .A2(KEYINPUT21), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT21), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n209_), .B1(G197gat), .B2(G204gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(new_n203_), .B2(G204gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(new_n205_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n207_), .B1(new_n208_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  XOR2_X1   g016(.A(new_n217_), .B(KEYINPUT3), .Z(new_n218_));
  NAND2_X1  g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  XOR2_X1   g018(.A(new_n219_), .B(KEYINPUT2), .Z(new_n220_));
  OAI211_X1 g019(.A(new_n215_), .B(new_n216_), .C1(new_n218_), .C2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n217_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT93), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(new_n215_), .B2(KEYINPUT1), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n215_), .A2(KEYINPUT1), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n216_), .ZN(new_n226_));
  NOR3_X1   g025(.A1(new_n215_), .A2(new_n223_), .A3(KEYINPUT1), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n222_), .B(new_n219_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n221_), .A2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n214_), .B1(KEYINPUT29), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G228gat), .A2(G233gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n232_), .A2(KEYINPUT95), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G78gat), .B(G106gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n229_), .A2(KEYINPUT29), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G22gat), .B(G50gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT28), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n237_), .B(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n234_), .B1(new_n232_), .B2(KEYINPUT95), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n236_), .B(new_n240_), .C1(new_n233_), .C2(new_n241_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n234_), .A2(KEYINPUT96), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n240_), .B1(new_n232_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n244_), .B1(new_n232_), .B2(new_n243_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G71gat), .B(G99gat), .ZN(new_n247_));
  INV_X1    g046(.A(G169gat), .ZN(new_n248_));
  INV_X1    g047(.A(G176gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT22), .B1(new_n248_), .B2(KEYINPUT87), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT87), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT22), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(G169gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n254_), .A3(new_n249_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n250_), .B1(new_n255_), .B2(KEYINPUT88), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n256_), .B1(KEYINPUT88), .B2(new_n255_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT89), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT23), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(G183gat), .B2(G190gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n258_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n261_), .B(new_n266_), .C1(new_n250_), .C2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G190gat), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n271_), .A2(KEYINPUT86), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT25), .B(G183gat), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT26), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(G190gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(KEYINPUT86), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n269_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n264_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT90), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT90), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n264_), .A2(new_n280_), .A3(new_n277_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n279_), .A2(KEYINPUT30), .A3(new_n281_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G15gat), .B(G43gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n286_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n247_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G127gat), .B(G134gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT92), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G113gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G120gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n293_), .B(G113gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(G120gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT31), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT91), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G227gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n284_), .A2(new_n285_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n286_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n247_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(new_n308_), .A3(new_n287_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n290_), .A2(new_n304_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n304_), .B1(new_n290_), .B2(new_n309_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n246_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n304_), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n288_), .A2(new_n289_), .A3(new_n247_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n308_), .B1(new_n307_), .B2(new_n287_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n290_), .A2(new_n304_), .A3(new_n309_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n246_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G226gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT19), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n279_), .A2(new_n281_), .A3(new_n214_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT20), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT22), .B(G169gat), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n250_), .B1(new_n326_), .B2(new_n249_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n262_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n273_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(new_n271_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n268_), .B2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n325_), .B1(new_n331_), .B2(new_n213_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n323_), .B1(new_n324_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n282_), .A2(new_n213_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT20), .B1(new_n331_), .B2(new_n213_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n323_), .A3(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G8gat), .B(G36gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT18), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(G64gat), .ZN(new_n341_));
  INV_X1    g140(.A(G92gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n334_), .A2(new_n338_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT27), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n214_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n322_), .B1(new_n346_), .B2(new_n336_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n324_), .A2(new_n323_), .A3(new_n332_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n343_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT103), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(KEYINPUT103), .A3(new_n350_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n345_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n229_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n298_), .A2(G120gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n295_), .A2(new_n296_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n229_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(KEYINPUT4), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT98), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n364_), .B(new_n229_), .C1(new_n297_), .C2(new_n299_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n356_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G1gat), .B(G29gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G57gat), .B(G85gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n373_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n366_), .A2(new_n367_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n346_), .A2(new_n322_), .A3(new_n336_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n350_), .B1(new_n378_), .B2(new_n333_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT27), .B1(new_n344_), .B2(new_n379_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n355_), .A2(new_n377_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n320_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n343_), .A2(KEYINPUT32), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n334_), .A2(new_n338_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT101), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT102), .ZN(new_n387_));
  INV_X1    g186(.A(new_n383_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n349_), .B2(new_n388_), .ZN(new_n389_));
  AOI211_X1 g188(.A(KEYINPUT102), .B(new_n383_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n377_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT33), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n376_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n361_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n356_), .A2(new_n360_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT100), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n363_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n395_), .A2(new_n396_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n373_), .B(new_n394_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n366_), .A2(KEYINPUT33), .A3(new_n367_), .A4(new_n375_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n393_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT97), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n344_), .A2(new_n379_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n344_), .B2(new_n379_), .ZN(new_n406_));
  OAI22_X1  g205(.A1(new_n386_), .A2(new_n391_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n246_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n382_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT85), .ZN(new_n411_));
  INV_X1    g210(.A(G36gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(G29gat), .ZN(new_n413_));
  INV_X1    g212(.A(G29gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(G36gat), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n413_), .A2(new_n415_), .A3(KEYINPUT71), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT71), .B1(new_n413_), .B2(new_n415_), .ZN(new_n417_));
  OAI21_X1  g216(.A(G43gat), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT71), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n414_), .A2(G36gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n412_), .A2(G29gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(G43gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n413_), .A2(new_n415_), .A3(KEYINPUT71), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n418_), .A2(G50gat), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(G50gat), .B1(new_n418_), .B2(new_n425_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT72), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G50gat), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n416_), .A2(new_n417_), .A3(G43gat), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n423_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT72), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n418_), .A2(new_n425_), .A3(G50gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n428_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT15), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(KEYINPUT76), .B(G1gat), .Z(new_n439_));
  INV_X1    g238(.A(G8gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT14), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G15gat), .B(G22gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G1gat), .B(G8gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT77), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n443_), .B(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n428_), .A2(KEYINPUT15), .A3(new_n435_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n438_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G229gat), .A2(G233gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT80), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n432_), .A2(KEYINPUT80), .A3(new_n434_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n445_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(new_n443_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n450_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n448_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n426_), .A2(new_n427_), .A3(new_n451_), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT80), .B1(new_n432_), .B2(new_n434_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n456_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n452_), .A2(new_n446_), .A3(new_n453_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(KEYINPUT81), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT81), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n452_), .A2(new_n446_), .A3(new_n465_), .A4(new_n453_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n450_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n464_), .A2(KEYINPUT82), .A3(new_n450_), .A4(new_n466_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n459_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G113gat), .B(G141gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT84), .B(G197gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT83), .B(G169gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n411_), .B1(new_n471_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n469_), .A2(new_n470_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n458_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n476_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n411_), .A3(new_n476_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT8), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NOR3_X1   g287(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(KEYINPUT65), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT65), .ZN(new_n496_));
  AND3_X1   g295(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n490_), .A2(new_n495_), .A3(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G85gat), .B(G92gat), .Z(new_n501_));
  AOI21_X1  g300(.A(new_n486_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT66), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT66), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n497_), .A2(new_n498_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n490_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(new_n486_), .A3(new_n501_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n504_), .A2(new_n506_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT67), .ZN(new_n511_));
  XOR2_X1   g310(.A(G71gat), .B(G78gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(G57gat), .B(G64gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n512_), .B1(KEYINPUT11), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(KEYINPUT11), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT9), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT64), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n518_), .A2(KEYINPUT64), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n501_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT10), .B(G99gat), .Z(new_n522_));
  INV_X1    g321(.A(G106gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n518_), .A2(KEYINPUT64), .A3(G85gat), .A4(G92gat), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n521_), .A2(new_n524_), .A3(new_n525_), .A4(new_n507_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n510_), .A2(new_n511_), .A3(new_n517_), .A4(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n509_), .B1(new_n502_), .B2(new_n505_), .ZN(new_n528_));
  AOI211_X1 g327(.A(KEYINPUT66), .B(new_n486_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n517_), .B(new_n526_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT67), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n526_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n516_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n527_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G230gat), .A2(G233gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n530_), .A2(new_n535_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n533_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT68), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(KEYINPUT12), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n532_), .A2(new_n516_), .A3(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n539_), .A2(new_n542_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n537_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G120gat), .B(G148gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT70), .ZN(new_n550_));
  XOR2_X1   g349(.A(G176gat), .B(G204gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n548_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n537_), .A2(new_n547_), .A3(new_n554_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT13), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n485_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT73), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(G134gat), .ZN(new_n564_));
  INV_X1    g363(.A(G162gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT36), .Z(new_n567_));
  INV_X1    g366(.A(new_n532_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n426_), .A2(new_n427_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT34), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n568_), .A2(new_n569_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n438_), .A2(new_n532_), .A3(new_n447_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n573_), .A2(new_n570_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n577_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n574_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n567_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n574_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n579_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n585_));
  AND2_X1   g384(.A1(new_n566_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(KEYINPUT75), .A3(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n578_), .A2(new_n580_), .A3(new_n586_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT75), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n581_), .B1(new_n587_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT37), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AOI211_X1 g392(.A(KEYINPUT37), .B(new_n581_), .C1(new_n587_), .C2(new_n590_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n456_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(new_n516_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT78), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n597_), .B(new_n517_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT78), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G127gat), .B(G155gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT16), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(G183gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(G211gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT17), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n599_), .A2(new_n602_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT79), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT17), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n606_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n600_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n595_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n410_), .A2(new_n561_), .A3(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT104), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(new_n377_), .A3(new_n439_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT38), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n616_), .A2(new_n591_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n410_), .A2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT105), .B1(new_n623_), .B2(new_n560_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT105), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n410_), .A2(new_n625_), .A3(new_n561_), .A4(new_n622_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n377_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(G1gat), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n621_), .A2(new_n628_), .ZN(G1324gat));
  NOR2_X1   g428(.A1(new_n355_), .A2(new_n380_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n619_), .A2(new_n440_), .A3(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n410_), .A2(new_n561_), .A3(new_n631_), .A4(new_n622_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n633_), .A2(new_n634_), .A3(G8gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n633_), .B2(G8gat), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n632_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(G1325gat));
  NOR2_X1   g438(.A1(new_n310_), .A2(new_n311_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n624_), .A2(new_n640_), .A3(new_n626_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G15gat), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT106), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n641_), .A2(new_n644_), .A3(G15gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT41), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(G15gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n619_), .A2(new_n649_), .A3(new_n640_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n643_), .A2(KEYINPUT41), .A3(new_n645_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n650_), .A3(new_n651_), .ZN(G1326gat));
  INV_X1    g451(.A(G22gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n619_), .A2(new_n653_), .A3(new_n246_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n624_), .A2(new_n246_), .A3(new_n626_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n655_), .A2(new_n656_), .A3(G22gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n655_), .B2(G22gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(G1327gat));
  AOI22_X1  g458(.A1(new_n610_), .A2(new_n611_), .B1(new_n614_), .B2(new_n600_), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT75), .B1(new_n584_), .B2(new_n586_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n588_), .A2(new_n589_), .ZN(new_n662_));
  OAI22_X1  g461(.A1(new_n661_), .A2(new_n662_), .B1(new_n584_), .B2(new_n567_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n660_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n410_), .A2(new_n561_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G29gat), .B1(new_n666_), .B2(new_n377_), .ZN(new_n667_));
  AOI22_X1  g466(.A1(new_n320_), .A2(new_n381_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n663_), .A2(KEYINPUT37), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n591_), .A2(new_n592_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(KEYINPUT43), .B1(new_n668_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n353_), .A2(new_n354_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n345_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n377_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n380_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n676_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n312_), .B2(new_n319_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n407_), .A2(new_n408_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n673_), .B(new_n595_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n672_), .A2(new_n682_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n683_), .A2(KEYINPUT44), .A3(new_n561_), .A4(new_n616_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n684_), .A2(G29gat), .A3(new_n377_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n683_), .A2(new_n561_), .A3(new_n616_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n667_), .B1(new_n685_), .B2(new_n688_), .ZN(G1328gat));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  AOI211_X1 g489(.A(new_n560_), .B(new_n660_), .C1(new_n672_), .C2(new_n682_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n630_), .B1(new_n691_), .B2(KEYINPUT44), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n412_), .B1(new_n692_), .B2(new_n688_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT45), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n630_), .A2(G36gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT107), .B1(new_n665_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n665_), .A2(KEYINPUT107), .A3(new_n696_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n699_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(KEYINPUT45), .A3(new_n697_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n690_), .B1(new_n693_), .B2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n691_), .A2(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n684_), .A2(new_n631_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G36gat), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n707_), .A2(KEYINPUT46), .A3(new_n702_), .A4(new_n700_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n704_), .A2(new_n708_), .ZN(G1329gat));
  INV_X1    g508(.A(new_n640_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n423_), .B1(new_n665_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT108), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n684_), .A2(G43gat), .A3(new_n640_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n705_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n712_), .B(new_n715_), .C1(new_n713_), .C2(new_n705_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1330gat));
  NAND3_X1  g518(.A1(new_n666_), .A2(new_n429_), .A3(new_n246_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n684_), .A2(new_n246_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n705_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G50gat), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n705_), .A2(new_n722_), .A3(new_n721_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n720_), .B1(new_n724_), .B2(new_n725_), .ZN(G1331gat));
  NOR2_X1   g525(.A1(new_n485_), .A2(new_n559_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n671_), .A2(new_n660_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n410_), .A2(new_n730_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(KEYINPUT111), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(KEYINPUT111), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n377_), .A3(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(G57gat), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n623_), .A2(new_n728_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n677_), .A2(new_n735_), .ZN(new_n737_));
  AOI22_X1  g536(.A1(new_n734_), .A2(new_n735_), .B1(new_n736_), .B2(new_n737_), .ZN(G1332gat));
  INV_X1    g537(.A(G64gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n736_), .B2(new_n631_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT48), .Z(new_n741_));
  INV_X1    g540(.A(new_n731_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(new_n739_), .A3(new_n631_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n736_), .B2(new_n640_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT49), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n742_), .A2(new_n745_), .A3(new_n640_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1334gat));
  INV_X1    g548(.A(G78gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n736_), .B2(new_n246_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT50), .Z(new_n752_));
  NAND2_X1  g551(.A1(new_n246_), .A2(new_n750_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT112), .Z(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n731_), .B2(new_n754_), .ZN(G1335gat));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n683_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n672_), .A2(KEYINPUT113), .A3(new_n682_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n728_), .A2(new_n660_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n677_), .ZN(new_n761_));
  NOR4_X1   g560(.A1(new_n668_), .A2(new_n663_), .A3(new_n660_), .A4(new_n728_), .ZN(new_n762_));
  INV_X1    g561(.A(G85gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(new_n377_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(new_n764_), .ZN(G1336gat));
  OAI21_X1  g564(.A(G92gat), .B1(new_n760_), .B2(new_n630_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(new_n342_), .A3(new_n631_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT114), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n766_), .A2(new_n770_), .A3(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n760_), .B2(new_n710_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n762_), .A2(new_n522_), .A3(new_n640_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT51), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n773_), .A2(new_n777_), .A3(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1338gat));
  NAND3_X1  g578(.A1(new_n762_), .A2(new_n523_), .A3(new_n246_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n683_), .A2(new_n246_), .A3(new_n616_), .A4(new_n727_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n781_), .A2(new_n782_), .A3(G106gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n781_), .B2(G106gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT53), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n787_), .B(new_n780_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1339gat));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n484_), .A2(new_n559_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n790_), .B1(new_n617_), .B2(new_n792_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n729_), .A2(KEYINPUT54), .A3(new_n791_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n449_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n448_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n464_), .A2(new_n449_), .A3(new_n466_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n476_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n799_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(KEYINPUT116), .A3(new_n476_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n471_), .A2(new_n477_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT117), .B1(new_n805_), .B2(new_n558_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n471_), .A2(new_n477_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n801_), .A2(new_n802_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n799_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n804_), .A3(new_n809_), .ZN(new_n810_));
  AND4_X1   g609(.A1(KEYINPUT117), .A2(new_n807_), .A3(new_n558_), .A4(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n806_), .A2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n539_), .A2(new_n542_), .A3(KEYINPUT55), .A4(new_n546_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n532_), .A2(new_n516_), .A3(new_n545_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n540_), .B1(new_n532_), .B2(new_n516_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n538_), .ZN(new_n816_));
  XOR2_X1   g615(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n817_));
  OAI21_X1  g616(.A(new_n813_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n527_), .A2(new_n531_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n814_), .A2(new_n815_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n535_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n555_), .B1(new_n818_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n542_), .A2(new_n546_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n527_), .A2(new_n531_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n536_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n817_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n547_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n827_), .A2(new_n829_), .A3(new_n813_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n555_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n824_), .A2(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n832_), .A2(new_n482_), .A3(new_n557_), .A4(new_n483_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n591_), .B1(new_n812_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n797_), .B1(new_n834_), .B2(KEYINPUT118), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836_));
  AOI211_X1 g635(.A(new_n836_), .B(new_n591_), .C1(new_n812_), .C2(new_n833_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n796_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n833_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n807_), .A2(new_n558_), .A3(new_n810_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n805_), .A2(KEYINPUT117), .A3(new_n558_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n663_), .B1(new_n839_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n836_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n834_), .A2(KEYINPUT118), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(KEYINPUT119), .A4(new_n797_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n807_), .A2(new_n557_), .A3(new_n810_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n832_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n849_), .A2(new_n832_), .A3(KEYINPUT58), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n595_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n595_), .A2(new_n852_), .A3(KEYINPUT121), .A4(new_n853_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n856_), .A2(new_n857_), .B1(KEYINPUT57), .B2(new_n834_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n838_), .A2(new_n848_), .A3(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n795_), .B1(new_n859_), .B2(new_n616_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n630_), .A2(new_n377_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n319_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT59), .B1(new_n860_), .B2(new_n863_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n853_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n834_), .A2(KEYINPUT57), .B1(new_n865_), .B2(new_n852_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n795_), .B1(new_n867_), .B2(new_n616_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n863_), .A2(KEYINPUT59), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT123), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n846_), .A2(new_n797_), .A3(new_n847_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n660_), .B1(new_n873_), .B2(new_n866_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n869_), .B(new_n872_), .C1(new_n874_), .C2(new_n795_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n484_), .A2(new_n294_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n864_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n860_), .A2(new_n484_), .A3(new_n863_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(G113gat), .ZN(new_n881_));
  INV_X1    g680(.A(new_n860_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(new_n485_), .A3(new_n862_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(KEYINPUT122), .A3(new_n294_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n878_), .B1(new_n881_), .B2(new_n884_), .ZN(G1340gat));
  INV_X1    g684(.A(new_n559_), .ZN(new_n886_));
  AOI21_X1  g685(.A(KEYINPUT60), .B1(new_n886_), .B2(new_n296_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(KEYINPUT60), .B2(new_n296_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n882_), .A2(new_n862_), .A3(new_n888_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n864_), .A2(new_n876_), .A3(new_n886_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n296_), .ZN(G1341gat));
  NAND3_X1  g690(.A1(new_n864_), .A2(new_n876_), .A3(new_n660_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G127gat), .ZN(new_n893_));
  OR4_X1    g692(.A1(G127gat), .A2(new_n860_), .A3(new_n616_), .A4(new_n863_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1342gat));
  NAND3_X1  g694(.A1(new_n864_), .A2(new_n876_), .A3(new_n595_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(G134gat), .ZN(new_n897_));
  OR4_X1    g696(.A1(G134gat), .A2(new_n860_), .A3(new_n663_), .A4(new_n863_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1343gat));
  NOR2_X1   g698(.A1(new_n861_), .A2(new_n312_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n860_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n485_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n886_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT124), .B(G148gat), .Z(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1345gat));
  NAND2_X1  g706(.A1(new_n902_), .A2(new_n660_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G155gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT126), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n908_), .B(new_n911_), .ZN(G1346gat));
  NAND3_X1  g711(.A1(new_n902_), .A2(new_n565_), .A3(new_n591_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n860_), .A2(new_n671_), .A3(new_n901_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n565_), .B2(new_n914_), .ZN(G1347gat));
  NAND2_X1  g714(.A1(new_n631_), .A2(new_n677_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n710_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n318_), .ZN(new_n918_));
  OR3_X1    g717(.A1(new_n868_), .A2(KEYINPUT127), .A3(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT127), .B1(new_n868_), .B2(new_n918_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n919_), .A2(new_n485_), .A3(new_n326_), .A4(new_n920_), .ZN(new_n921_));
  OR3_X1    g720(.A1(new_n868_), .A2(new_n484_), .A3(new_n918_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n922_), .A2(new_n923_), .A3(G169gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n922_), .B2(G169gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n921_), .B1(new_n924_), .B2(new_n925_), .ZN(G1348gat));
  NAND3_X1  g725(.A1(new_n919_), .A2(new_n886_), .A3(new_n920_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n860_), .A2(new_n246_), .ZN(new_n928_));
  NOR4_X1   g727(.A1(new_n916_), .A2(new_n710_), .A3(new_n249_), .A4(new_n559_), .ZN(new_n929_));
  AOI22_X1  g728(.A1(new_n927_), .A2(new_n249_), .B1(new_n928_), .B2(new_n929_), .ZN(G1349gat));
  AND4_X1   g729(.A1(new_n329_), .A2(new_n919_), .A3(new_n660_), .A4(new_n920_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n916_), .A2(new_n710_), .A3(new_n616_), .ZN(new_n932_));
  AOI21_X1  g731(.A(G183gat), .B1(new_n928_), .B2(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n931_), .A2(new_n933_), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n919_), .A2(new_n595_), .A3(new_n920_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(G190gat), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n919_), .A2(new_n270_), .A3(new_n591_), .A4(new_n920_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1351gat));
  NOR2_X1   g737(.A1(new_n916_), .A2(new_n312_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n860_), .A2(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n485_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n886_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  NAND2_X1  g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  AND4_X1   g746(.A1(new_n660_), .A2(new_n941_), .A3(new_n946_), .A4(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n946_), .B1(new_n941_), .B2(new_n660_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n948_), .A2(new_n949_), .ZN(G1354gat));
  INV_X1    g749(.A(G218gat), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n941_), .A2(new_n951_), .A3(new_n591_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n860_), .A2(new_n671_), .A3(new_n940_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n951_), .B2(new_n953_), .ZN(G1355gat));
endmodule


