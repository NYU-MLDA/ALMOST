//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203_));
  INV_X1    g002(.A(G71gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G99gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G15gat), .B(G43gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n207_), .B(new_n210_), .Z(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT23), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n216_), .A3(KEYINPUT82), .ZN(new_n217_));
  INV_X1    g016(.A(G183gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT80), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G183gat), .ZN(new_n221_));
  INV_X1    g020(.A(G190gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n219_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT82), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n213_), .A2(new_n224_), .A3(KEYINPUT23), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n217_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT81), .ZN(new_n227_));
  INV_X1    g026(.A(G169gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT22), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G169gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n227_), .B1(new_n232_), .B2(G176gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G169gat), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n235_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n226_), .B(new_n233_), .C1(new_n227_), .C2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT83), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n222_), .A2(KEYINPUT26), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G190gat), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n245_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n244_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n228_), .A2(new_n237_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(KEYINPUT24), .A3(new_n234_), .ZN(new_n250_));
  OR3_X1    g049(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n214_), .A2(new_n216_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n248_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n239_), .A2(new_n240_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n240_), .B1(new_n239_), .B2(new_n254_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT30), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n239_), .A2(new_n254_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT83), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n239_), .A2(new_n254_), .A3(new_n240_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n258_), .A2(new_n264_), .A3(KEYINPUT86), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT86), .B1(new_n258_), .B2(new_n264_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n212_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n212_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G127gat), .B(G134gat), .Z(new_n271_));
  XOR2_X1   g070(.A(G113gat), .B(G120gat), .Z(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT87), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G127gat), .B(G134gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G113gat), .B(G120gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n276_), .A3(KEYINPUT87), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT31), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n268_), .A2(new_n270_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n281_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT86), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n257_), .A2(KEYINPUT30), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n262_), .A2(new_n263_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n284_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n211_), .B1(new_n287_), .B2(new_n265_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n283_), .B1(new_n288_), .B2(new_n269_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n282_), .A2(new_n289_), .ZN(new_n290_));
  OR3_X1    g089(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n291_), .A2(new_n294_), .A3(new_n295_), .A4(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(G155gat), .ZN(new_n298_));
  INV_X1    g097(.A(G162gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n299_), .A3(KEYINPUT88), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT88), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(G155gat), .B2(G162gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT89), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT89), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(G155gat), .A3(G162gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n297_), .A2(new_n304_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n306_), .A2(new_n308_), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n303_), .ZN(new_n314_));
  INV_X1    g113(.A(G141gat), .ZN(new_n315_));
  INV_X1    g114(.A(G148gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n292_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n310_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n319_), .A2(KEYINPUT29), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n322_));
  OR2_X1    g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n322_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G228gat), .A2(G233gat), .ZN(new_n326_));
  INV_X1    g125(.A(G78gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(G106gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n323_), .A2(new_n332_), .A3(new_n324_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G197gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G204gat), .ZN(new_n336_));
  INV_X1    g135(.A(G204gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G197gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n339_), .A2(KEYINPUT21), .ZN(new_n340_));
  XOR2_X1   g139(.A(G211gat), .B(G218gat), .Z(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n335_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n343_));
  OAI211_X1 g142(.A(KEYINPUT21), .B(new_n343_), .C1(new_n339_), .C2(KEYINPUT91), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT92), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n339_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n336_), .A2(new_n338_), .A3(KEYINPUT92), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n347_), .A2(KEYINPUT21), .A3(new_n341_), .A4(new_n348_), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n350_), .B1(new_n319_), .B2(KEYINPUT29), .ZN(new_n351_));
  XOR2_X1   g150(.A(G22gat), .B(G50gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n334_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n331_), .A2(new_n353_), .A3(new_n333_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n290_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT27), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT18), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G64gat), .B(G92gat), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  NAND2_X1  g162(.A1(G226gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT19), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n345_), .A2(new_n349_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n255_), .A2(new_n256_), .A3(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n241_), .B(new_n243_), .C1(new_n368_), .C2(new_n247_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n369_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT93), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n217_), .A2(new_n225_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n369_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n217_), .A2(new_n225_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT93), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n232_), .A2(KEYINPUT94), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n232_), .A2(KEYINPUT94), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n237_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n218_), .A2(new_n222_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n235_), .B1(new_n253_), .B2(new_n380_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n373_), .A2(new_n376_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT20), .B1(new_n382_), .B2(new_n350_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n365_), .B1(new_n367_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT95), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT20), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n379_), .A2(new_n381_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n371_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(new_n374_), .A2(new_n375_), .A3(KEYINPUT93), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n386_), .B1(new_n390_), .B2(new_n366_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n260_), .A2(new_n261_), .A3(new_n350_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT95), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(new_n365_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n385_), .A2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n366_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n365_), .B1(new_n382_), .B2(new_n350_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n397_), .A2(new_n398_), .A3(KEYINPUT20), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n363_), .B1(new_n396_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n363_), .ZN(new_n402_));
  AOI211_X1 g201(.A(new_n399_), .B(new_n402_), .C1(new_n385_), .C2(new_n395_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n359_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n399_), .B1(new_n385_), .B2(new_n395_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n363_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n350_), .B(new_n387_), .C1(new_n375_), .C2(new_n374_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n397_), .A2(new_n407_), .A3(KEYINPUT20), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n365_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n365_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n391_), .A2(new_n392_), .A3(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n406_), .B(KEYINPUT27), .C1(new_n363_), .C2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n358_), .A2(new_n404_), .A3(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(G85gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT0), .B(G57gat), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n416_), .B(new_n417_), .Z(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n278_), .A2(new_n279_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n319_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n273_), .A2(new_n277_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n310_), .B(new_n422_), .C1(new_n314_), .C2(new_n318_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n421_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n309_), .A2(KEYINPUT1), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n306_), .A2(new_n308_), .A3(new_n311_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n304_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n318_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n303_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n429_), .A2(new_n430_), .B1(new_n431_), .B2(new_n297_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n423_), .B(KEYINPUT4), .C1(new_n280_), .C2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT96), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT96), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n421_), .A2(new_n435_), .A3(KEYINPUT4), .A4(new_n423_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n424_), .B(KEYINPUT97), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n421_), .B2(KEYINPUT4), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT98), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n426_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n439_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n444_), .A2(KEYINPUT98), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n419_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT100), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n441_), .A2(new_n442_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n425_), .B1(new_n444_), .B2(KEYINPUT98), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n418_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n451_));
  OAI211_X1 g250(.A(KEYINPUT100), .B(new_n419_), .C1(new_n443_), .C2(new_n445_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n202_), .B1(new_n414_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n413_), .A2(new_n404_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n457_), .A2(KEYINPUT102), .A3(new_n453_), .A4(new_n358_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT99), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n450_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT33), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n450_), .A2(new_n460_), .A3(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n401_), .A2(new_n403_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n437_), .B(new_n424_), .C1(KEYINPUT4), .C2(new_n421_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n421_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n423_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n418_), .B1(new_n469_), .B2(new_n438_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n462_), .A2(new_n464_), .A3(new_n465_), .A4(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n363_), .A2(KEYINPUT32), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n473_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n474_), .B1(new_n405_), .B2(new_n473_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n451_), .A2(new_n452_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n357_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT101), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n357_), .B1(new_n472_), .B2(new_n476_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT101), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n457_), .A2(new_n357_), .A3(new_n453_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n459_), .B1(new_n485_), .B2(new_n290_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT14), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT74), .B(G1gat), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n487_), .B1(new_n488_), .B2(G8gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT75), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G15gat), .B(G22gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G1gat), .B(G8gat), .Z(new_n494_));
  OR2_X1    g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n494_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G29gat), .B(G36gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G43gat), .B(G50gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n497_), .B(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G229gat), .A2(G233gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n497_), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT68), .B(KEYINPUT15), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n500_), .B(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n497_), .A2(new_n500_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(new_n502_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n504_), .A2(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G113gat), .B(G141gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT79), .ZN(new_n513_));
  XOR2_X1   g312(.A(G169gat), .B(G197gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n511_), .B(new_n515_), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n486_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT13), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G230gat), .A2(G233gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G85gat), .B(G92gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT9), .ZN(new_n524_));
  XOR2_X1   g323(.A(KEYINPUT10), .B(G99gat), .Z(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n329_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT6), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT64), .B(G92gat), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT9), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(G85gat), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n524_), .A2(new_n526_), .A3(new_n528_), .A4(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT8), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT65), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n528_), .A2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(G99gat), .A2(G106gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT7), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n528_), .A2(new_n534_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n533_), .B1(new_n539_), .B2(new_n523_), .ZN(new_n540_));
  AOI211_X1 g339(.A(KEYINPUT8), .B(new_n522_), .C1(new_n537_), .C2(new_n528_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n532_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G71gat), .B(G78gat), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(KEYINPUT11), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n546_), .A2(new_n544_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n545_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n542_), .A2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n549_), .B(new_n532_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(KEYINPUT12), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT12), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n542_), .A2(new_n554_), .A3(new_n550_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n521_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT66), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n551_), .A2(new_n552_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n521_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G120gat), .B(G148gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT5), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G176gat), .B(G204gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n558_), .A2(new_n560_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n519_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT13), .A3(new_n566_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(KEYINPUT67), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(KEYINPUT67), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT69), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n542_), .A2(new_n578_), .A3(new_n507_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n542_), .B2(new_n507_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT71), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n500_), .B(new_n532_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT34), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT70), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n587_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n581_), .A2(new_n588_), .A3(KEYINPUT35), .A4(new_n584_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(KEYINPUT36), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n594_));
  OAI221_X1 g393(.A(new_n587_), .B1(KEYINPUT71), .B2(new_n594_), .C1(new_n579_), .C2(new_n580_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(new_n593_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT72), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT72), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n589_), .A2(new_n598_), .A3(new_n593_), .A4(new_n595_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n589_), .A2(new_n595_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n592_), .B(KEYINPUT36), .Z(new_n601_));
  AOI22_X1  g400(.A1(new_n597_), .A2(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(KEYINPUT73), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(KEYINPUT73), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n602_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT78), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT76), .Z(new_n613_));
  OR2_X1    g412(.A1(new_n497_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n497_), .A2(new_n613_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n549_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(new_n550_), .A3(new_n615_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G127gat), .B(G155gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT16), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n621_), .B(new_n622_), .Z(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT17), .Z(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n611_), .B1(new_n619_), .B2(new_n625_), .ZN(new_n626_));
  AOI211_X1 g425(.A(KEYINPUT78), .B(new_n624_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n623_), .A2(new_n628_), .ZN(new_n629_));
  OAI22_X1  g428(.A1(new_n626_), .A2(new_n627_), .B1(new_n619_), .B2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n610_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n518_), .A2(new_n577_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT103), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT103), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n518_), .A2(new_n577_), .A3(new_n634_), .A4(new_n631_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n488_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n454_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT38), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n636_), .A2(KEYINPUT38), .A3(new_n454_), .A4(new_n637_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n486_), .A2(new_n602_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n572_), .A2(new_n517_), .A3(new_n630_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n453_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(new_n641_), .A3(new_n645_), .ZN(G1324gat));
  NOR2_X1   g445(.A1(new_n457_), .A2(G8gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n633_), .A2(new_n635_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n484_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n651_));
  AOI211_X1 g450(.A(KEYINPUT101), .B(new_n357_), .C1(new_n472_), .C2(new_n476_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n290_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n455_), .A2(new_n458_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n602_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n655_), .A2(new_n456_), .A3(new_n656_), .A4(new_n643_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n650_), .B1(new_n657_), .B2(G8gat), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n657_), .A2(new_n650_), .A3(G8gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n649_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n660_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n662_), .A2(new_n658_), .A3(KEYINPUT39), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n648_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n648_), .B(new_n665_), .C1(new_n661_), .C2(new_n663_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1325gat));
  OAI21_X1  g468(.A(G15gat), .B1(new_n644_), .B2(new_n290_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT41), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n632_), .A2(G15gat), .A3(new_n290_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1326gat));
  XNOR2_X1  g472(.A(new_n357_), .B(KEYINPUT106), .ZN(new_n674_));
  OAI21_X1  g473(.A(G22gat), .B1(new_n644_), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT42), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n674_), .A2(G22gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n632_), .B2(new_n677_), .ZN(G1327gat));
  INV_X1    g477(.A(new_n630_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n572_), .A2(new_n517_), .A3(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n655_), .B2(new_n610_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(KEYINPUT107), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n609_), .B(new_n684_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n685_));
  OAI211_X1 g484(.A(KEYINPUT44), .B(new_n680_), .C1(new_n682_), .C2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n680_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n681_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n688_), .B1(new_n486_), .B2(new_n609_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n684_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n655_), .A2(new_n610_), .A3(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n687_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n693_));
  OAI21_X1  g492(.A(new_n686_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694_), .B2(new_n453_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n656_), .A2(new_n679_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n572_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n655_), .A2(new_n516_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT109), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n655_), .A2(new_n701_), .A3(new_n516_), .A4(new_n698_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n453_), .A2(G29gat), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT110), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n695_), .A2(new_n706_), .ZN(G1328gat));
  OAI211_X1 g506(.A(new_n686_), .B(new_n456_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G36gat), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n457_), .A2(KEYINPUT111), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n457_), .A2(KEYINPUT111), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(G36gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n700_), .A2(new_n702_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT45), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n700_), .A2(new_n717_), .A3(new_n702_), .A4(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n709_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n709_), .A2(KEYINPUT46), .A3(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1329gat));
  INV_X1    g523(.A(new_n290_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n700_), .A2(new_n725_), .A3(new_n702_), .ZN(new_n726_));
  INV_X1    g525(.A(G43gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(G43gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n694_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g530(.A(G50gat), .ZN(new_n732_));
  INV_X1    g531(.A(new_n674_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n703_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n686_), .B(new_n357_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(KEYINPUT112), .ZN(new_n736_));
  OAI21_X1  g535(.A(G50gat), .B1(new_n735_), .B2(KEYINPUT112), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n734_), .B1(new_n736_), .B2(new_n737_), .ZN(G1331gat));
  NOR2_X1   g537(.A1(new_n486_), .A2(new_n516_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(new_n572_), .A3(new_n631_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT113), .ZN(new_n741_));
  INV_X1    g540(.A(G57gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n454_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n630_), .A2(new_n516_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n576_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n454_), .A3(new_n642_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G57gat), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n743_), .A2(new_n747_), .ZN(G1332gat));
  INV_X1    g547(.A(G64gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n741_), .A2(new_n749_), .A3(new_n712_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n745_), .A2(new_n642_), .A3(new_n712_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n751_), .A2(G64gat), .A3(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n751_), .B2(G64gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(G1333gat));
  NAND3_X1  g554(.A1(new_n741_), .A2(new_n204_), .A3(new_n725_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n745_), .A2(new_n725_), .A3(new_n642_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(G71gat), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n758_), .A2(KEYINPUT49), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n758_), .A2(KEYINPUT49), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(G1334gat));
  NAND3_X1  g560(.A1(new_n741_), .A2(new_n327_), .A3(new_n733_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n745_), .A2(new_n642_), .A3(new_n733_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(G78gat), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n764_), .A2(KEYINPUT50), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n764_), .A2(KEYINPUT50), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(G1335gat));
  NOR2_X1   g566(.A1(new_n577_), .A2(new_n697_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n739_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(G85gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(new_n454_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n679_), .A2(new_n516_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n572_), .A2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT115), .B1(new_n682_), .B2(new_n685_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n689_), .A2(new_n776_), .A3(new_n691_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n774_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n778_), .A2(new_n454_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n772_), .B1(new_n779_), .B2(new_n771_), .ZN(G1336gat));
  AOI21_X1  g579(.A(G92gat), .B1(new_n770_), .B2(new_n456_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n712_), .A2(new_n529_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT116), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n781_), .B1(new_n778_), .B2(new_n783_), .ZN(G1337gat));
  AOI21_X1  g583(.A(new_n206_), .B1(new_n778_), .B2(new_n725_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n725_), .A2(new_n525_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n769_), .A2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT51), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789_));
  INV_X1    g588(.A(new_n787_), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n290_), .B(new_n774_), .C1(new_n775_), .C2(new_n777_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n789_), .B(new_n790_), .C1(new_n791_), .C2(new_n206_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n788_), .A2(new_n792_), .ZN(G1338gat));
  AND2_X1   g592(.A1(new_n572_), .A2(new_n773_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n357_), .B(new_n794_), .C1(new_n682_), .C2(new_n685_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(new_n796_), .A3(G106gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n795_), .B2(G106gat), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n357_), .A2(new_n329_), .ZN(new_n799_));
  OAI22_X1  g598(.A1(new_n797_), .A2(new_n798_), .B1(new_n769_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT53), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802_));
  OAI221_X1 g601(.A(new_n802_), .B1(new_n769_), .B2(new_n799_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1339gat));
  INV_X1    g603(.A(G113gat), .ZN(new_n805_));
  INV_X1    g604(.A(new_n414_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n553_), .A2(new_n555_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n520_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n557_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n556_), .A2(KEYINPUT66), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n807_), .A2(new_n520_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n556_), .B2(KEYINPUT55), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n815_), .C2(new_n565_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n565_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n816_), .A2(new_n516_), .A3(new_n820_), .A4(new_n566_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n504_), .A2(new_n510_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n508_), .A2(new_n509_), .A3(new_n503_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n515_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n822_), .A2(new_n515_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n821_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT57), .B1(new_n827_), .B2(new_n656_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n829_), .B(new_n602_), .C1(new_n821_), .C2(new_n826_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n818_), .A2(KEYINPUT56), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n835_), .B(new_n817_), .C1(new_n815_), .C2(new_n565_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT120), .B1(new_n818_), .B2(KEYINPUT56), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n818_), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n834_), .A2(new_n836_), .A3(new_n837_), .A4(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n825_), .A2(new_n566_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n839_), .A2(KEYINPUT58), .A3(new_n840_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n610_), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n679_), .B1(new_n831_), .B2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n744_), .A2(new_n569_), .A3(new_n571_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n744_), .A2(new_n569_), .A3(new_n571_), .A4(KEYINPUT117), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n609_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n851_), .B2(new_n609_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n454_), .B(new_n806_), .C1(new_n846_), .C2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n805_), .B1(new_n856_), .B2(new_n517_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT121), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n859_), .B(new_n805_), .C1(new_n856_), .C2(new_n517_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n831_), .A2(new_n845_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n630_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n853_), .A2(new_n854_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n864_), .A2(KEYINPUT59), .A3(new_n454_), .A4(new_n806_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n856_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n517_), .A2(new_n805_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n858_), .A2(new_n860_), .B1(new_n868_), .B2(new_n869_), .ZN(G1340gat));
  AOI21_X1  g669(.A(new_n577_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n871_));
  INV_X1    g670(.A(G120gat), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n873_));
  AOI21_X1  g672(.A(G120gat), .B1(new_n572_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(KEYINPUT122), .B1(new_n873_), .B2(G120gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n874_), .B2(new_n877_), .ZN(new_n878_));
  OAI22_X1  g677(.A1(new_n871_), .A2(new_n872_), .B1(new_n856_), .B2(new_n878_), .ZN(G1341gat));
  INV_X1    g678(.A(G127gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n679_), .B2(KEYINPUT123), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(KEYINPUT123), .B2(new_n880_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n453_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(new_n806_), .A3(new_n679_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n868_), .A2(new_n882_), .B1(new_n884_), .B2(new_n880_), .ZN(G1342gat));
  AOI21_X1  g684(.A(new_n609_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n886_));
  INV_X1    g685(.A(G134gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n602_), .A2(new_n887_), .ZN(new_n888_));
  OAI22_X1  g687(.A1(new_n886_), .A2(new_n887_), .B1(new_n856_), .B2(new_n888_), .ZN(G1343gat));
  NOR2_X1   g688(.A1(new_n725_), .A2(new_n478_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n713_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n883_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(new_n315_), .A3(new_n516_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G141gat), .B1(new_n893_), .B2(new_n517_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1344gat));
  NAND3_X1  g696(.A1(new_n894_), .A2(new_n316_), .A3(new_n576_), .ZN(new_n898_));
  OAI21_X1  g697(.A(G148gat), .B1(new_n893_), .B2(new_n577_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1345gat));
  XNOR2_X1  g699(.A(KEYINPUT61), .B(G155gat), .ZN(new_n901_));
  OR3_X1    g700(.A1(new_n893_), .A2(new_n630_), .A3(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n893_), .B2(new_n630_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1346gat));
  NOR2_X1   g703(.A1(new_n609_), .A2(new_n299_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT124), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n883_), .A2(new_n602_), .A3(new_n892_), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n894_), .A2(new_n906_), .B1(new_n907_), .B2(new_n299_), .ZN(G1347gat));
  NOR2_X1   g707(.A1(new_n454_), .A2(new_n290_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n712_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n674_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n516_), .B(new_n913_), .C1(new_n846_), .C2(new_n855_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(G169gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT125), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n914_), .A2(new_n917_), .A3(G169gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n916_), .A2(KEYINPUT62), .A3(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n377_), .A2(new_n378_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n914_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n917_), .B1(new_n914_), .B2(G169gat), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n919_), .A2(new_n924_), .ZN(G1348gat));
  OAI211_X1 g724(.A(new_n572_), .B(new_n913_), .C1(new_n846_), .C2(new_n855_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n237_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n926_), .A2(KEYINPUT126), .A3(new_n237_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n357_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n577_), .A2(new_n237_), .A3(new_n910_), .ZN(new_n932_));
  AOI22_X1  g731(.A1(new_n929_), .A2(new_n930_), .B1(new_n931_), .B2(new_n932_), .ZN(G1349gat));
  NAND3_X1  g732(.A1(new_n931_), .A2(new_n679_), .A3(new_n911_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n219_), .A2(new_n221_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n912_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n630_), .A2(new_n247_), .A3(new_n368_), .ZN(new_n937_));
  AOI22_X1  g736(.A1(new_n934_), .A2(new_n935_), .B1(new_n936_), .B2(new_n937_), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n936_), .A2(new_n244_), .A3(new_n602_), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n936_), .A2(new_n610_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(new_n222_), .ZN(G1351gat));
  AND3_X1   g740(.A1(new_n712_), .A2(new_n453_), .A3(new_n890_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n864_), .A2(new_n516_), .A3(new_n942_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g743(.A1(new_n864_), .A2(new_n942_), .ZN(new_n945_));
  OAI21_X1  g744(.A(G204gat), .B1(new_n945_), .B2(new_n577_), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n864_), .A2(new_n337_), .A3(new_n576_), .A4(new_n942_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1353gat));
  NAND3_X1  g747(.A1(new_n864_), .A2(new_n679_), .A3(new_n942_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  AND2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n949_), .A2(new_n950_), .A3(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n952_), .B1(new_n949_), .B2(new_n950_), .ZN(G1354gat));
  OAI21_X1  g752(.A(G218gat), .B1(new_n945_), .B2(new_n609_), .ZN(new_n954_));
  OR2_X1    g753(.A1(new_n656_), .A2(G218gat), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n945_), .B2(new_n955_), .ZN(G1355gat));
endmodule


