//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n962_, new_n963_, new_n965_, new_n966_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n982_,
    new_n983_;
  NAND2_X1  g000(.A1(G127gat), .A2(G134gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G127gat), .A2(G134gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT82), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G113gat), .B(G120gat), .Z(new_n206_));
  INV_X1    g005(.A(G127gat), .ZN(new_n207_));
  INV_X1    g006(.A(G134gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(new_n202_), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n205_), .A2(new_n206_), .A3(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n206_), .B1(new_n205_), .B2(new_n211_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT83), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT30), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n205_), .A2(new_n206_), .A3(new_n211_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT83), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n214_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT25), .B(G183gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  AOI22_X1  g022(.A1(new_n220_), .A2(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n223_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT24), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT76), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT76), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n225_), .A2(new_n229_), .A3(KEYINPUT24), .A4(new_n226_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT23), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(G183gat), .A3(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n224_), .A2(new_n228_), .A3(new_n230_), .A4(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT77), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT22), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT78), .A4(G169gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G169gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT22), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(G169gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(new_n237_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT78), .B1(new_n242_), .B2(KEYINPUT77), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n240_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n226_), .B1(new_n247_), .B2(G176gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n232_), .A2(new_n234_), .A3(KEYINPUT79), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n231_), .A2(new_n252_), .A3(KEYINPUT23), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT80), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n249_), .A2(KEYINPUT80), .A3(new_n251_), .A4(new_n253_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n236_), .B1(new_n248_), .B2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n215_), .B1(new_n214_), .B2(new_n218_), .ZN(new_n260_));
  OR3_X1    g059(.A1(new_n219_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n219_), .B2(new_n260_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G71gat), .B(G99gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G227gat), .A2(G233gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n264_), .B(new_n265_), .Z(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n266_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n261_), .A2(new_n262_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT81), .B(G43gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT31), .B(G15gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n267_), .A2(new_n273_), .A3(new_n269_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n278_));
  INV_X1    g077(.A(G141gat), .ZN(new_n279_));
  INV_X1    g078(.A(G148gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT3), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n281_), .A2(new_n283_), .A3(new_n284_), .A4(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NOR3_X1   g088(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n286_), .B(new_n287_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G141gat), .B(G148gat), .Z(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(KEYINPUT1), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT85), .B1(new_n287_), .B2(KEYINPUT1), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT85), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(G155gat), .A4(G162gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n292_), .B1(new_n294_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n291_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n214_), .A2(new_n301_), .A3(new_n218_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n291_), .B(new_n300_), .C1(new_n212_), .C2(new_n213_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT94), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n214_), .A2(new_n301_), .A3(new_n305_), .A4(new_n218_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(KEYINPUT4), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT4), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n308_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G1gat), .B(G29gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(G85gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT0), .ZN(new_n316_));
  INV_X1    g115(.A(G57gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n304_), .A2(new_n312_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n313_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n312_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n304_), .A2(new_n311_), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n322_), .A2(new_n318_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT33), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n321_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT20), .ZN(new_n327_));
  INV_X1    g126(.A(new_n236_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n256_), .A2(new_n257_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n226_), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT77), .B1(new_n242_), .B2(new_n243_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT77), .B1(new_n238_), .B2(G169gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT78), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n239_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G176gat), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n330_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n328_), .B1(new_n329_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT89), .ZN(new_n339_));
  AND2_X1   g138(.A1(G211gat), .A2(G218gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G211gat), .A2(G218gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(G211gat), .ZN(new_n343_));
  INV_X1    g142(.A(G218gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G211gat), .A2(G218gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(KEYINPUT89), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(G197gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n349_), .A2(G204gat), .ZN(new_n350_));
  INV_X1    g149(.A(G204gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n351_), .A2(G197gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT21), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G197gat), .B(G204gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT21), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AND4_X1   g155(.A1(KEYINPUT88), .A2(new_n348_), .A3(new_n353_), .A4(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT88), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n342_), .B2(new_n347_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n353_), .B1(new_n359_), .B2(new_n356_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n327_), .B1(new_n338_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G226gat), .A2(G233gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT19), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT92), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n227_), .A2(new_n249_), .A3(new_n253_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n367_));
  AND2_X1   g166(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n368_));
  AND2_X1   g167(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n370_));
  OAI22_X1  g169(.A1(new_n367_), .A2(new_n368_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n223_), .A2(new_n222_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n366_), .A2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n250_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT91), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n226_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  AOI211_X1 g176(.A(KEYINPUT91), .B(new_n250_), .C1(new_n232_), .C2(new_n234_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n242_), .A2(new_n243_), .A3(new_n336_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n374_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n365_), .B1(new_n381_), .B2(new_n361_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n235_), .A2(new_n251_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n330_), .B1(new_n383_), .B2(KEYINPUT91), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n375_), .A2(new_n376_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n380_), .A3(new_n385_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n366_), .A2(new_n373_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n348_), .A2(KEYINPUT88), .ZN(new_n389_));
  INV_X1    g188(.A(new_n354_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(KEYINPUT21), .A3(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n359_), .A2(new_n353_), .A3(new_n356_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n388_), .A2(new_n393_), .A3(KEYINPUT92), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n362_), .A2(new_n364_), .A3(new_n382_), .A4(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT20), .B1(new_n388_), .B2(new_n393_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT93), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(new_n338_), .B2(new_n361_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n259_), .A2(KEYINPUT93), .A3(new_n393_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n396_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n395_), .B1(new_n400_), .B2(new_n364_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT18), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(G64gat), .ZN(new_n404_));
  INV_X1    g203(.A(G92gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n406_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n408_), .B(new_n395_), .C1(new_n400_), .C2(new_n364_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n319_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(KEYINPUT33), .A3(new_n318_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n326_), .A2(new_n407_), .A3(new_n409_), .A4(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n406_), .A2(KEYINPUT32), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT95), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n401_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n396_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n335_), .A2(new_n336_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n417_), .A2(new_n226_), .A3(new_n256_), .A4(new_n257_), .ZN(new_n418_));
  AOI221_X4 g217(.A(new_n397_), .B1(new_n391_), .B2(new_n392_), .C1(new_n418_), .C2(new_n236_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT93), .B1(new_n259_), .B2(new_n393_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n416_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n364_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT96), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n361_), .A2(new_n236_), .A3(new_n418_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n382_), .A2(KEYINPUT20), .A3(new_n394_), .A4(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n423_), .B1(new_n425_), .B2(new_n364_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n388_), .A2(new_n393_), .A3(KEYINPUT92), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT92), .B1(new_n388_), .B2(new_n393_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n364_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n429_), .A2(KEYINPUT96), .A3(new_n430_), .A4(new_n362_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n422_), .A2(new_n426_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n401_), .A2(KEYINPUT95), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n415_), .A2(new_n432_), .B1(new_n433_), .B2(new_n413_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT97), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n410_), .B2(new_n318_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n318_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n311_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n438_));
  OAI211_X1 g237(.A(KEYINPUT97), .B(new_n437_), .C1(new_n438_), .C2(new_n319_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n436_), .A2(new_n321_), .A3(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n412_), .B1(new_n434_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n301_), .A2(KEYINPUT29), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n393_), .ZN(new_n443_));
  INV_X1    g242(.A(G228gat), .ZN(new_n444_));
  INV_X1    g243(.A(G233gat), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n442_), .B(new_n393_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G78gat), .B(G106gat), .Z(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n453_), .B1(new_n301_), .B2(KEYINPUT29), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G22gat), .B(G50gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT29), .ZN(new_n456_));
  INV_X1    g255(.A(new_n453_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n291_), .A2(new_n300_), .A3(new_n456_), .A4(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(new_n455_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n455_), .B1(new_n454_), .B2(new_n458_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n447_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n452_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT90), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n452_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n449_), .A2(new_n465_), .A3(new_n451_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n462_), .A2(KEYINPUT87), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n460_), .A2(new_n471_), .A3(new_n461_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n464_), .B1(new_n469_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n441_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n436_), .A2(new_n321_), .A3(new_n439_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n476_), .A2(new_n474_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n422_), .A2(new_n426_), .A3(new_n431_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n408_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(KEYINPUT27), .A3(new_n407_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n407_), .A2(new_n409_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT27), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT98), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT98), .ZN(new_n484_));
  AOI211_X1 g283(.A(new_n484_), .B(KEYINPUT27), .C1(new_n407_), .C2(new_n409_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n477_), .B(new_n480_), .C1(new_n483_), .C2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n277_), .B1(new_n475_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT99), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AOI211_X1 g288(.A(KEYINPUT99), .B(new_n277_), .C1(new_n475_), .C2(new_n486_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n479_), .A2(KEYINPUT27), .A3(new_n407_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n409_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n421_), .A2(new_n430_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n408_), .B1(new_n493_), .B2(new_n395_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n482_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n484_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n481_), .A2(KEYINPUT98), .A3(new_n482_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n491_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n277_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n474_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n498_), .A2(new_n501_), .A3(new_n440_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n489_), .A2(new_n490_), .A3(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(G57gat), .A2(G64gat), .ZN(new_n505_));
  NOR2_X1   g304(.A1(G57gat), .A2(G64gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT11), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n507_), .A2(new_n508_), .B1(G71gat), .B2(G78gat), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT67), .B1(new_n507_), .B2(new_n508_), .ZN(new_n510_));
  INV_X1    g309(.A(G71gat), .ZN(new_n511_));
  INV_X1    g310(.A(G78gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT67), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n514_), .B(KEYINPUT11), .C1(new_n505_), .C2(new_n506_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n509_), .A2(new_n510_), .A3(new_n513_), .A4(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G71gat), .A2(G78gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G57gat), .B(G64gat), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n513_), .B(new_n517_), .C1(new_n518_), .C2(KEYINPUT11), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n514_), .B1(new_n518_), .B2(KEYINPUT11), .ZN(new_n520_));
  INV_X1    g319(.A(new_n515_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n516_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G85gat), .B(G92gat), .Z(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT9), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT6), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT6), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(G99gat), .A3(G106gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G106gat), .ZN(new_n532_));
  INV_X1    g331(.A(G99gat), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n533_), .A2(KEYINPUT10), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(KEYINPUT10), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n532_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n405_), .A2(KEYINPUT9), .ZN(new_n537_));
  OR2_X1    g336(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n526_), .A2(new_n531_), .A3(new_n536_), .A4(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT66), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT10), .B(G99gat), .Z(new_n544_));
  AOI22_X1  g343(.A1(new_n544_), .A2(new_n532_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n545_), .A2(KEYINPUT66), .A3(new_n526_), .A4(new_n540_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n548_));
  OR3_X1    g347(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n531_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT8), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n550_), .A2(new_n551_), .A3(new_n525_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n551_), .B1(new_n550_), .B2(new_n525_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n524_), .B1(new_n547_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n525_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT8), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n550_), .A2(new_n551_), .A3(new_n525_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n559_), .A2(new_n523_), .A3(new_n546_), .A4(new_n543_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n555_), .A2(KEYINPUT12), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT12), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n562_), .B(new_n524_), .C1(new_n547_), .C2(new_n554_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT64), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n555_), .A2(KEYINPUT68), .A3(new_n560_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n569_), .B(new_n566_), .C1(KEYINPUT68), .C2(new_n560_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G120gat), .B(G148gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT5), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G176gat), .B(G204gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n575_), .B(new_n576_), .Z(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n571_), .B(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT13), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT13), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT75), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G29gat), .B(G36gat), .ZN(new_n584_));
  INV_X1    g383(.A(G43gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(G50gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT15), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G15gat), .B(G22gat), .ZN(new_n590_));
  INV_X1    g389(.A(G1gat), .ZN(new_n591_));
  INV_X1    g390(.A(G8gat), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT14), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n590_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G1gat), .B(G8gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n589_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598_));
  INV_X1    g397(.A(new_n596_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n588_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n597_), .A2(new_n598_), .A3(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n588_), .B(new_n599_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(G229gat), .A3(G233gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT74), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(new_n241_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(new_n349_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n601_), .A2(new_n603_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n607_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n583_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n610_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(KEYINPUT75), .A3(new_n608_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n504_), .A2(new_n582_), .A3(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n547_), .A2(new_n554_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n589_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n588_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT34), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(KEYINPUT35), .A3(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n622_), .B(KEYINPUT35), .Z(new_n624_));
  NAND3_X1  g423(.A1(new_n618_), .A2(new_n619_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT71), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT71), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n618_), .A2(new_n627_), .A3(new_n619_), .A4(new_n624_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n623_), .A2(new_n626_), .A3(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G190gat), .B(G218gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(G134gat), .ZN(new_n631_));
  INV_X1    g430(.A(G162gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(KEYINPUT36), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n629_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n633_), .B(KEYINPUT36), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n629_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(KEYINPUT37), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT72), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n629_), .A2(KEYINPUT72), .A3(new_n638_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n642_), .A2(new_n637_), .A3(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n644_), .B2(KEYINPUT37), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n523_), .B(new_n596_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(G231gat), .A2(G233gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G127gat), .B(G155gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT16), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(G183gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(new_n343_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n648_), .B1(KEYINPUT17), .B2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT73), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT17), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n656_), .B2(new_n652_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n654_), .A2(KEYINPUT73), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n654_), .A2(KEYINPUT73), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n658_), .A2(KEYINPUT17), .A3(new_n653_), .A4(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n657_), .A2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n645_), .A2(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n615_), .A2(new_n662_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n663_), .A2(new_n591_), .A3(new_n476_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT38), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(KEYINPUT38), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n666_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n504_), .A2(new_n644_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n661_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n612_), .A2(new_n608_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n582_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n670_), .A2(new_n671_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G1gat), .B1(new_n675_), .B2(new_n440_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .A4(new_n676_), .ZN(G1324gat));
  INV_X1    g476(.A(new_n498_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n663_), .A2(new_n592_), .A3(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G8gat), .B1(new_n675_), .B2(new_n498_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT101), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT39), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n683_), .B(G8gat), .C1(new_n675_), .C2(new_n498_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n681_), .A2(new_n682_), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n682_), .B1(new_n681_), .B2(new_n684_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n679_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT40), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT40), .B(new_n679_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1325gat));
  INV_X1    g490(.A(G15gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n674_), .ZN(new_n693_));
  NOR4_X1   g492(.A1(new_n504_), .A2(new_n644_), .A3(new_n661_), .A4(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n692_), .B1(new_n694_), .B2(new_n277_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT41), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n663_), .A2(new_n692_), .A3(new_n277_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT102), .ZN(G1326gat));
  INV_X1    g498(.A(G22gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n694_), .B2(new_n500_), .ZN(new_n701_));
  XOR2_X1   g500(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n663_), .A2(new_n700_), .A3(new_n500_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT104), .Z(G1327gat));
  OAI211_X1 g505(.A(new_n642_), .B(new_n643_), .C1(new_n636_), .C2(new_n629_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n671_), .A2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n615_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(G29gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n476_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n640_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT37), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n707_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT43), .B1(new_n504_), .B2(new_n714_), .ZN(new_n715_));
  AOI22_X1  g514(.A1(new_n498_), .A2(new_n477_), .B1(new_n474_), .B2(new_n441_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT99), .B1(new_n716_), .B2(new_n277_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n487_), .A2(new_n488_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n502_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n645_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n715_), .A2(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n693_), .A2(new_n671_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n722_), .A2(KEYINPUT44), .A3(new_n723_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(new_n476_), .A3(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n711_), .B1(new_n728_), .B2(new_n710_), .ZN(G1328gat));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n730_));
  XOR2_X1   g529(.A(KEYINPUT106), .B(KEYINPUT46), .Z(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n726_), .A2(new_n678_), .A3(new_n727_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(G36gat), .ZN(new_n734_));
  INV_X1    g533(.A(G36gat), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n709_), .A2(new_n735_), .A3(new_n678_), .A4(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n615_), .A2(new_n735_), .A3(new_n708_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n736_), .B1(new_n739_), .B2(new_n498_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n730_), .B(new_n732_), .C1(new_n734_), .C2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(G36gat), .B2(new_n733_), .ZN(new_n743_));
  OAI21_X1  g542(.A(KEYINPUT107), .B1(new_n743_), .B2(new_n731_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(KEYINPUT46), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n742_), .A2(new_n744_), .A3(new_n745_), .ZN(G1329gat));
  NAND3_X1  g545(.A1(new_n709_), .A2(new_n585_), .A3(new_n277_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n726_), .A2(new_n277_), .A3(new_n727_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n585_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(G1330gat));
  NAND3_X1  g550(.A1(new_n709_), .A2(new_n587_), .A3(new_n500_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n726_), .A2(new_n500_), .A3(new_n727_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(new_n754_), .A3(G50gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n753_), .B2(G50gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(G1331gat));
  AND3_X1   g556(.A1(new_n657_), .A2(new_n614_), .A3(new_n660_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n670_), .A2(new_n582_), .A3(new_n758_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n759_), .A2(new_n317_), .A3(new_n440_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n582_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n504_), .A2(new_n761_), .A3(new_n672_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(new_n662_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n476_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n760_), .B1(new_n317_), .B2(new_n764_), .ZN(G1332gat));
  OAI21_X1  g564(.A(G64gat), .B1(new_n759_), .B2(new_n498_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT48), .ZN(new_n767_));
  INV_X1    g566(.A(G64gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n763_), .A2(new_n768_), .A3(new_n678_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1333gat));
  OAI21_X1  g569(.A(G71gat), .B1(new_n759_), .B2(new_n499_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT49), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n763_), .A2(new_n511_), .A3(new_n277_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1334gat));
  NAND3_X1  g573(.A1(new_n763_), .A2(new_n512_), .A3(new_n500_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G78gat), .B1(new_n759_), .B2(new_n474_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT109), .Z(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(KEYINPUT50), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(KEYINPUT50), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1335gat));
  AND2_X1   g579(.A1(new_n762_), .A2(new_n708_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G85gat), .B1(new_n781_), .B2(new_n476_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n761_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n722_), .A2(new_n783_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n476_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n782_), .B1(new_n784_), .B2(new_n785_), .ZN(G1336gat));
  AOI21_X1  g585(.A(new_n405_), .B1(new_n784_), .B2(new_n678_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n498_), .A2(G92gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n781_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(G1337gat));
  AOI21_X1  g590(.A(new_n533_), .B1(new_n784_), .B2(new_n277_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n277_), .A2(new_n544_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n781_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n794_), .B(new_n795_), .ZN(G1338gat));
  AND3_X1   g595(.A1(new_n719_), .A2(new_n720_), .A3(new_n645_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n720_), .B1(new_n719_), .B2(new_n645_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n500_), .B(new_n783_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT111), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n722_), .A2(new_n801_), .A3(new_n500_), .A4(new_n783_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n802_), .A3(G106gat), .ZN(new_n803_));
  XOR2_X1   g602(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n804_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n800_), .A2(new_n802_), .A3(G106gat), .A4(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n781_), .A2(new_n532_), .A3(new_n500_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT53), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n808_), .A2(new_n812_), .A3(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1339gat));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n611_), .A2(new_n613_), .A3(G113gat), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n498_), .A2(new_n476_), .A3(new_n501_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n568_), .A2(new_n821_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n566_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT115), .B1(new_n825_), .B2(new_n822_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n561_), .A2(new_n566_), .A3(new_n563_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(KEYINPUT55), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n824_), .A2(new_n826_), .A3(new_n827_), .A4(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(KEYINPUT56), .A3(new_n578_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n578_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT117), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n832_), .A2(new_n836_), .A3(new_n833_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n831_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n607_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n602_), .A2(new_n598_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n597_), .A2(new_n600_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n839_), .B(new_n840_), .C1(new_n841_), .C2(new_n598_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n842_), .A2(new_n608_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n571_), .A2(new_n577_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT116), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n843_), .A2(new_n847_), .A3(new_n844_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n820_), .B1(new_n838_), .B2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n836_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n851_));
  AOI211_X1 g650(.A(KEYINPUT117), .B(KEYINPUT56), .C1(new_n829_), .C2(new_n578_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n830_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n846_), .A2(new_n848_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(KEYINPUT58), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n850_), .A2(new_n645_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n672_), .A2(new_n844_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n834_), .B2(new_n830_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n843_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n579_), .A2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n707_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n856_), .A2(KEYINPUT120), .A3(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n861_), .A2(new_n862_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT120), .B1(new_n856_), .B2(new_n863_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n661_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n758_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT113), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n761_), .A2(new_n872_), .A3(new_n758_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n645_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n819_), .B1(new_n869_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n850_), .A2(new_n879_), .A3(new_n645_), .A4(new_n855_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n880_), .A2(new_n863_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n865_), .B1(new_n856_), .B2(KEYINPUT118), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n671_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n871_), .A2(new_n873_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n875_), .B1(new_n884_), .B2(new_n714_), .ZN(new_n885_));
  AOI211_X1 g684(.A(KEYINPUT54), .B(new_n645_), .C1(new_n871_), .C2(new_n873_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n878_), .B1(new_n883_), .B2(new_n887_), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n853_), .A2(KEYINPUT58), .A3(new_n854_), .ZN(new_n889_));
  AOI21_X1  g688(.A(KEYINPUT58), .B1(new_n853_), .B2(new_n854_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n889_), .A2(new_n890_), .A3(new_n714_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n866_), .B1(new_n891_), .B2(new_n879_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n880_), .A2(new_n863_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n661_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(new_n876_), .A3(KEYINPUT119), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n888_), .A2(new_n895_), .A3(new_n817_), .ZN(new_n896_));
  AOI211_X1 g695(.A(new_n816_), .B(new_n877_), .C1(new_n896_), .C2(KEYINPUT59), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n888_), .A2(new_n895_), .A3(new_n672_), .A4(new_n817_), .ZN(new_n898_));
  INV_X1    g697(.A(G113gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n815_), .B1(new_n897_), .B2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n896_), .A2(KEYINPUT59), .ZN(new_n903_));
  INV_X1    g702(.A(new_n877_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  OAI211_X1 g704(.A(KEYINPUT121), .B(new_n900_), .C1(new_n905_), .C2(new_n816_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n902_), .A2(new_n906_), .ZN(G1340gat));
  AOI21_X1  g706(.A(new_n877_), .B1(new_n896_), .B2(KEYINPUT59), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n761_), .B2(G120gat), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n888_), .A2(new_n895_), .A3(new_n817_), .A4(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n908_), .A2(new_n582_), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(G120gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(KEYINPUT60), .B2(new_n911_), .ZN(G1341gat));
  OAI21_X1  g713(.A(G127gat), .B1(new_n905_), .B2(new_n661_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n896_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n916_), .A2(new_n207_), .A3(new_n671_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(G1342gat));
  AOI21_X1  g717(.A(G134gat), .B1(new_n916_), .B2(new_n644_), .ZN(new_n919_));
  XOR2_X1   g718(.A(KEYINPUT122), .B(G134gat), .Z(new_n920_));
  NOR2_X1   g719(.A1(new_n714_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n908_), .B2(new_n921_), .ZN(G1343gat));
  AND2_X1   g721(.A1(new_n888_), .A2(new_n895_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n277_), .A2(new_n474_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n498_), .A2(new_n476_), .A3(new_n924_), .ZN(new_n925_));
  XOR2_X1   g724(.A(new_n925_), .B(KEYINPUT123), .Z(new_n926_));
  AND2_X1   g725(.A1(new_n923_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n672_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(G141gat), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n927_), .A2(new_n279_), .A3(new_n672_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1344gat));
  NAND2_X1  g730(.A1(new_n927_), .A2(new_n582_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(G148gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n927_), .A2(new_n280_), .A3(new_n582_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1345gat));
  NAND3_X1  g734(.A1(new_n923_), .A2(new_n671_), .A3(new_n926_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT61), .B(G155gat), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n936_), .B(new_n937_), .ZN(G1346gat));
  NAND2_X1  g737(.A1(new_n927_), .A2(new_n644_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n714_), .A2(new_n632_), .ZN(new_n940_));
  AOI22_X1  g739(.A1(new_n939_), .A2(new_n632_), .B1(new_n927_), .B2(new_n940_), .ZN(G1347gat));
  NOR2_X1   g740(.A1(new_n498_), .A2(new_n476_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n501_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n943_), .B1(new_n869_), .B2(new_n876_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n672_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(G169gat), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n946_), .A2(KEYINPUT124), .A3(new_n947_), .ZN(new_n948_));
  OR2_X1    g747(.A1(new_n947_), .A2(KEYINPUT124), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n947_), .A2(KEYINPUT124), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n945_), .A2(G169gat), .A3(new_n949_), .A4(new_n950_), .ZN(new_n951_));
  OAI211_X1 g750(.A(new_n948_), .B(new_n951_), .C1(new_n244_), .C2(new_n945_), .ZN(G1348gat));
  AOI21_X1  g751(.A(G176gat), .B1(new_n944_), .B2(new_n582_), .ZN(new_n953_));
  AND2_X1   g752(.A1(new_n923_), .A2(new_n582_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n943_), .A2(new_n336_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n953_), .B1(new_n954_), .B2(new_n955_), .ZN(G1349gat));
  INV_X1    g755(.A(new_n944_), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n957_), .A2(new_n661_), .A3(new_n220_), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n923_), .A2(new_n671_), .A3(new_n501_), .A4(new_n942_), .ZN(new_n959_));
  INV_X1    g758(.A(G183gat), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n958_), .B1(new_n959_), .B2(new_n960_), .ZN(G1350gat));
  OAI21_X1  g760(.A(G190gat), .B1(new_n957_), .B2(new_n714_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n944_), .A2(new_n644_), .A3(new_n221_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(G1351gat));
  NAND4_X1  g763(.A1(new_n888_), .A2(new_n895_), .A3(new_n924_), .A4(new_n942_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n965_), .A2(new_n673_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(new_n349_), .ZN(G1352gat));
  NOR2_X1   g766(.A1(new_n965_), .A2(new_n761_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(new_n351_), .ZN(G1353gat));
  AND3_X1   g768(.A1(new_n888_), .A2(new_n895_), .A3(new_n924_), .ZN(new_n970_));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971_));
  INV_X1    g770(.A(KEYINPUT63), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n671_), .B1(new_n972_), .B2(new_n343_), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n973_), .B(KEYINPUT125), .ZN(new_n974_));
  INV_X1    g773(.A(new_n974_), .ZN(new_n975_));
  NAND4_X1  g774(.A1(new_n970_), .A2(new_n971_), .A3(new_n942_), .A4(new_n975_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n977_));
  OAI21_X1  g776(.A(KEYINPUT126), .B1(new_n965_), .B2(new_n974_), .ZN(new_n978_));
  AND3_X1   g777(.A1(new_n976_), .A2(new_n977_), .A3(new_n978_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n977_), .B1(new_n976_), .B2(new_n978_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n979_), .A2(new_n980_), .ZN(G1354gat));
  NOR3_X1   g780(.A1(new_n965_), .A2(new_n344_), .A3(new_n714_), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n970_), .A2(new_n644_), .A3(new_n942_), .ZN(new_n983_));
  AOI21_X1  g782(.A(new_n982_), .B1(new_n983_), .B2(new_n344_), .ZN(G1355gat));
endmodule


