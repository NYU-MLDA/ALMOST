//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n844_, new_n845_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(G85gat), .B(G92gat), .Z(new_n204_));
  INV_X1    g003(.A(KEYINPUT7), .ZN(new_n205_));
  INV_X1    g004(.A(G99gat), .ZN(new_n206_));
  INV_X1    g005(.A(G106gat), .ZN(new_n207_));
  NAND4_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .A4(KEYINPUT64), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209_));
  OAI22_X1  g008(.A1(new_n209_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n209_), .A2(KEYINPUT7), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n204_), .B1(new_n211_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT8), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n204_), .B(new_n220_), .C1(new_n211_), .C2(new_n217_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n204_), .A2(KEYINPUT9), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT10), .B(G99gat), .Z(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n207_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n214_), .A2(new_n215_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT9), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(G85gat), .A3(G92gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .A4(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n235_));
  XOR2_X1   g034(.A(G71gat), .B(G78gat), .Z(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n235_), .A2(new_n236_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n224_), .A2(new_n231_), .A3(new_n239_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(KEYINPUT12), .A3(new_n242_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n227_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n222_), .A2(new_n223_), .B1(new_n244_), .B2(new_n225_), .ZN(new_n245_));
  OR3_X1    g044(.A1(new_n245_), .A2(KEYINPUT12), .A3(new_n239_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n203_), .B1(new_n243_), .B2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n202_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G120gat), .B(G148gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G204gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT5), .B(G176gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n249_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT13), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n249_), .A2(new_n254_), .ZN(new_n258_));
  OR3_X1    g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n257_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT66), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G15gat), .B(G22gat), .ZN(new_n268_));
  INV_X1    g067(.A(G1gat), .ZN(new_n269_));
  INV_X1    g068(.A(G8gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT14), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G1gat), .B(G8gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G29gat), .B(G36gat), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G43gat), .B(G50gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G43gat), .B(G50gat), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n275_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n274_), .A2(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n278_), .A2(new_n280_), .A3(KEYINPUT15), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT15), .B1(new_n278_), .B2(new_n280_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n282_), .B1(new_n286_), .B2(new_n274_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G229gat), .A2(G233gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n288_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n274_), .A2(new_n281_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(new_n282_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G169gat), .B(G197gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G113gat), .B(G141gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n295_), .B(new_n296_), .Z(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n289_), .A2(new_n292_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT78), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n298_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n302_));
  OR3_X1    g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n301_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G127gat), .B(G155gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G211gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(KEYINPUT16), .B(G183gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G231gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n274_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(new_n239_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n310_), .B1(new_n314_), .B2(KEYINPUT17), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(KEYINPUT17), .B2(new_n310_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(KEYINPUT75), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n267_), .A2(new_n306_), .A3(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(KEYINPUT67), .B(KEYINPUT34), .Z(new_n321_));
  NAND2_X1  g120(.A1(G232gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n245_), .A2(new_n285_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n232_), .A2(new_n281_), .ZN(new_n325_));
  OAI211_X1 g124(.A(KEYINPUT35), .B(new_n323_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n245_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n286_), .A2(new_n232_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(KEYINPUT35), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n323_), .A2(KEYINPUT35), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .A4(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n326_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT72), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G190gat), .B(G218gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(G134gat), .B(G162gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT36), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT36), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(KEYINPUT68), .B(KEYINPUT69), .Z(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n326_), .A2(new_n331_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT70), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n326_), .A2(new_n331_), .A3(KEYINPUT70), .A4(new_n342_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n334_), .A2(new_n338_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n346_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT71), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n332_), .A2(new_n338_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT71), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n345_), .A2(new_n353_), .A3(new_n346_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n351_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT37), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n349_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT74), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n349_), .B(new_n359_), .C1(new_n355_), .C2(new_n356_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT1), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT85), .ZN(new_n364_));
  OR2_X1    g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT85), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n362_), .A2(new_n366_), .A3(KEYINPUT1), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT86), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n362_), .A2(KEYINPUT1), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT86), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n364_), .A2(new_n371_), .A3(new_n365_), .A4(new_n367_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n369_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G141gat), .A2(G148gat), .ZN(new_n374_));
  OR2_X1    g173(.A1(G141gat), .A2(G148gat), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT87), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n365_), .A2(new_n362_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT90), .B1(new_n374_), .B2(KEYINPUT89), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT2), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n374_), .B2(KEYINPUT90), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n381_), .B1(new_n383_), .B2(new_n380_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT88), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n375_), .B(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n379_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT91), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  OAI211_X1 g189(.A(KEYINPUT91), .B(new_n379_), .C1(new_n384_), .C2(new_n387_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n373_), .A2(KEYINPUT87), .A3(new_n374_), .A4(new_n375_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n378_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G127gat), .B(G134gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G113gat), .B(G120gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n397_), .A2(KEYINPUT83), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n396_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n394_), .A2(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n378_), .A2(new_n392_), .A3(new_n397_), .A4(new_n393_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT4), .B1(new_n394_), .B2(new_n401_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n408_), .B1(new_n404_), .B2(KEYINPUT4), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n409_), .B2(new_n406_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411_));
  INV_X1    g210(.A(G85gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT0), .B(G57gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n413_), .B(new_n414_), .Z(new_n415_));
  NAND2_X1  g214(.A1(new_n410_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT105), .ZN(new_n417_));
  INV_X1    g216(.A(new_n415_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n407_), .B(new_n418_), .C1(new_n409_), .C2(new_n406_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n416_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  OR3_X1    g219(.A1(new_n410_), .A2(new_n417_), .A3(new_n415_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT25), .B(G183gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT26), .B(G190gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G183gat), .A2(G190gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT23), .ZN(new_n427_));
  INV_X1    g226(.A(G169gat), .ZN(new_n428_));
  INV_X1    g227(.A(G176gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n430_), .A2(KEYINPUT24), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n425_), .A2(new_n427_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G169gat), .A2(G176gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT24), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n432_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n427_), .B1(G183gat), .B2(G190gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(G176gat), .B1(KEYINPUT79), .B2(KEYINPUT22), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(G169gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G197gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G204gat), .ZN(new_n443_));
  INV_X1    g242(.A(G204gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G197gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT21), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT93), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT92), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n445_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n443_), .A2(new_n449_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT21), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G211gat), .B(G218gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n448_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n454_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT21), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n441_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT97), .B1(new_n434_), .B2(KEYINPUT24), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT97), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n430_), .B1(new_n435_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n432_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT22), .B(G169gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT98), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n464_), .A2(new_n429_), .B1(new_n465_), .B2(new_n434_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n437_), .B(new_n466_), .C1(new_n465_), .C2(new_n434_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n458_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n459_), .B(KEYINPUT20), .C1(new_n468_), .C2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G226gat), .A2(G233gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT19), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n468_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT99), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n441_), .B2(new_n458_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n475_), .A2(KEYINPUT99), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n473_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n474_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G64gat), .B(G92gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT101), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT102), .B(G36gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(new_n270_), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n486_), .B(new_n488_), .Z(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n482_), .B(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(KEYINPUT27), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT27), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n475_), .A2(new_n478_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n472_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n496_), .A2(new_n490_), .ZN(new_n497_));
  AOI211_X1 g296(.A(new_n493_), .B(new_n497_), .C1(new_n489_), .C2(new_n482_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n492_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT96), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n394_), .A2(KEYINPUT29), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n458_), .ZN(new_n502_));
  INV_X1    g301(.A(G228gat), .ZN(new_n503_));
  INV_X1    g302(.A(G233gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n505_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n501_), .A2(new_n458_), .A3(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G78gat), .B(G106gat), .Z(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(KEYINPUT95), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n506_), .A2(new_n508_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n507_), .B1(new_n501_), .B2(new_n458_), .ZN(new_n513_));
  AOI211_X1 g312(.A(new_n469_), .B(new_n505_), .C1(new_n394_), .C2(KEYINPUT29), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n510_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n512_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT28), .B(G22gat), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT29), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n378_), .A2(new_n392_), .A3(new_n519_), .A4(new_n393_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(G50gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n520_), .A2(G50gat), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n518_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n523_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(new_n517_), .A3(new_n521_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n500_), .B1(new_n516_), .B2(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n524_), .A2(new_n526_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n529_), .A2(KEYINPUT96), .A3(new_n512_), .A4(new_n515_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G227gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT81), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT82), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G15gat), .B(G43gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n536_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G71gat), .B(G99gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n441_), .B(new_n540_), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n441_), .B(new_n540_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n536_), .A2(new_n538_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n536_), .A2(new_n538_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n542_), .A2(KEYINPUT84), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT31), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT31), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n542_), .A2(KEYINPUT84), .A3(new_n549_), .A4(new_n546_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n401_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n401_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n548_), .A2(new_n553_), .A3(new_n550_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n506_), .A2(KEYINPUT94), .A3(new_n508_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT94), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n509_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n556_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n557_), .B(new_n509_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n527_), .A3(new_n561_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n531_), .A2(new_n555_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n555_), .B1(new_n531_), .B2(new_n562_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n422_), .B(new_n499_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n406_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n405_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n409_), .A2(new_n566_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT104), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT4), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n571_));
  OAI211_X1 g370(.A(KEYINPUT104), .B(new_n406_), .C1(new_n571_), .C2(new_n408_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n415_), .B(new_n567_), .C1(new_n569_), .C2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n419_), .A2(KEYINPUT103), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT33), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT33), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n419_), .A2(KEYINPUT103), .A3(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n574_), .A2(new_n576_), .A3(new_n578_), .A4(new_n491_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT32), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n482_), .B1(new_n580_), .B2(new_n490_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n496_), .A2(KEYINPUT32), .A3(new_n489_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n420_), .A2(new_n421_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n531_), .A2(new_n562_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(new_n555_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n565_), .A2(new_n587_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n320_), .A2(new_n361_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n422_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n269_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT107), .Z(new_n594_));
  NOR2_X1   g393(.A1(new_n591_), .A2(new_n592_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT106), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n320_), .A2(new_n588_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n347_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n599_), .A2(new_n590_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n594_), .B(new_n596_), .C1(new_n269_), .C2(new_n600_), .ZN(G1324gat));
  INV_X1    g400(.A(new_n499_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n589_), .A2(new_n270_), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n597_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n604_), .A2(new_n605_), .A3(G8gat), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n605_), .B1(new_n604_), .B2(G8gat), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n603_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g408(.A(G15gat), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n589_), .A2(new_n610_), .A3(new_n555_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n599_), .A2(new_n555_), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n612_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT41), .B1(new_n612_), .B2(G15gat), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n611_), .B1(new_n613_), .B2(new_n614_), .ZN(G1326gat));
  INV_X1    g414(.A(G22gat), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n589_), .A2(new_n616_), .A3(new_n585_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n599_), .A2(new_n585_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(G22gat), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n619_), .A2(KEYINPUT42), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(KEYINPUT42), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n617_), .B1(new_n620_), .B2(new_n621_), .ZN(G1327gat));
  AOI21_X1  g421(.A(new_n598_), .B1(new_n565_), .B2(new_n587_), .ZN(new_n623_));
  AOI211_X1 g422(.A(new_n306_), .B(new_n318_), .C1(new_n263_), .C2(new_n265_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT110), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT110), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n623_), .A2(new_n624_), .A3(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(G29gat), .B1(new_n629_), .B2(new_n590_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT108), .ZN(new_n631_));
  AOI221_X4 g430(.A(new_n361_), .B1(new_n631_), .B2(KEYINPUT43), .C1(new_n565_), .C2(new_n587_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n358_), .A2(KEYINPUT108), .A3(new_n360_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT43), .ZN(new_n634_));
  INV_X1    g433(.A(new_n361_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n588_), .B2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n624_), .B1(new_n632_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT109), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n637_), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n422_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n630_), .B1(new_n642_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g442(.A(G36gat), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n626_), .A2(new_n644_), .A3(new_n628_), .A4(new_n602_), .ZN(new_n645_));
  XOR2_X1   g444(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n499_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n648_), .B2(new_n644_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT46), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(KEYINPUT46), .B(new_n647_), .C1(new_n648_), .C2(new_n644_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1329gat));
  INV_X1    g452(.A(KEYINPUT47), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n637_), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT44), .B1(new_n637_), .B2(KEYINPUT109), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n555_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(G43gat), .ZN(new_n658_));
  INV_X1    g457(.A(G43gat), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n629_), .A2(new_n659_), .A3(new_n555_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n654_), .B1(new_n658_), .B2(new_n661_), .ZN(new_n662_));
  AOI211_X1 g461(.A(KEYINPUT47), .B(new_n660_), .C1(new_n657_), .C2(G43gat), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1330gat));
  INV_X1    g463(.A(G50gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n629_), .A2(new_n665_), .A3(new_n585_), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n640_), .A2(new_n641_), .B1(new_n562_), .B2(new_n531_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n667_), .B2(new_n665_), .ZN(G1331gat));
  NAND3_X1  g467(.A1(new_n267_), .A2(new_n361_), .A3(new_n318_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT112), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n305_), .B1(new_n565_), .B2(new_n587_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT113), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n670_), .A2(KEYINPUT113), .A3(new_n671_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G57gat), .B1(new_n676_), .B2(new_n590_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n319_), .A2(new_n305_), .ZN(new_n678_));
  AND4_X1   g477(.A1(new_n598_), .A2(new_n588_), .A3(new_n267_), .A4(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(G57gat), .A3(new_n590_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT114), .Z(new_n681_));
  NOR2_X1   g480(.A1(new_n677_), .A2(new_n681_), .ZN(G1332gat));
  NOR2_X1   g481(.A1(new_n499_), .A2(G64gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n674_), .A2(new_n675_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n679_), .A2(new_n602_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G64gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(KEYINPUT48), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(KEYINPUT48), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT115), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1333gat));
  INV_X1    g490(.A(G71gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n676_), .A2(new_n692_), .A3(new_n555_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n679_), .B2(new_n555_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT49), .Z(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1334gat));
  INV_X1    g495(.A(G78gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n676_), .A2(new_n697_), .A3(new_n585_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n679_), .B2(new_n585_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT50), .Z(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1335gat));
  NOR3_X1   g500(.A1(new_n266_), .A2(new_n305_), .A3(new_n318_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n623_), .A2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G85gat), .B1(new_n703_), .B2(new_n590_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n632_), .A2(new_n636_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(new_n702_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n422_), .A2(new_n412_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(G1336gat));
  AOI21_X1  g507(.A(G92gat), .B1(new_n703_), .B2(new_n602_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n602_), .A2(G92gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n706_), .B2(new_n710_), .ZN(G1337gat));
  AOI21_X1  g510(.A(new_n206_), .B1(new_n706_), .B2(new_n555_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n703_), .A2(new_n226_), .A3(new_n555_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT51), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(G1338gat));
  OAI211_X1 g516(.A(new_n585_), .B(new_n702_), .C1(new_n632_), .C2(new_n636_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G106gat), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT52), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n703_), .A2(new_n207_), .A3(new_n585_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n720_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1339gat));
  NAND3_X1  g525(.A1(new_n361_), .A2(new_n262_), .A3(new_n678_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT54), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT120), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT55), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n243_), .A2(new_n246_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(new_n202_), .ZN(new_n732_));
  AOI211_X1 g531(.A(KEYINPUT55), .B(new_n203_), .C1(new_n243_), .C2(new_n246_), .ZN(new_n733_));
  OAI22_X1  g532(.A1(new_n732_), .A2(new_n733_), .B1(new_n202_), .B2(new_n731_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n253_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT56), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT56), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n734_), .A2(new_n737_), .A3(new_n253_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n736_), .A2(new_n305_), .A3(new_n255_), .A4(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n287_), .A2(new_n290_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n288_), .B1(new_n291_), .B2(new_n282_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n297_), .A3(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n299_), .A2(new_n742_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT117), .Z(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n739_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n598_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT57), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n736_), .A2(new_n255_), .A3(new_n744_), .A4(new_n738_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT58), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n635_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT119), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT118), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n746_), .B2(new_n598_), .ZN(new_n755_));
  AOI211_X1 g554(.A(KEYINPUT118), .B(new_n347_), .C1(new_n739_), .C2(new_n745_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n753_), .B1(new_n757_), .B2(new_n748_), .ZN(new_n758_));
  NOR4_X1   g557(.A1(new_n755_), .A2(new_n756_), .A3(KEYINPUT119), .A4(KEYINPUT57), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n729_), .B(new_n752_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n319_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n747_), .A2(KEYINPUT118), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n746_), .A2(new_n754_), .A3(new_n598_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n748_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT119), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n757_), .A2(new_n753_), .A3(new_n748_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n729_), .B1(new_n767_), .B2(new_n752_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n728_), .B1(new_n761_), .B2(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n602_), .A2(new_n422_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(new_n563_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(G113gat), .B1(new_n772_), .B2(new_n305_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT59), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n752_), .A2(new_n764_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n319_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n728_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n778_), .A2(new_n774_), .A3(new_n771_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n775_), .A2(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n305_), .A2(G113gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n773_), .B1(new_n780_), .B2(new_n781_), .ZN(G1340gat));
  INV_X1    g581(.A(G120gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n266_), .B2(KEYINPUT60), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n772_), .B(new_n784_), .C1(KEYINPUT60), .C2(new_n783_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n775_), .A2(new_n266_), .A3(new_n779_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(new_n783_), .ZN(G1341gat));
  AOI21_X1  g586(.A(G127gat), .B1(new_n772_), .B2(new_n318_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n318_), .A2(G127gat), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT121), .Z(new_n790_));
  AOI21_X1  g589(.A(new_n788_), .B1(new_n780_), .B2(new_n790_), .ZN(G1342gat));
  AOI21_X1  g590(.A(G134gat), .B1(new_n772_), .B2(new_n347_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n635_), .A2(G134gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n780_), .B2(new_n793_), .ZN(G1343gat));
  NAND4_X1  g593(.A1(new_n769_), .A2(new_n305_), .A3(new_n564_), .A4(new_n770_), .ZN(new_n795_));
  XOR2_X1   g594(.A(KEYINPUT122), .B(G141gat), .Z(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(G1344gat));
  NAND4_X1  g596(.A1(new_n769_), .A2(new_n267_), .A3(new_n564_), .A4(new_n770_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(KEYINPUT123), .B(G148gat), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n798_), .B(new_n799_), .ZN(G1345gat));
  NAND4_X1  g599(.A1(new_n769_), .A2(new_n318_), .A3(new_n564_), .A4(new_n770_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT61), .B(G155gat), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n801_), .B(new_n802_), .ZN(G1346gat));
  NAND2_X1  g602(.A1(new_n769_), .A2(new_n564_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n804_), .A2(new_n422_), .A3(new_n602_), .ZN(new_n805_));
  INV_X1    g604(.A(G162gat), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n361_), .A2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n769_), .A2(new_n347_), .A3(new_n564_), .A4(new_n770_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n805_), .A2(new_n807_), .B1(new_n806_), .B2(new_n808_), .ZN(G1347gat));
  INV_X1    g608(.A(KEYINPUT124), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n499_), .A2(new_n590_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n563_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n778_), .A2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n306_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n810_), .B1(new_n815_), .B2(new_n428_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT124), .B(G169gat), .C1(new_n814_), .C2(new_n306_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(KEYINPUT62), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n815_), .A2(new_n464_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT62), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n810_), .B(new_n820_), .C1(new_n815_), .C2(new_n428_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n819_), .A3(new_n821_), .ZN(G1348gat));
  INV_X1    g621(.A(new_n814_), .ZN(new_n823_));
  AOI21_X1  g622(.A(G176gat), .B1(new_n823_), .B2(new_n267_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n752_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT120), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(new_n319_), .A3(new_n760_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n812_), .B1(new_n827_), .B2(new_n728_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n266_), .A2(new_n429_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n824_), .B1(new_n828_), .B2(new_n829_), .ZN(G1349gat));
  AOI21_X1  g629(.A(G183gat), .B1(new_n828_), .B2(new_n318_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n814_), .A2(new_n319_), .A3(new_n423_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT125), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(G183gat), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n769_), .A2(new_n813_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n319_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT125), .ZN(new_n837_));
  INV_X1    g636(.A(new_n832_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n833_), .A2(new_n839_), .ZN(G1350gat));
  OAI21_X1  g639(.A(G190gat), .B1(new_n814_), .B2(new_n361_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n347_), .A2(new_n424_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n814_), .B2(new_n842_), .ZN(G1351gat));
  NAND4_X1  g642(.A1(new_n769_), .A2(new_n305_), .A3(new_n564_), .A4(new_n811_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT126), .B(G197gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1352gat));
  NAND4_X1  g645(.A1(new_n769_), .A2(new_n267_), .A3(new_n564_), .A4(new_n811_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g647(.A1(new_n769_), .A2(new_n318_), .A3(new_n564_), .A4(new_n811_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n850_));
  AND2_X1   g649(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n849_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n850_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT127), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n849_), .A2(KEYINPUT127), .A3(new_n850_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n852_), .B1(new_n855_), .B2(new_n856_), .ZN(G1354gat));
  NOR3_X1   g656(.A1(new_n804_), .A2(new_n590_), .A3(new_n499_), .ZN(new_n858_));
  INV_X1    g657(.A(G218gat), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n361_), .A2(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n769_), .A2(new_n347_), .A3(new_n564_), .A4(new_n811_), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n858_), .A2(new_n860_), .B1(new_n859_), .B2(new_n861_), .ZN(G1355gat));
endmodule


