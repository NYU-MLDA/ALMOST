//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT78), .B(KEYINPUT23), .Z(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(KEYINPUT79), .A3(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT79), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT78), .B(KEYINPUT23), .ZN(new_n207_));
  INV_X1    g006(.A(new_n204_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(KEYINPUT80), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT80), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n205_), .B(new_n209_), .C1(KEYINPUT23), .C2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT25), .B(G183gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT26), .B(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n218_), .A2(KEYINPUT24), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n217_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n214_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n207_), .A2(new_n208_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n210_), .A2(new_n212_), .A3(KEYINPUT23), .ZN(new_n226_));
  INV_X1    g025(.A(G183gat), .ZN(new_n227_));
  INV_X1    g026(.A(G190gat), .ZN(new_n228_));
  AOI22_X1  g027(.A1(new_n225_), .A2(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G169gat), .ZN(new_n232_));
  INV_X1    g031(.A(G176gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n219_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n236_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n224_), .B1(new_n231_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT30), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  OAI211_X1 g039(.A(KEYINPUT30), .B(new_n224_), .C1(new_n231_), .C2(new_n237_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n240_), .A2(KEYINPUT83), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT83), .B1(new_n240_), .B2(new_n241_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT82), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G15gat), .B(G43gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G71gat), .B(G99gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n242_), .A2(new_n243_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n243_), .A2(new_n249_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n202_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n249_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n240_), .A2(new_n241_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(new_n255_), .B2(KEYINPUT83), .ZN(new_n256_));
  OAI211_X1 g055(.A(KEYINPUT84), .B(new_n251_), .C1(new_n256_), .C2(new_n242_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G127gat), .B(G134gat), .Z(new_n258_));
  XOR2_X1   g057(.A(G113gat), .B(G120gat), .Z(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  XOR2_X1   g059(.A(new_n260_), .B(KEYINPUT31), .Z(new_n261_));
  NAND3_X1  g060(.A1(new_n253_), .A2(new_n257_), .A3(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n250_), .A2(new_n252_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n261_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(KEYINPUT84), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT3), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT2), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272_));
  OR2_X1    g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n267_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n276_), .B1(new_n272_), .B2(KEYINPUT1), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(KEYINPUT1), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n273_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(new_n272_), .A2(new_n276_), .A3(KEYINPUT1), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n275_), .B(new_n269_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n274_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT86), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT86), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n274_), .A2(new_n284_), .A3(new_n281_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(KEYINPUT29), .A3(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G197gat), .B(G204gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT21), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(G197gat), .A2(G204gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G197gat), .A2(G204gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(KEYINPUT21), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n289_), .A2(KEYINPUT87), .A3(new_n292_), .A4(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(KEYINPUT87), .ZN(new_n295_));
  INV_X1    g094(.A(new_n287_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(KEYINPUT21), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT88), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n294_), .A2(KEYINPUT88), .A3(new_n297_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(G228gat), .A2(G233gat), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n286_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n282_), .A2(KEYINPUT29), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n298_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n303_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G78gat), .B(G106gat), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT89), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n283_), .A2(new_n285_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G22gat), .B(G50gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n315_), .B(KEYINPUT28), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n314_), .B(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n309_), .A2(new_n310_), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n286_), .A2(new_n304_), .B1(new_n307_), .B2(new_n303_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n310_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  OAI22_X1  g121(.A1(new_n311_), .A2(new_n318_), .B1(new_n319_), .B2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n314_), .B(new_n316_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n309_), .A2(new_n310_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n321_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(KEYINPUT89), .A4(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n266_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n283_), .A2(new_n285_), .A3(new_n260_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n282_), .A2(new_n260_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(KEYINPUT4), .A3(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT93), .B(KEYINPUT4), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n283_), .A2(new_n285_), .A3(new_n260_), .A4(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n330_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT0), .ZN(new_n338_));
  INV_X1    g137(.A(G57gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G85gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n330_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n345_));
  OR3_X1    g144(.A1(new_n336_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n343_), .B1(new_n336_), .B2(new_n345_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n227_), .A2(new_n228_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n235_), .B1(new_n214_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n225_), .A2(new_n226_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(new_n222_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n298_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT20), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT95), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT19), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n302_), .B(new_n224_), .C1(new_n231_), .C2(new_n237_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n356_), .A2(new_n357_), .A3(new_n360_), .A4(new_n361_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n361_), .A2(KEYINPUT20), .A3(new_n360_), .A4(new_n354_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT95), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n214_), .A2(new_n349_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n353_), .B1(new_n365_), .B2(new_n236_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n298_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n301_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT88), .B1(new_n294_), .B2(new_n297_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n238_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n368_), .A2(new_n372_), .A3(KEYINPUT20), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n359_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n362_), .A2(new_n364_), .A3(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G64gat), .B(G92gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(G8gat), .B(G36gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n375_), .A2(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n238_), .A2(new_n371_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n359_), .B1(new_n355_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n360_), .A2(KEYINPUT20), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(new_n238_), .B2(new_n371_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT90), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n388_));
  NOR4_X1   g187(.A1(new_n350_), .A2(KEYINPUT90), .A3(new_n353_), .A4(new_n298_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n386_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n384_), .A2(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n348_), .B(new_n382_), .C1(new_n381_), .C2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT92), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n384_), .A2(new_n390_), .A3(new_n380_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n380_), .B1(new_n384_), .B2(new_n390_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n380_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n391_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n384_), .A2(new_n390_), .A3(new_n380_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(KEYINPUT92), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(KEYINPUT33), .B(new_n343_), .C1(new_n336_), .C2(new_n345_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n333_), .A2(new_n330_), .A3(new_n335_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n331_), .A2(new_n344_), .A3(new_n332_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n342_), .A3(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT94), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT33), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n347_), .B2(new_n408_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n347_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n401_), .B(new_n406_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n329_), .B1(new_n392_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n375_), .A2(new_n397_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT96), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n394_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n399_), .B2(KEYINPUT96), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n413_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n346_), .A2(new_n347_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n416_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n328_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n266_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n262_), .A2(new_n328_), .A3(new_n265_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n412_), .A2(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(KEYINPUT10), .B(G99gat), .Z(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT64), .B(G106gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G85gat), .B(G92gat), .Z(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT9), .ZN(new_n431_));
  INV_X1    g230(.A(G92gat), .ZN(new_n432_));
  OR3_X1    g231(.A1(new_n341_), .A2(new_n432_), .A3(KEYINPUT9), .ZN(new_n433_));
  AND3_X1   g232(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n429_), .A2(new_n431_), .A3(new_n433_), .A4(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(G99gat), .ZN(new_n438_));
  INV_X1    g237(.A(G106gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(KEYINPUT65), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT7), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT7), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n442_), .A2(new_n438_), .A3(new_n439_), .A4(KEYINPUT65), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n436_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT8), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n430_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n445_), .B1(new_n444_), .B2(new_n430_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n437_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G57gat), .B(G64gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT11), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT11), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n339_), .A2(G64gat), .ZN(new_n452_));
  INV_X1    g251(.A(G64gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(G57gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n451_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G71gat), .B(G78gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n450_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n449_), .A2(new_n456_), .A3(KEYINPUT11), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n448_), .A2(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n437_), .B(new_n460_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(KEYINPUT66), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G230gat), .A2(G233gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n464_), .B(new_n466_), .C1(KEYINPUT66), .C2(new_n462_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n465_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT67), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT67), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n463_), .A2(new_n470_), .A3(new_n465_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(new_n448_), .B2(new_n461_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n448_), .A2(new_n472_), .A3(new_n461_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n469_), .B(new_n471_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G120gat), .B(G148gat), .Z(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(G204gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT5), .B(G176gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  NAND3_X1  g278(.A1(new_n467_), .A2(new_n475_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n479_), .B1(new_n467_), .B2(new_n475_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT68), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n467_), .A2(new_n475_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n479_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT68), .B1(new_n487_), .B2(new_n480_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n489_), .A2(KEYINPUT13), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(KEYINPUT13), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G229gat), .A2(G233gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G15gat), .B(G22gat), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(KEYINPUT71), .A2(G1gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(KEYINPUT71), .A2(G1gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(G8gat), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n499_), .A2(KEYINPUT72), .A3(KEYINPUT14), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT72), .B1(new_n499_), .B2(KEYINPUT14), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n496_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G1gat), .B(G8gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G29gat), .B(G36gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G43gat), .B(G50gat), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n507_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n503_), .B(new_n496_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n505_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n511_), .B1(new_n505_), .B2(new_n512_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n494_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n499_), .A2(KEYINPUT14), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT72), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n499_), .A2(KEYINPUT72), .A3(KEYINPUT14), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n503_), .B1(new_n520_), .B2(new_n496_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n512_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n510_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n508_), .A2(KEYINPUT15), .A3(new_n509_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT15), .B1(new_n508_), .B2(new_n509_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(new_n512_), .A3(new_n505_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n523_), .A2(new_n527_), .A3(new_n493_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G169gat), .B(G197gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT75), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n530_), .B(new_n531_), .Z(new_n532_));
  NAND3_X1  g331(.A1(new_n515_), .A2(new_n528_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT76), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT76), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n515_), .A2(new_n528_), .A3(new_n535_), .A4(new_n532_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n515_), .A2(new_n528_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n532_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT77), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n426_), .A2(new_n492_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n505_), .A2(new_n512_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G231gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(new_n461_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n547_), .A2(KEYINPUT73), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G127gat), .B(G155gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT16), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(G183gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(G211gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT17), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT74), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n548_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n547_), .A2(KEYINPUT73), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n552_), .B(KEYINPUT17), .Z(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n547_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n563_), .B(KEYINPUT36), .Z(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n448_), .A2(new_n526_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT34), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n571_), .B1(new_n448_), .B2(new_n511_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n566_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT69), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n574_), .B(new_n571_), .C1(new_n448_), .C2(new_n511_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n569_), .A2(new_n570_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n575_), .B(new_n576_), .C1(new_n566_), .C2(new_n572_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n565_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n563_), .A2(KEYINPUT36), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n578_), .A2(new_n579_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n580_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT70), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n584_), .A3(KEYINPUT37), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n578_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n584_), .B(new_n586_), .C1(new_n582_), .C2(new_n565_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n585_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n560_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n543_), .A2(new_n591_), .ZN(new_n592_));
  NOR4_X1   g391(.A1(new_n592_), .A2(new_n419_), .A3(new_n498_), .A4(new_n497_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n583_), .B(KEYINPUT98), .Z(new_n596_));
  NOR2_X1   g395(.A1(new_n426_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n541_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n492_), .A2(new_n560_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(G1gat), .B1(new_n600_), .B2(new_n419_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n601_), .ZN(G1324gat));
  NAND2_X1  g401(.A1(new_n418_), .A2(new_n420_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G8gat), .B1(new_n600_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT39), .ZN(new_n606_));
  OR3_X1    g405(.A1(new_n592_), .A2(G8gat), .A3(new_n604_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT40), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(G1325gat));
  NOR3_X1   g409(.A1(new_n592_), .A2(G15gat), .A3(new_n266_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT100), .ZN(new_n612_));
  INV_X1    g411(.A(new_n266_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n597_), .A2(new_n613_), .A3(new_n599_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(G15gat), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(KEYINPUT99), .A3(G15gat), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT41), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT41), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n617_), .A2(new_n621_), .A3(new_n618_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n612_), .A2(new_n620_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT101), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n612_), .A2(new_n620_), .A3(new_n625_), .A4(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(G1326gat));
  OAI21_X1  g426(.A(G22gat), .B1(new_n600_), .B2(new_n328_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT42), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n328_), .A2(G22gat), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n592_), .B2(new_n630_), .ZN(G1327gat));
  NAND2_X1  g430(.A1(new_n560_), .A2(new_n583_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT102), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n543_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(G29gat), .B1(new_n635_), .B2(new_n348_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n590_), .B1(new_n412_), .B2(new_n425_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT43), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n394_), .A2(new_n395_), .A3(new_n393_), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT92), .B1(new_n398_), .B2(new_n399_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n406_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n410_), .A2(new_n409_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n392_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n422_), .B1(new_n265_), .B2(new_n262_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n262_), .A2(new_n328_), .A3(new_n265_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n328_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n645_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n590_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n638_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n560_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n492_), .A2(new_n654_), .A3(new_n598_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT44), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  INV_X1    g456(.A(new_n492_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n560_), .A3(new_n541_), .ZN(new_n659_));
  AOI211_X1 g458(.A(new_n657_), .B(new_n659_), .C1(new_n638_), .C2(new_n652_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n656_), .A2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n348_), .A2(G29gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n636_), .B1(new_n661_), .B2(new_n662_), .ZN(G1328gat));
  AOI21_X1  g462(.A(new_n651_), .B1(new_n650_), .B2(new_n590_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n590_), .ZN(new_n665_));
  AOI211_X1 g464(.A(KEYINPUT43), .B(new_n665_), .C1(new_n645_), .C2(new_n649_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n655_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n657_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n653_), .A2(KEYINPUT44), .A3(new_n655_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n603_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n668_), .A2(new_n669_), .A3(KEYINPUT103), .A4(new_n603_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(G36gat), .A3(new_n673_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n634_), .A2(G36gat), .A3(new_n604_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT45), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT46), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n674_), .A2(KEYINPUT46), .A3(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1329gat));
  INV_X1    g481(.A(G43gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n683_), .B1(new_n634_), .B2(new_n266_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n266_), .A2(new_n683_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT104), .B1(new_n661_), .B2(new_n685_), .ZN(new_n686_));
  AND4_X1   g485(.A1(KEYINPUT104), .A2(new_n668_), .A3(new_n669_), .A4(new_n685_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n684_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n689_), .B(new_n684_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1330gat));
  AOI21_X1  g492(.A(G50gat), .B1(new_n635_), .B2(new_n422_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n422_), .A2(G50gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n661_), .B2(new_n695_), .ZN(G1331gat));
  AND3_X1   g495(.A1(new_n492_), .A2(new_n654_), .A3(new_n542_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n597_), .A2(new_n697_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n698_), .A2(new_n339_), .A3(new_n419_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT108), .Z(new_n700_));
  NAND2_X1  g499(.A1(new_n650_), .A2(new_n598_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT106), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(KEYINPUT106), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n658_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n591_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n705_), .A2(KEYINPUT107), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(KEYINPUT107), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n348_), .A3(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n700_), .B1(new_n708_), .B2(new_n339_), .ZN(G1332gat));
  OAI21_X1  g508(.A(G64gat), .B1(new_n698_), .B2(new_n604_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT48), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n706_), .A2(new_n707_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n603_), .A2(new_n453_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n711_), .B1(new_n712_), .B2(new_n713_), .ZN(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n698_), .B2(new_n266_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT49), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n266_), .A2(G71gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT109), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n712_), .B2(new_n718_), .ZN(G1334gat));
  OAI21_X1  g518(.A(G78gat), .B1(new_n698_), .B2(new_n328_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT50), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n328_), .A2(G78gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n712_), .B2(new_n722_), .ZN(G1335gat));
  NOR3_X1   g522(.A1(new_n658_), .A2(new_n654_), .A3(new_n541_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n653_), .A2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G85gat), .B1(new_n725_), .B2(new_n419_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n704_), .A2(new_n633_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n348_), .A2(new_n341_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n726_), .B1(new_n727_), .B2(new_n728_), .ZN(G1336gat));
  OAI21_X1  g528(.A(G92gat), .B1(new_n725_), .B2(new_n604_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n603_), .A2(new_n432_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n727_), .B2(new_n731_), .ZN(G1337gat));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  OAI21_X1  g532(.A(G99gat), .B1(new_n725_), .B2(new_n266_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n613_), .A2(new_n427_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n733_), .B(new_n734_), .C1(new_n727_), .C2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g536(.A1(new_n653_), .A2(new_n422_), .A3(new_n724_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(G106gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G106gat), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n422_), .A2(new_n428_), .ZN(new_n742_));
  OAI22_X1  g541(.A1(new_n740_), .A2(new_n741_), .B1(new_n727_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g543(.A1(new_n604_), .A2(new_n348_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n745_), .A2(new_n424_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n475_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n473_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n448_), .A2(new_n472_), .A3(new_n461_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n752_), .A2(KEYINPUT55), .A3(new_n471_), .A4(new_n469_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n463_), .B1(new_n474_), .B2(new_n473_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n466_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n749_), .A2(new_n753_), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n486_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT111), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n756_), .A2(KEYINPUT111), .A3(new_n758_), .A4(new_n486_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n481_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n760_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n505_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n494_), .B1(new_n523_), .B2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n766_), .B2(new_n532_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n493_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(KEYINPUT112), .A3(new_n539_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n523_), .A2(new_n527_), .A3(new_n494_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n537_), .A2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n484_), .B2(new_n488_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n763_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n583_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(KEYINPUT57), .A3(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n583_), .B1(new_n763_), .B2(new_n773_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT113), .B1(new_n779_), .B2(KEYINPUT57), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n757_), .A2(KEYINPUT56), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n537_), .A2(new_n480_), .A3(new_n771_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n756_), .A2(new_n758_), .A3(new_n486_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n782_), .A2(new_n783_), .A3(KEYINPUT58), .A4(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n590_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n758_), .B1(new_n756_), .B2(new_n486_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n537_), .A2(new_n480_), .A3(new_n771_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT58), .B1(new_n789_), .B2(new_n784_), .ZN(new_n790_));
  OAI22_X1  g589(.A1(new_n779_), .A2(KEYINPUT57), .B1(new_n786_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT114), .B1(new_n781_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n776_), .A2(new_n777_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n779_), .A2(KEYINPUT113), .A3(KEYINPUT57), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n791_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n792_), .A2(new_n560_), .A3(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n591_), .A2(new_n490_), .A3(new_n491_), .A4(new_n542_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT54), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n747_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(G113gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n541_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT59), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n560_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n793_), .A2(new_n794_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n791_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n806_), .A2(new_n796_), .A3(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n800_), .B1(new_n805_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n804_), .B1(new_n809_), .B2(new_n746_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n800_), .B1(new_n654_), .B2(new_n795_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n747_), .A2(KEYINPUT115), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n747_), .A2(KEYINPUT115), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n812_), .A2(new_n813_), .A3(KEYINPUT59), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n811_), .A2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT116), .B1(new_n810_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n811_), .A2(new_n814_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n817_), .B(new_n818_), .C1(new_n801_), .C2(new_n804_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n542_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n803_), .B1(new_n820_), .B2(new_n802_), .ZN(G1340gat));
  XOR2_X1   g620(.A(KEYINPUT117), .B(G120gat), .Z(new_n822_));
  NOR2_X1   g621(.A1(new_n822_), .A2(KEYINPUT60), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n658_), .B2(KEYINPUT60), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n801_), .B(new_n826_), .C1(new_n825_), .C2(new_n824_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n810_), .A2(new_n815_), .A3(new_n658_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n828_), .B2(new_n822_), .ZN(G1341gat));
  AOI21_X1  g628(.A(G127gat), .B1(new_n801_), .B2(new_n654_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n816_), .A2(new_n819_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n654_), .A2(G127gat), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT119), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n830_), .B1(new_n831_), .B2(new_n833_), .ZN(G1342gat));
  INV_X1    g633(.A(G134gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n801_), .A2(new_n835_), .A3(new_n596_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n665_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n835_), .ZN(G1343gat));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n745_), .A2(new_n423_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n809_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n839_), .B1(new_n809_), .B2(new_n840_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n541_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G141gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n809_), .A2(new_n840_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT120), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n841_), .ZN(new_n848_));
  INV_X1    g647(.A(G141gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n541_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n845_), .A2(new_n850_), .ZN(G1344gat));
  XNOR2_X1  g650(.A(KEYINPUT121), .B(G148gat), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT122), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n848_), .B2(new_n492_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n853_), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n658_), .B(new_n855_), .C1(new_n847_), .C2(new_n841_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1345gat));
  XNOR2_X1  g656(.A(KEYINPUT61), .B(G155gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT123), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n848_), .B2(new_n654_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n859_), .ZN(new_n861_));
  AOI211_X1 g660(.A(new_n560_), .B(new_n861_), .C1(new_n847_), .C2(new_n841_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1346gat));
  NAND2_X1  g662(.A1(new_n848_), .A2(new_n596_), .ZN(new_n864_));
  INV_X1    g663(.A(G162gat), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n590_), .A2(G162gat), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(KEYINPUT124), .Z(new_n867_));
  AOI22_X1  g666(.A1(new_n864_), .A2(new_n865_), .B1(new_n848_), .B2(new_n867_), .ZN(G1347gat));
  NOR3_X1   g667(.A1(new_n604_), .A2(new_n348_), .A3(new_n424_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n811_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G169gat), .B1(new_n870_), .B2(new_n598_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT62), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n870_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n232_), .A3(new_n541_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n872_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(new_n875_), .A3(new_n876_), .ZN(G1348gat));
  AOI21_X1  g676(.A(G176gat), .B1(new_n874_), .B2(new_n492_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n422_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n613_), .A2(new_n419_), .A3(new_n603_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n658_), .A2(new_n233_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n878_), .B1(new_n879_), .B2(new_n881_), .ZN(G1349gat));
  NOR2_X1   g681(.A1(new_n880_), .A2(new_n560_), .ZN(new_n883_));
  AOI21_X1  g682(.A(G183gat), .B1(new_n879_), .B2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n560_), .A2(new_n215_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n874_), .B2(new_n885_), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n870_), .B2(new_n665_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n596_), .A2(new_n216_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n870_), .B2(new_n888_), .ZN(G1351gat));
  NOR2_X1   g688(.A1(new_n423_), .A2(new_n348_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n890_), .A2(KEYINPUT125), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(KEYINPUT125), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n604_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n809_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n541_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g696(.A1(new_n894_), .A2(new_n658_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT126), .B(G204gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1353gat));
  INV_X1    g699(.A(KEYINPUT127), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n894_), .A2(new_n560_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n903_));
  INV_X1    g702(.A(G211gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n901_), .B1(new_n902_), .B2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  OAI211_X1 g706(.A(KEYINPUT127), .B(new_n907_), .C1(new_n894_), .C2(new_n560_), .ZN(new_n908_));
  XOR2_X1   g707(.A(KEYINPUT63), .B(G211gat), .Z(new_n909_));
  AOI22_X1  g708(.A1(new_n906_), .A2(new_n908_), .B1(new_n902_), .B2(new_n909_), .ZN(G1354gat));
  OAI21_X1  g709(.A(G218gat), .B1(new_n894_), .B2(new_n665_), .ZN(new_n911_));
  INV_X1    g710(.A(G218gat), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n596_), .A2(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n911_), .B1(new_n894_), .B2(new_n913_), .ZN(G1355gat));
endmodule


