//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n957_, new_n958_, new_n959_,
    new_n961_, new_n962_, new_n963_, new_n965_, new_n966_, new_n967_,
    new_n969_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_, new_n978_, new_n979_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT72), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT36), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT15), .ZN(new_n207_));
  INV_X1    g006(.A(G36gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G29gat), .ZN(new_n209_));
  INV_X1    g008(.A(G29gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G36gat), .ZN(new_n211_));
  INV_X1    g010(.A(G43gat), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n209_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n212_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT67), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n210_), .A2(G36gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n208_), .A2(G29gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(G43gat), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n209_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n215_), .A2(G50gat), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(G50gat), .B1(new_n215_), .B2(new_n221_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n207_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT6), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n230_));
  INV_X1    g029(.A(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G85gat), .A2(G92gat), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n234_), .A2(KEYINPUT9), .ZN(new_n235_));
  INV_X1    g034(.A(G85gat), .ZN(new_n236_));
  INV_X1    g035(.A(G92gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(KEYINPUT9), .A3(new_n234_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n229_), .A2(new_n233_), .A3(new_n235_), .A4(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n241_));
  INV_X1    g040(.A(G99gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(new_n231_), .ZN(new_n243_));
  OAI22_X1  g042(.A1(KEYINPUT64), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n243_), .A2(new_n227_), .A3(new_n228_), .A4(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT8), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n238_), .A2(new_n234_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n246_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n240_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G50gat), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT67), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n219_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n215_), .A2(new_n221_), .A3(G50gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(KEYINPUT15), .A3(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n224_), .A2(new_n251_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n255_), .A2(new_n256_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n240_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n245_), .A2(new_n247_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT8), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n262_), .B1(new_n264_), .B2(new_n248_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n260_), .B1(new_n261_), .B2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n258_), .A2(new_n259_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G232gat), .A2(G233gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n268_), .B(KEYINPUT34), .Z(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n258_), .A2(new_n259_), .A3(new_n266_), .A4(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT35), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n258_), .A2(new_n274_), .A3(new_n266_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n270_), .A2(KEYINPUT35), .A3(new_n272_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n206_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n278_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n206_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n280_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(KEYINPUT69), .B(KEYINPUT36), .Z(new_n285_));
  NOR2_X1   g084(.A1(new_n204_), .A2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n286_), .B(KEYINPUT70), .Z(new_n287_));
  NAND3_X1  g086(.A1(new_n277_), .A2(new_n278_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT37), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n284_), .A2(new_n289_), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n270_), .A2(KEYINPUT35), .A3(new_n272_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n275_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n283_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT74), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n295_), .B(new_n283_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n296_), .A3(new_n288_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT37), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n281_), .A2(new_n290_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G57gat), .B(G64gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(KEYINPUT11), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G71gat), .B(G78gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(KEYINPUT11), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n300_), .A2(new_n302_), .A3(KEYINPUT11), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G231gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G1gat), .B(G8gat), .Z(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G15gat), .B(G22gat), .ZN(new_n312_));
  INV_X1    g111(.A(G1gat), .ZN(new_n313_));
  INV_X1    g112(.A(G8gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT14), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT75), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n316_), .A2(KEYINPUT75), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n311_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n319_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(new_n310_), .A3(new_n317_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n309_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n325_), .A2(KEYINPUT77), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(KEYINPUT77), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G127gat), .B(G155gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G183gat), .B(G211gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n332_), .B(KEYINPUT17), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT78), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n326_), .A2(new_n327_), .A3(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n325_), .A2(KEYINPUT17), .A3(new_n332_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n299_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n251_), .A2(new_n306_), .A3(new_n305_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT12), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(KEYINPUT65), .A3(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT65), .B1(new_n265_), .B2(new_n307_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT12), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G230gat), .A2(G233gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n265_), .A2(new_n307_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n343_), .A2(new_n345_), .A3(new_n346_), .A4(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT66), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n344_), .A2(KEYINPUT12), .B1(new_n265_), .B2(new_n307_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n351_), .A2(KEYINPUT66), .A3(new_n346_), .A4(new_n343_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n341_), .A2(new_n347_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(G230gat), .A3(G233gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G120gat), .B(G148gat), .ZN(new_n356_));
  INV_X1    g155(.A(G204gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT5), .B(G176gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n355_), .B(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT13), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n362_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G229gat), .A2(G233gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n224_), .A2(new_n323_), .A3(new_n257_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n323_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n255_), .A2(KEYINPUT79), .A3(new_n256_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT79), .B1(new_n255_), .B2(new_n256_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n368_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n372_), .A2(KEYINPUT80), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n374_));
  INV_X1    g173(.A(new_n371_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n369_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n374_), .B1(new_n376_), .B2(new_n368_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n366_), .B(new_n367_), .C1(new_n373_), .C2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n376_), .A2(new_n368_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n372_), .A2(KEYINPUT80), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(new_n374_), .A3(new_n368_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n378_), .B1(new_n382_), .B2(new_n366_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G113gat), .B(G141gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G169gat), .ZN(new_n385_));
  INV_X1    g184(.A(G197gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n378_), .B(new_n387_), .C1(new_n382_), .C2(new_n366_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(KEYINPUT81), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n383_), .A2(new_n392_), .A3(new_n388_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n365_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G225gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n398_));
  INV_X1    g197(.A(G134gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(G127gat), .ZN(new_n400_));
  INV_X1    g199(.A(G127gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(G134gat), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n400_), .A2(new_n402_), .A3(KEYINPUT86), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT86), .B1(new_n400_), .B2(new_n402_), .ZN(new_n404_));
  OAI21_X1  g203(.A(G113gat), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT86), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n401_), .A2(G134gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n399_), .A2(G127gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n406_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G113gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n400_), .A2(new_n402_), .A3(KEYINPUT86), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n405_), .A2(G120gat), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(G120gat), .B1(new_n405_), .B2(new_n412_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n398_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(G155gat), .ZN(new_n416_));
  INV_X1    g215(.A(G162gat), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT1), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT1), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(G155gat), .A3(G162gat), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .A4(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G141gat), .A2(G148gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT87), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT87), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(G141gat), .A3(G148gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(G141gat), .A2(G148gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n424_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT2), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n429_), .A2(new_n434_), .B1(KEYINPUT3), .B2(new_n431_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT91), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT90), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT3), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(new_n430_), .B2(KEYINPUT89), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n441_), .A2(G141gat), .A3(G148gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n438_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n430_), .A2(KEYINPUT89), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n441_), .B1(G141gat), .B2(G148gat), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n444_), .A2(KEYINPUT90), .A3(new_n445_), .A4(new_n439_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n435_), .A2(new_n437_), .A3(new_n443_), .A4(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n420_), .A2(new_n421_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n448_), .B1(G155gat), .B2(G162gat), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n433_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n415_), .A2(KEYINPUT99), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT99), .ZN(new_n452_));
  INV_X1    g251(.A(G120gat), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n403_), .A2(new_n404_), .A3(G113gat), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n410_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n453_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n405_), .A2(new_n412_), .A3(G120gat), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT4), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n429_), .A2(new_n434_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n431_), .A2(KEYINPUT3), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n437_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n443_), .A2(new_n446_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n449_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n432_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n452_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n397_), .B1(new_n451_), .B2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n413_), .A2(new_n414_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT98), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n450_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n463_), .A2(new_n468_), .A3(new_n432_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n456_), .A2(new_n457_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n469_), .A2(new_n472_), .A3(KEYINPUT4), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT100), .B1(new_n466_), .B2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT99), .B1(new_n415_), .B2(new_n450_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n458_), .A2(new_n452_), .A3(new_n464_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n469_), .A2(new_n472_), .A3(KEYINPUT4), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT100), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .A4(new_n397_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n469_), .A2(new_n472_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(new_n397_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n474_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G1gat), .B(G29gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT102), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G57gat), .B(G85gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n486_), .B(new_n489_), .Z(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n484_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT103), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n474_), .A2(new_n480_), .A3(new_n490_), .A4(new_n483_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n484_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(KEYINPUT103), .A3(new_n490_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G226gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT19), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT25), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n501_), .A2(G183gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(G183gat), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G190gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT26), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT26), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(G190gat), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(G169gat), .A2(G176gat), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT24), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(G169gat), .A2(G176gat), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n514_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n510_), .A2(new_n513_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G183gat), .A2(G190gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT23), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n519_), .B1(new_n520_), .B2(new_n518_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT22), .B(G169gat), .ZN(new_n522_));
  INV_X1    g321(.A(G176gat), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n514_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n525_));
  NOR2_X1   g324(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n518_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT23), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n528_), .A2(KEYINPUT84), .A3(G183gat), .A4(G190gat), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT84), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n530_), .B1(new_n518_), .B2(KEYINPUT23), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(G183gat), .A2(G190gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n517_), .A2(new_n521_), .B1(new_n524_), .B2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G211gat), .B(G218gat), .Z(new_n537_));
  NAND2_X1  g336(.A1(new_n386_), .A2(G204gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n357_), .A2(G197gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n537_), .A2(KEYINPUT21), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT95), .B1(new_n540_), .B2(KEYINPUT21), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT21), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n538_), .A2(new_n539_), .A3(new_n544_), .A4(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n357_), .B2(G197gat), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n386_), .A2(KEYINPUT94), .A3(G204gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n539_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n537_), .B1(new_n551_), .B2(KEYINPUT21), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n542_), .B1(new_n547_), .B2(new_n552_), .ZN(new_n553_));
  OR3_X1    g352(.A1(new_n536_), .A2(KEYINPUT96), .A3(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT96), .B1(new_n536_), .B2(new_n553_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n532_), .A2(new_n513_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT85), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n532_), .A2(KEYINPUT85), .A3(new_n513_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT82), .B1(new_n501_), .B2(G183gat), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n561_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT82), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n563_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n515_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n559_), .A2(new_n560_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n521_), .A2(new_n534_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n524_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n553_), .A3(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n569_), .A2(KEYINPUT20), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n500_), .B1(new_n556_), .B2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(KEYINPUT97), .B(KEYINPUT18), .Z(new_n572_));
  XNOR2_X1  g371(.A(G8gat), .B(G36gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G64gat), .B(G92gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n577_), .A2(KEYINPUT32), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n536_), .A2(new_n553_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT20), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n553_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n580_), .A2(new_n581_), .A3(new_n499_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n571_), .A2(new_n578_), .A3(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n556_), .A2(new_n500_), .A3(new_n570_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n499_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n583_), .B1(new_n578_), .B2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n495_), .A2(new_n497_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n582_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n556_), .A2(new_n570_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n577_), .B(new_n589_), .C1(new_n590_), .C2(new_n500_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n477_), .A2(new_n478_), .A3(new_n396_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n592_), .B(new_n491_), .C1(new_n481_), .C2(new_n396_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n576_), .B1(new_n571_), .B2(new_n582_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n591_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n494_), .A2(KEYINPUT33), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n494_), .A2(KEYINPUT33), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n588_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n560_), .A2(new_n565_), .ZN(new_n600_));
  AOI21_X1  g399(.A(KEYINPUT85), .B1(new_n532_), .B2(new_n513_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n568_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT30), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  OAI211_X1 g403(.A(KEYINPUT30), .B(new_n568_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G15gat), .B(G43gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G71gat), .B(G99gat), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n610_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n604_), .A2(new_n605_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n606_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n612_), .B1(new_n615_), .B2(new_n607_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n467_), .A2(KEYINPUT31), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT31), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n471_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G227gat), .A2(G233gat), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n617_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n620_), .B1(new_n617_), .B2(new_n619_), .ZN(new_n622_));
  OAI22_X1  g421(.A1(new_n611_), .A2(new_n616_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n610_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n621_), .A2(new_n622_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n615_), .A2(new_n612_), .A3(new_n607_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n623_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n553_), .B1(new_n464_), .B2(KEYINPUT29), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT93), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n547_), .A2(new_n552_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n633_), .B2(new_n541_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G228gat), .A2(G233gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G78gat), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(G78gat), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n638_), .B(new_n635_), .C1(new_n553_), .C2(new_n632_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n637_), .A2(G106gat), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(G106gat), .B1(new_n637_), .B2(new_n639_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n631_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n637_), .A2(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n231_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n637_), .A2(G106gat), .A3(new_n639_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n630_), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT92), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n642_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n464_), .A2(KEYINPUT29), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G22gat), .B(G50gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT28), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n649_), .B(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n648_), .A2(new_n653_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n642_), .A2(new_n646_), .A3(new_n652_), .A4(new_n647_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n629_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n599_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n640_), .A2(new_n641_), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT92), .B1(new_n660_), .B2(new_n630_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n652_), .B1(new_n661_), .B2(new_n642_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n655_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n628_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n654_), .A2(new_n627_), .A3(new_n623_), .A4(new_n655_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n577_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n668_), .A2(KEYINPUT27), .A3(new_n591_), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT27), .B1(new_n591_), .B2(new_n594_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n495_), .A2(new_n497_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n666_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n659_), .A2(new_n673_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n340_), .A2(new_n395_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n672_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(new_n313_), .A3(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT38), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n297_), .B(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(new_n337_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n395_), .A3(new_n674_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G1gat), .B1(new_n682_), .B2(new_n672_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n678_), .A2(new_n683_), .ZN(G1324gat));
  INV_X1    g483(.A(new_n671_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n675_), .A2(new_n314_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT39), .ZN(new_n687_));
  INV_X1    g486(.A(new_n682_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n685_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n687_), .B1(new_n689_), .B2(G8gat), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n687_), .B(G8gat), .C1(new_n682_), .C2(new_n671_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n686_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT105), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n695_), .B(new_n686_), .C1(new_n690_), .C2(new_n692_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n694_), .A2(KEYINPUT40), .A3(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT40), .B1(new_n694_), .B2(new_n696_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1325gat));
  OAI21_X1  g498(.A(G15gat), .B1(new_n682_), .B2(new_n629_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT41), .Z(new_n701_));
  INV_X1    g500(.A(G15gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n675_), .A2(new_n702_), .A3(new_n628_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT106), .ZN(G1326gat));
  OAI21_X1  g504(.A(G22gat), .B1(new_n682_), .B2(new_n656_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT42), .ZN(new_n707_));
  INV_X1    g506(.A(G22gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n656_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n675_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(G1327gat));
  XNOR2_X1  g510(.A(new_n297_), .B(KEYINPUT104), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n659_), .B2(new_n673_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n365_), .A2(new_n394_), .A3(new_n338_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G29gat), .B1(new_n716_), .B2(new_n676_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718_));
  INV_X1    g517(.A(new_n714_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n288_), .B1(new_n279_), .B2(new_n295_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n296_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n298_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n293_), .A2(KEYINPUT73), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n281_), .A2(new_n723_), .A3(KEYINPUT37), .A4(new_n288_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n666_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n657_), .B1(new_n588_), .B2(new_n598_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n725_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n725_), .B2(KEYINPUT107), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  OAI221_X1 g530(.A(new_n725_), .B1(KEYINPUT107), .B2(new_n729_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n719_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n718_), .B1(new_n733_), .B2(KEYINPUT108), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735_));
  AOI211_X1 g534(.A(new_n735_), .B(new_n719_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT109), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n299_), .B1(new_n659_), .B2(new_n673_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT43), .B1(new_n299_), .B2(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n728_), .A2(new_n730_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n714_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n735_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n733_), .A2(KEYINPUT108), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n744_), .A2(new_n745_), .A3(new_n718_), .A4(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n737_), .A2(new_n747_), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n210_), .B(new_n672_), .C1(new_n733_), .C2(KEYINPUT44), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n717_), .B1(new_n748_), .B2(new_n749_), .ZN(G1328gat));
  INV_X1    g549(.A(KEYINPUT46), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n733_), .A2(KEYINPUT44), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n685_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n208_), .B1(new_n748_), .B2(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n671_), .A2(G36gat), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OR3_X1    g556(.A1(new_n715_), .A2(KEYINPUT110), .A3(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT110), .B1(new_n715_), .B2(new_n757_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n760_), .B(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n751_), .B1(new_n755_), .B2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n760_), .B(KEYINPUT45), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n753_), .B1(new_n737_), .B2(new_n747_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n764_), .B(KEYINPUT46), .C1(new_n765_), .C2(new_n208_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n763_), .A2(new_n766_), .ZN(G1329gat));
  NAND3_X1  g566(.A1(new_n752_), .A2(G43gat), .A3(new_n628_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n737_), .B2(new_n747_), .ZN(new_n769_));
  XOR2_X1   g568(.A(KEYINPUT111), .B(G43gat), .Z(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n716_), .B2(new_n628_), .ZN(new_n771_));
  OR3_X1    g570(.A1(new_n769_), .A2(KEYINPUT47), .A3(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT47), .B1(new_n769_), .B2(new_n771_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1330gat));
  AOI21_X1  g573(.A(G50gat), .B1(new_n716_), .B2(new_n709_), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n252_), .B(new_n656_), .C1(new_n733_), .C2(KEYINPUT44), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n748_), .B2(new_n776_), .ZN(G1331gat));
  INV_X1    g576(.A(new_n365_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n394_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(new_n340_), .A3(new_n674_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT112), .Z(new_n782_));
  INV_X1    g581(.A(G57gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n676_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n681_), .A2(new_n780_), .A3(new_n674_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G57gat), .B1(new_n785_), .B2(new_n672_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1332gat));
  INV_X1    g586(.A(G64gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n782_), .A2(new_n788_), .A3(new_n685_), .ZN(new_n789_));
  OAI21_X1  g588(.A(G64gat), .B1(new_n785_), .B2(new_n671_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT48), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1333gat));
  INV_X1    g591(.A(G71gat), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n782_), .A2(new_n793_), .A3(new_n628_), .ZN(new_n794_));
  OAI21_X1  g593(.A(G71gat), .B1(new_n785_), .B2(new_n629_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT49), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1334gat));
  NAND3_X1  g596(.A1(new_n782_), .A2(new_n638_), .A3(new_n709_), .ZN(new_n798_));
  OAI21_X1  g597(.A(G78gat), .B1(new_n785_), .B2(new_n656_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT50), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1335gat));
  NAND3_X1  g600(.A1(new_n365_), .A2(new_n394_), .A3(new_n337_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n713_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n236_), .A3(new_n676_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n802_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n807_), .A2(new_n676_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n806_), .B1(new_n808_), .B2(new_n236_), .ZN(G1336gat));
  AND2_X1   g608(.A1(new_n807_), .A2(new_n685_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n685_), .A2(new_n237_), .ZN(new_n811_));
  OAI22_X1  g610(.A1(new_n810_), .A2(new_n237_), .B1(new_n804_), .B2(new_n811_), .ZN(new_n812_));
  XOR2_X1   g611(.A(new_n812_), .B(KEYINPUT113), .Z(G1337gat));
  AOI21_X1  g612(.A(new_n242_), .B1(new_n807_), .B2(new_n628_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n628_), .A2(new_n230_), .A3(new_n232_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n805_), .B2(new_n815_), .ZN(new_n816_));
  XOR2_X1   g615(.A(new_n816_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g616(.A1(new_n805_), .A2(new_n231_), .A3(new_n709_), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n656_), .B(new_n802_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT114), .B1(new_n819_), .B2(new_n231_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n807_), .A2(new_n709_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(G106gat), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n820_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n820_), .B2(new_n823_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n818_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT53), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n829_), .B(new_n818_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1339gat));
  INV_X1    g630(.A(new_n390_), .ZN(new_n832_));
  OAI22_X1  g631(.A1(new_n373_), .A2(new_n377_), .B1(new_n376_), .B2(new_n368_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n387_), .B1(new_n833_), .B2(new_n366_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n367_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n836_));
  OAI211_X1 g635(.A(G229gat), .B(G233gat), .C1(new_n836_), .C2(KEYINPUT118), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n836_), .A2(KEYINPUT118), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n834_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n832_), .B1(new_n839_), .B2(KEYINPUT119), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n355_), .A2(new_n360_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n834_), .B(new_n842_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n840_), .A2(new_n841_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n350_), .A2(new_n352_), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n350_), .A2(new_n352_), .A3(KEYINPUT116), .A4(new_n845_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n348_), .A2(new_n845_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n351_), .A2(new_n343_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(G230gat), .A3(G233gat), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .A4(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n360_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT56), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n853_), .A2(new_n856_), .A3(new_n360_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n844_), .A2(KEYINPUT58), .A3(new_n855_), .A4(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n299_), .B1(new_n858_), .B2(KEYINPUT121), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n844_), .A2(KEYINPUT120), .A3(new_n855_), .A4(new_n857_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n840_), .A2(new_n857_), .A3(new_n841_), .A4(new_n843_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n855_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n861_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n860_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n862_), .A2(new_n863_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(new_n868_), .A3(KEYINPUT58), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n859_), .A2(new_n866_), .A3(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n840_), .A2(new_n361_), .A3(new_n843_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n853_), .A2(KEYINPUT117), .A3(new_n856_), .A4(new_n360_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n872_), .A2(new_n841_), .A3(new_n393_), .A4(new_n391_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n853_), .A2(new_n360_), .B1(KEYINPUT117), .B2(new_n856_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n871_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n712_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n875_), .A2(KEYINPUT57), .A3(new_n712_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n337_), .B1(new_n870_), .B2(new_n880_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n339_), .A2(new_n365_), .A3(new_n779_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n881_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n685_), .A2(new_n664_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n886_), .A2(new_n887_), .A3(new_n676_), .A4(new_n888_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n875_), .A2(KEYINPUT57), .A3(new_n712_), .ZN(new_n890_));
  AOI21_X1  g689(.A(KEYINPUT57), .B1(new_n875_), .B2(new_n712_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n859_), .A2(new_n866_), .A3(new_n869_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n338_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n676_), .B(new_n888_), .C1(new_n894_), .C2(new_n884_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(KEYINPUT59), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n889_), .A2(new_n896_), .A3(new_n779_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G113gat), .ZN(new_n898_));
  INV_X1    g697(.A(new_n895_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n410_), .A3(new_n779_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1340gat));
  NAND3_X1  g700(.A1(new_n889_), .A2(new_n896_), .A3(new_n365_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G120gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(KEYINPUT60), .B1(new_n365_), .B2(new_n453_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n453_), .A2(KEYINPUT60), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n899_), .A2(KEYINPUT122), .A3(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n908_));
  INV_X1    g707(.A(new_n906_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n895_), .B2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n907_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n903_), .A2(new_n911_), .ZN(G1341gat));
  AOI21_X1  g711(.A(G127gat), .B1(new_n899_), .B2(new_n338_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n889_), .A2(new_n896_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n337_), .A2(new_n401_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT123), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n913_), .B1(new_n914_), .B2(new_n916_), .ZN(G1342gat));
  NAND3_X1  g716(.A1(new_n889_), .A2(new_n896_), .A3(new_n725_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(G134gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n899_), .A2(new_n399_), .A3(new_n680_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1343gat));
  NOR2_X1   g720(.A1(new_n685_), .A2(new_n665_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n676_), .B(new_n922_), .C1(new_n894_), .C2(new_n884_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n779_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n365_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g727(.A1(new_n923_), .A2(new_n337_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT61), .B(G155gat), .Z(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT124), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n929_), .B(new_n931_), .ZN(G1346gat));
  NOR3_X1   g731(.A1(new_n923_), .A2(new_n417_), .A3(new_n299_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n417_), .B1(new_n923_), .B2(new_n712_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(KEYINPUT125), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n936_), .B(new_n417_), .C1(new_n923_), .C2(new_n712_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n933_), .B1(new_n935_), .B2(new_n937_), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n894_), .A2(new_n884_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n676_), .A2(new_n671_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n664_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  OAI21_X1  g741(.A(KEYINPUT126), .B1(new_n939_), .B2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n944_));
  INV_X1    g743(.A(new_n942_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n886_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n943_), .A2(new_n946_), .A3(new_n779_), .A4(new_n522_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n886_), .A2(new_n779_), .A3(new_n945_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n948_), .A2(new_n949_), .A3(G169gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n948_), .B2(G169gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n947_), .B1(new_n950_), .B2(new_n951_), .ZN(G1348gat));
  NAND3_X1  g751(.A1(new_n943_), .A2(new_n946_), .A3(new_n365_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n939_), .A2(new_n942_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n778_), .A2(new_n523_), .ZN(new_n955_));
  AOI22_X1  g754(.A1(new_n953_), .A2(new_n523_), .B1(new_n954_), .B2(new_n955_), .ZN(G1349gat));
  AOI21_X1  g755(.A(G183gat), .B1(new_n954_), .B2(new_n338_), .ZN(new_n957_));
  AND2_X1   g756(.A1(new_n943_), .A2(new_n946_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n337_), .A2(new_n504_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n957_), .B1(new_n958_), .B2(new_n959_), .ZN(G1350gat));
  NAND3_X1  g759(.A1(new_n943_), .A2(new_n946_), .A3(new_n725_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(G190gat), .ZN(new_n962_));
  NAND4_X1  g761(.A1(new_n943_), .A2(new_n946_), .A3(new_n509_), .A4(new_n680_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(G1351gat));
  NAND3_X1  g763(.A1(new_n940_), .A2(new_n629_), .A3(new_n709_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n939_), .A2(new_n965_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(new_n779_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g767(.A1(new_n966_), .A2(new_n365_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g769(.A(new_n337_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n966_), .A2(new_n971_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n973_));
  XOR2_X1   g772(.A(new_n973_), .B(KEYINPUT127), .Z(new_n974_));
  XNOR2_X1  g773(.A(new_n972_), .B(new_n974_), .ZN(G1354gat));
  INV_X1    g774(.A(G218gat), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n966_), .A2(new_n976_), .A3(new_n680_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n966_), .A2(new_n725_), .ZN(new_n978_));
  INV_X1    g777(.A(new_n978_), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n977_), .B1(new_n979_), .B2(new_n976_), .ZN(G1355gat));
endmodule


