//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_;
  XOR2_X1   g000(.A(G141gat), .B(G148gat), .Z(new_n202_));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT82), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT82), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G155gat), .A3(G162gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT83), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n204_), .B(new_n210_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n213_));
  AOI211_X1 g012(.A(KEYINPUT83), .B(new_n209_), .C1(new_n206_), .C2(new_n208_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n202_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT84), .ZN(new_n216_));
  INV_X1    g015(.A(G141gat), .ZN(new_n217_));
  INV_X1    g016(.A(G148gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT3), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n216_), .B1(new_n222_), .B2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n207_), .B1(G155gat), .B2(G162gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n205_), .A2(KEYINPUT82), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n204_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT85), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n206_), .A2(new_n208_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT85), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n204_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n219_), .A2(new_n221_), .ZN(new_n235_));
  AND3_X1   g034(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(new_n223_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n237_), .A3(KEYINPUT84), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n227_), .A2(new_n231_), .A3(new_n234_), .A4(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n215_), .A2(new_n239_), .A3(KEYINPUT93), .ZN(new_n240_));
  XOR2_X1   g039(.A(G127gat), .B(G134gat), .Z(new_n241_));
  XOR2_X1   g040(.A(G113gat), .B(G120gat), .Z(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G225gat), .A2(G233gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n243_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n215_), .A2(new_n246_), .A3(new_n239_), .A4(KEYINPUT93), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n244_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n244_), .A2(new_n247_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n215_), .A2(new_n239_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n243_), .A2(KEYINPUT4), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n249_), .A2(KEYINPUT4), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n248_), .B1(new_n252_), .B2(new_n245_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G1gat), .B(G29gat), .Z(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT94), .B(G85gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT0), .B(G57gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT96), .ZN(new_n260_));
  INV_X1    g059(.A(new_n258_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n248_), .B(new_n261_), .C1(new_n252_), .C2(new_n245_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n259_), .A2(new_n260_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n253_), .A2(KEYINPUT96), .A3(new_n258_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G226gat), .A2(G233gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT19), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT23), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT23), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(G183gat), .A3(G190gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n271_), .A3(KEYINPUT79), .ZN(new_n272_));
  INV_X1    g071(.A(G183gat), .ZN(new_n273_));
  INV_X1    g072(.A(G190gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT79), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n276_), .A2(new_n270_), .A3(G183gat), .A4(G190gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n272_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(KEYINPUT78), .A2(G169gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(G176gat), .B1(new_n279_), .B2(KEYINPUT22), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT22), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(KEYINPUT78), .A3(G169gat), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n280_), .A2(new_n282_), .B1(G169gat), .B2(G176gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT77), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT26), .B1(new_n285_), .B2(new_n274_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n273_), .A2(KEYINPUT25), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(G183gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT26), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(KEYINPUT77), .A3(G190gat), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n286_), .A2(new_n287_), .A3(new_n289_), .A4(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n269_), .A2(new_n271_), .ZN(new_n293_));
  INV_X1    g092(.A(G169gat), .ZN(new_n294_));
  INV_X1    g093(.A(G176gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(KEYINPUT24), .A3(new_n297_), .ZN(new_n298_));
  OR3_X1    g097(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n292_), .A2(new_n293_), .A3(new_n298_), .A4(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(KEYINPUT87), .A2(KEYINPUT21), .ZN(new_n301_));
  INV_X1    g100(.A(G204gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G197gat), .ZN(new_n303_));
  INV_X1    g102(.A(G197gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G204gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(KEYINPUT87), .A2(KEYINPUT21), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n301_), .A2(new_n303_), .A3(new_n305_), .A4(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G211gat), .B(G218gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT86), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n303_), .A2(new_n305_), .A3(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n302_), .A2(KEYINPUT86), .A3(G197gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT21), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n307_), .B(new_n308_), .C1(new_n310_), .C2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n308_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n303_), .A2(new_n305_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(KEYINPUT21), .A3(new_n315_), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n284_), .A2(new_n300_), .B1(new_n313_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n293_), .A2(new_n275_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n281_), .A2(G169gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n294_), .A2(KEYINPUT22), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n295_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n297_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n287_), .A2(new_n289_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n274_), .A2(KEYINPUT26), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n290_), .A2(G190gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT91), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n290_), .A2(G190gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n274_), .A2(KEYINPUT26), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT91), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n323_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n272_), .A2(new_n298_), .A3(new_n277_), .A4(new_n299_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n322_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n313_), .A2(new_n316_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT20), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT95), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n317_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  OAI211_X1 g136(.A(KEYINPUT95), .B(KEYINPUT20), .C1(new_n333_), .C2(new_n334_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n267_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n284_), .A2(new_n300_), .A3(new_n313_), .A4(new_n316_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n321_), .A2(new_n297_), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n269_), .A2(new_n271_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n332_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n323_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n330_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n329_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n343_), .B1(new_n344_), .B2(new_n348_), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n307_), .A2(new_n308_), .ZN(new_n350_));
  OAI211_X1 g149(.A(KEYINPUT21), .B(new_n311_), .C1(new_n315_), .C2(KEYINPUT86), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n315_), .A2(KEYINPUT21), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n350_), .A2(new_n351_), .B1(new_n314_), .B2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n340_), .B(KEYINPUT20), .C1(new_n349_), .C2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(new_n266_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n339_), .A2(new_n355_), .ZN(new_n356_));
  OR3_X1    g155(.A1(new_n335_), .A2(new_n266_), .A3(new_n317_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT92), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT20), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n359_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n360_));
  AOI211_X1 g159(.A(new_n358_), .B(new_n267_), .C1(new_n360_), .C2(new_n340_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT92), .B1(new_n354_), .B2(new_n266_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n357_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G8gat), .B(G36gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT18), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT32), .ZN(new_n368_));
  MUX2_X1   g167(.A(new_n356_), .B(new_n363_), .S(new_n368_), .Z(new_n369_));
  NAND3_X1  g168(.A1(new_n263_), .A2(new_n264_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT33), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n259_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n249_), .A2(KEYINPUT4), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n250_), .A2(new_n251_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n245_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n245_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n258_), .B1(new_n249_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n367_), .B(new_n357_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n367_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n363_), .A2(new_n380_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n378_), .A2(new_n379_), .A3(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n253_), .A2(KEYINPUT33), .A3(new_n258_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n372_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n370_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(KEYINPUT88), .A2(G228gat), .A3(G233gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n334_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT88), .B1(G228gat), .B2(G233gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n232_), .A2(KEYINPUT1), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT83), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n211_), .A2(new_n212_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n392_), .A2(new_n393_), .A3(new_n204_), .A4(new_n210_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n235_), .A2(new_n237_), .A3(KEYINPUT84), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT84), .B1(new_n235_), .B2(new_n237_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n233_), .B1(new_n232_), .B2(new_n204_), .ZN(new_n398_));
  AOI211_X1 g197(.A(KEYINPUT85), .B(new_n203_), .C1(new_n206_), .C2(new_n208_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n394_), .A2(new_n202_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT29), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n388_), .B(new_n390_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n402_), .B1(new_n215_), .B2(new_n239_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n389_), .B1(new_n404_), .B2(new_n387_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G78gat), .B(G106gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n403_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n406_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n250_), .A2(KEYINPUT29), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n390_), .B1(new_n410_), .B2(new_n388_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n404_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n409_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT89), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n403_), .A2(new_n405_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT89), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(new_n409_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n408_), .B1(new_n414_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT28), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n401_), .A2(new_n419_), .A3(new_n402_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT28), .B1(new_n250_), .B2(KEYINPUT29), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G22gat), .B(G50gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT90), .B1(new_n418_), .B2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n416_), .B1(new_n415_), .B2(new_n409_), .ZN(new_n426_));
  AOI211_X1 g225(.A(KEYINPUT89), .B(new_n406_), .C1(new_n403_), .C2(new_n405_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n407_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n429_));
  INV_X1    g228(.A(new_n424_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n408_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n425_), .A2(new_n431_), .B1(new_n413_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n385_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n354_), .A2(new_n266_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n358_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n354_), .A2(KEYINPUT92), .A3(new_n266_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n367_), .B1(new_n439_), .B2(new_n357_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n379_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n435_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n380_), .B1(new_n339_), .B2(new_n355_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(KEYINPUT27), .A3(new_n379_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n445_), .B1(new_n264_), .B2(new_n263_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n424_), .A2(new_n407_), .A3(new_n413_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n429_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n446_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n434_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n284_), .A2(new_n300_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT30), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n246_), .A2(KEYINPUT31), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT31), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT81), .B1(new_n243_), .B2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n455_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G71gat), .B(G99gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(G43gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G227gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(G15gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n463_), .B(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(new_n454_), .B2(KEYINPUT80), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n456_), .A2(new_n458_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n454_), .B2(KEYINPUT80), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n461_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n468_), .B1(new_n461_), .B2(new_n470_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n425_), .A2(new_n431_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n263_), .A2(new_n264_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT27), .B1(new_n381_), .B2(new_n379_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n443_), .A2(KEYINPUT27), .A3(new_n379_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n476_), .A2(new_n477_), .A3(new_n473_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n474_), .A2(new_n475_), .A3(new_n478_), .A4(new_n447_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT97), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n433_), .A2(KEYINPUT97), .A3(new_n475_), .A4(new_n478_), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n452_), .A2(new_n473_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G1gat), .B(G8gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT73), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G22gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n465_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G15gat), .A2(G22gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G1gat), .A2(G8gat), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n488_), .A2(new_n489_), .B1(KEYINPUT14), .B2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n486_), .B(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G29gat), .B(G36gat), .Z(new_n493_));
  XOR2_X1   g292(.A(G43gat), .B(G50gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT75), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n492_), .A2(new_n495_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G229gat), .A2(G233gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n492_), .A2(new_n495_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT15), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n495_), .B(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n504_), .B2(new_n492_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n505_), .A2(new_n500_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n501_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G113gat), .B(G141gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G169gat), .B(G197gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n501_), .A2(new_n506_), .A3(new_n510_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT76), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n512_), .A2(KEYINPUT76), .A3(new_n513_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n483_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT98), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT70), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT13), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G57gat), .B(G64gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT11), .ZN(new_n527_));
  XOR2_X1   g326(.A(G71gat), .B(G78gat), .Z(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n526_), .A2(KEYINPUT11), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n527_), .A2(new_n528_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT12), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n536_));
  NOR2_X1   g335(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n537_));
  OAI21_X1  g336(.A(G92gat), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT9), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT66), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT66), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n542_), .A3(new_n539_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(G85gat), .A2(G92gat), .ZN(new_n544_));
  AND2_X1   g343(.A1(G85gat), .A2(G92gat), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n544_), .B1(new_n545_), .B2(KEYINPUT9), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n541_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT10), .B(G99gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n549_), .A2(KEYINPUT6), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(KEYINPUT6), .ZN(new_n551_));
  OAI22_X1  g350(.A1(new_n548_), .A2(G106gat), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n545_), .A2(new_n544_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n550_), .A2(new_n551_), .ZN(new_n556_));
  OR3_X1    g355(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n555_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT8), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n558_), .B(new_n557_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT8), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n563_), .A3(new_n555_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n532_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(new_n530_), .B2(new_n529_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n554_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n554_), .B2(new_n565_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n535_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G230gat), .A2(G233gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT64), .Z(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT67), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n569_), .A2(new_n574_), .A3(KEYINPUT12), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n562_), .A2(new_n563_), .A3(new_n555_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n563_), .B1(new_n562_), .B2(new_n555_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n546_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n540_), .B2(KEYINPUT66), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n552_), .B1(new_n580_), .B2(new_n543_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n533_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT67), .B1(new_n582_), .B2(new_n534_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n570_), .B(new_n573_), .C1(new_n575_), .C2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n572_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G120gat), .B(G148gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT5), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G176gat), .B(G204gat), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n587_), .B(new_n588_), .Z(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n584_), .A2(new_n585_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT69), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(KEYINPUT68), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n592_), .B1(new_n591_), .B2(KEYINPUT68), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n584_), .A2(new_n585_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n589_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n594_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n597_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n591_), .A2(KEYINPUT68), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT69), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n601_), .B2(new_n593_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n524_), .B(new_n525_), .C1(new_n598_), .C2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n597_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(new_n599_), .A3(new_n593_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n522_), .A4(new_n523_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G134gat), .B(G162gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(KEYINPUT36), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n504_), .B1(new_n581_), .B2(new_n578_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n495_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n554_), .A2(new_n565_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT72), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT34), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n618_), .B(new_n619_), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n615_), .A2(new_n616_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n610_), .A2(KEYINPUT36), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n622_), .B(new_n623_), .C1(new_n615_), .C2(new_n618_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n621_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n611_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT37), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n624_), .A2(new_n625_), .A3(new_n611_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n629_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT37), .B1(new_n631_), .B2(new_n626_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n567_), .B(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(new_n492_), .ZN(new_n636_));
  XOR2_X1   g435(.A(G127gat), .B(G155gat), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT16), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G183gat), .B(G211gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT17), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n640_), .A2(new_n641_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n636_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n636_), .A2(new_n642_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n645_), .A2(KEYINPUT74), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(KEYINPUT74), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n644_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n607_), .A2(new_n633_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n521_), .A2(new_n650_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n651_), .A2(G1gat), .A3(new_n475_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT38), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT99), .Z(new_n654_));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n655_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n631_), .A2(KEYINPUT100), .A3(new_n626_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n481_), .A2(new_n482_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n473_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n434_), .B2(new_n451_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT101), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n607_), .A2(new_n519_), .A3(new_n649_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n475_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G1gat), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n654_), .B(new_n669_), .C1(KEYINPUT38), .C2(new_n652_), .ZN(G1324gat));
  INV_X1    g469(.A(new_n651_), .ZN(new_n671_));
  INV_X1    g470(.A(G8gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n445_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n666_), .A2(new_n445_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n675_), .B2(G8gat), .ZN(new_n676_));
  AOI211_X1 g475(.A(KEYINPUT39), .B(new_n672_), .C1(new_n666_), .C2(new_n445_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(G1325gat));
  AOI21_X1  g479(.A(new_n465_), .B1(new_n666_), .B2(new_n661_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT41), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n671_), .A2(new_n465_), .A3(new_n661_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1326gat));
  AOI21_X1  g483(.A(new_n487_), .B1(new_n666_), .B2(new_n450_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT42), .Z(new_n686_));
  NAND3_X1  g485(.A1(new_n671_), .A2(new_n487_), .A3(new_n450_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1327gat));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n630_), .A2(new_n632_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT43), .B1(new_n690_), .B2(KEYINPUT103), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n692_), .B1(new_n483_), .B2(new_n690_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n633_), .B(new_n691_), .C1(new_n660_), .C2(new_n662_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n603_), .A2(new_n518_), .A3(new_n649_), .A4(new_n606_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT102), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n603_), .A2(new_n606_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n518_), .A4(new_n649_), .ZN(new_n699_));
  AOI22_X1  g498(.A1(new_n693_), .A2(new_n694_), .B1(new_n696_), .B2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n689_), .B1(new_n700_), .B2(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n693_), .A2(new_n694_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n699_), .A2(new_n696_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(KEYINPUT104), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707_));
  AND4_X1   g506(.A1(new_n707_), .A2(new_n702_), .A3(KEYINPUT44), .A4(new_n703_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n700_), .B2(KEYINPUT44), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n701_), .B(new_n706_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT106), .B1(new_n710_), .B2(new_n475_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n706_), .A2(new_n701_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n713_));
  OAI21_X1  g512(.A(KEYINPUT105), .B1(new_n704_), .B2(new_n705_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n700_), .A2(new_n707_), .A3(KEYINPUT44), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n712_), .A2(new_n713_), .A3(new_n716_), .A4(new_n667_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n711_), .A2(G29gat), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n658_), .A2(new_n649_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n607_), .A2(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n521_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(G29gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n667_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n718_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT107), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n718_), .A2(new_n726_), .A3(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1328gat));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729_));
  INV_X1    g528(.A(new_n445_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n710_), .B2(new_n730_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n712_), .A2(KEYINPUT108), .A3(new_n716_), .A4(new_n445_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(G36gat), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(G36gat), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n445_), .B(KEYINPUT109), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n721_), .A2(new_n734_), .A3(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT45), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n733_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(KEYINPUT46), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n733_), .B(new_n738_), .C1(new_n740_), .C2(KEYINPUT46), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1329gat));
  OAI21_X1  g543(.A(G43gat), .B1(new_n710_), .B2(new_n473_), .ZN(new_n745_));
  INV_X1    g544(.A(G43gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n721_), .A2(new_n746_), .A3(new_n661_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g548(.A(G50gat), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n710_), .A2(new_n750_), .A3(new_n433_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G50gat), .B1(new_n721_), .B2(new_n450_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1331gat));
  AND4_X1   g552(.A1(new_n519_), .A2(new_n664_), .A3(new_n648_), .A4(new_n607_), .ZN(new_n754_));
  INV_X1    g553(.A(G57gat), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n475_), .A2(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n483_), .A2(new_n518_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n697_), .A2(new_n649_), .A3(new_n633_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n475_), .B1(new_n759_), .B2(KEYINPUT111), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(KEYINPUT111), .B2(new_n759_), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n754_), .A2(new_n756_), .B1(new_n761_), .B2(new_n755_), .ZN(G1332gat));
  INV_X1    g561(.A(G64gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n754_), .B2(new_n736_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT48), .Z(new_n765_));
  NAND2_X1  g564(.A1(new_n736_), .A2(new_n763_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT112), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n765_), .B1(new_n759_), .B2(new_n767_), .ZN(G1333gat));
  INV_X1    g567(.A(G71gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n754_), .B2(new_n661_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT49), .Z(new_n771_));
  INV_X1    g570(.A(new_n759_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n769_), .A3(new_n661_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1334gat));
  INV_X1    g573(.A(G78gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n754_), .B2(new_n450_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT50), .Z(new_n777_));
  NAND3_X1  g576(.A1(new_n772_), .A2(new_n775_), .A3(new_n450_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1335gat));
  OR2_X1    g578(.A1(new_n702_), .A2(KEYINPUT113), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n702_), .A2(KEYINPUT113), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n697_), .A2(new_n518_), .A3(new_n648_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n536_), .A2(new_n537_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n783_), .A2(new_n475_), .A3(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n697_), .A2(new_n719_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n757_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(G85gat), .B1(new_n788_), .B2(new_n667_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n785_), .A2(new_n789_), .ZN(G1336gat));
  OAI21_X1  g589(.A(G92gat), .B1(new_n783_), .B2(new_n735_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n730_), .A2(G92gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n787_), .B2(new_n792_), .ZN(G1337gat));
  OAI21_X1  g592(.A(G99gat), .B1(new_n783_), .B2(new_n473_), .ZN(new_n794_));
  OR3_X1    g593(.A1(new_n787_), .A2(new_n473_), .A3(new_n548_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g596(.A1(new_n702_), .A2(new_n450_), .A3(new_n782_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(G106gat), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n799_), .B(KEYINPUT52), .Z(new_n800_));
  NOR3_X1   g599(.A1(new_n787_), .A2(G106gat), .A3(new_n433_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n802_), .B(KEYINPUT53), .Z(G1339gat));
  NAND2_X1  g602(.A1(new_n650_), .A2(new_n519_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n584_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(KEYINPUT115), .A3(KEYINPUT55), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n584_), .B2(new_n810_), .ZN(new_n811_));
  XOR2_X1   g610(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n812_));
  OAI21_X1  g611(.A(new_n570_), .B1(new_n575_), .B2(new_n583_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n572_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n808_), .B(new_n811_), .C1(new_n814_), .C2(new_n807_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n589_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n815_), .A2(KEYINPUT56), .A3(new_n589_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(KEYINPUT119), .A3(new_n819_), .ZN(new_n820_));
  OR3_X1    g619(.A1(new_n816_), .A2(KEYINPUT119), .A3(new_n817_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n510_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n505_), .A2(KEYINPUT117), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n500_), .B1(new_n505_), .B2(KEYINPUT117), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n825_), .A2(KEYINPUT118), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(KEYINPUT118), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n826_), .A2(new_n513_), .A3(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n820_), .A2(new_n821_), .A3(new_n591_), .A4(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n830_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n633_), .A3(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n518_), .A2(new_n591_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n818_), .A2(new_n835_), .A3(new_n819_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n816_), .A2(KEYINPUT116), .A3(new_n817_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n828_), .A2(new_n605_), .A3(new_n604_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n659_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(KEYINPUT57), .A3(new_n659_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n833_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n806_), .B1(new_n845_), .B2(new_n649_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n433_), .A2(new_n667_), .A3(new_n478_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(G113gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n518_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n847_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n845_), .A2(new_n649_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT59), .B(new_n853_), .C1(new_n854_), .C2(new_n806_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n519_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n850_), .B1(new_n856_), .B2(new_n849_), .ZN(G1340gat));
  INV_X1    g656(.A(G120gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n697_), .B2(KEYINPUT60), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(KEYINPUT60), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(KEYINPUT120), .B2(new_n860_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n848_), .B(new_n861_), .C1(KEYINPUT120), .C2(new_n859_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n697_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n858_), .ZN(G1341gat));
  INV_X1    g663(.A(G127gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n848_), .A2(new_n865_), .A3(new_n648_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n649_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n865_), .ZN(G1342gat));
  INV_X1    g667(.A(G134gat), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n852_), .A2(new_n855_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n633_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n848_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n658_), .A2(new_n869_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT121), .B1(new_n871_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n690_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n877_));
  OAI221_X1 g676(.A(new_n876_), .B1(new_n872_), .B2(new_n873_), .C1(new_n877_), .C2(new_n869_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n878_), .ZN(G1343gat));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n735_), .A2(new_n473_), .A3(new_n450_), .A4(new_n667_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT122), .ZN(new_n882_));
  OR3_X1    g681(.A1(new_n846_), .A2(new_n880_), .A3(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n880_), .B1(new_n846_), .B2(new_n882_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n519_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n217_), .ZN(G1344gat));
  AOI21_X1  g685(.A(new_n697_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT124), .B(G148gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1345gat));
  AOI21_X1  g688(.A(new_n649_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n890_), .B(new_n892_), .ZN(G1346gat));
  NAND2_X1  g692(.A1(new_n883_), .A2(new_n884_), .ZN(new_n894_));
  INV_X1    g693(.A(G162gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n894_), .A2(new_n895_), .A3(new_n658_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n690_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n895_), .ZN(G1347gat));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n846_), .A2(new_n735_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n450_), .A2(new_n667_), .A3(new_n473_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n519_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n899_), .B1(new_n903_), .B2(new_n294_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n905_));
  OAI211_X1 g704(.A(KEYINPUT62), .B(G169gat), .C1(new_n902_), .C2(new_n519_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n904_), .A2(new_n905_), .A3(new_n906_), .ZN(G1348gat));
  NOR2_X1   g706(.A1(new_n902_), .A2(new_n697_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(new_n295_), .ZN(G1349gat));
  NAND3_X1  g708(.A1(new_n900_), .A2(new_n648_), .A3(new_n901_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n345_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(new_n273_), .B2(new_n910_), .ZN(G1350gat));
  NAND2_X1  g711(.A1(new_n326_), .A2(new_n330_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n900_), .A2(new_n913_), .A3(new_n658_), .A4(new_n901_), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n900_), .A2(new_n633_), .A3(new_n901_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n915_), .B2(new_n274_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(KEYINPUT125), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n918_), .B(new_n914_), .C1(new_n915_), .C2(new_n274_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1351gat));
  NOR3_X1   g719(.A1(new_n433_), .A2(new_n667_), .A3(new_n661_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n900_), .A2(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n519_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(new_n304_), .ZN(G1352gat));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n697_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n302_), .ZN(G1353gat));
  AND3_X1   g725(.A1(new_n900_), .A2(new_n648_), .A3(new_n921_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT63), .B(G211gat), .Z(new_n928_));
  AOI21_X1  g727(.A(KEYINPUT126), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n900_), .A2(new_n648_), .A3(new_n921_), .A4(new_n928_), .ZN(new_n930_));
  OR2_X1    g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n927_), .B2(new_n931_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n929_), .B1(KEYINPUT126), .B2(new_n932_), .ZN(G1354gat));
  INV_X1    g732(.A(G218gat), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n900_), .A2(new_n934_), .A3(new_n658_), .A4(new_n921_), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n900_), .A2(new_n633_), .A3(new_n921_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n936_), .B2(new_n934_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(KEYINPUT127), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n939_), .B(new_n935_), .C1(new_n936_), .C2(new_n934_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1355gat));
endmodule


