//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n957_, new_n958_, new_n960_,
    new_n961_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_, new_n985_, new_n986_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT36), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT66), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n212_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT7), .ZN(new_n215_));
  INV_X1    g014(.A(G99gat), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT6), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n218_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n209_), .B1(new_n214_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT8), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n226_), .B(new_n209_), .C1(new_n214_), .C2(new_n223_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT9), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n208_), .A2(new_n229_), .ZN(new_n230_));
  OAI211_X1 g029(.A(KEYINPUT65), .B(new_n230_), .C1(new_n209_), .C2(new_n229_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n221_), .A2(new_n222_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT10), .B(G99gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n232_), .B1(new_n234_), .B2(new_n217_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n229_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n230_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n231_), .A2(new_n235_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n228_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G36gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G29gat), .ZN(new_n243_));
  INV_X1    g042(.A(G29gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G36gat), .ZN(new_n245_));
  INV_X1    g044(.A(G43gat), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n243_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n246_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT68), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n244_), .A2(G36gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n242_), .A2(G29gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(G43gat), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n243_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n249_), .A2(G50gat), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(G50gat), .B1(new_n249_), .B2(new_n255_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT15), .ZN(new_n258_));
  NOR3_X1   g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G50gat), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n247_), .A2(new_n248_), .A3(KEYINPUT68), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n253_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n249_), .A2(new_n255_), .A3(G50gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT15), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n241_), .B1(new_n259_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n235_), .A2(new_n239_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n268_), .A2(new_n231_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(new_n264_), .A4(new_n263_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n228_), .A2(new_n264_), .A3(new_n263_), .A4(new_n240_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT69), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n266_), .A2(new_n267_), .A3(new_n271_), .A4(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G232gat), .A2(G233gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n275_), .B(KEYINPUT34), .Z(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n258_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n263_), .A2(KEYINPUT15), .A3(new_n264_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n280_), .A2(new_n241_), .B1(KEYINPUT69), .B2(new_n272_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n276_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n281_), .A2(new_n267_), .A3(new_n271_), .A4(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT35), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n281_), .A2(new_n285_), .A3(new_n271_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n277_), .A2(new_n283_), .A3(KEYINPUT35), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n206_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n277_), .A2(new_n283_), .A3(KEYINPUT35), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n286_), .B1(new_n277_), .B2(new_n283_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n292_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n288_), .A2(new_n292_), .A3(new_n289_), .A4(new_n296_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n291_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT37), .B1(new_n290_), .B2(KEYINPUT72), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n288_), .A2(new_n289_), .A3(new_n296_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT71), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n290_), .B1(new_n305_), .B2(new_n298_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n301_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G230gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT64), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G57gat), .B(G64gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT67), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n312_), .A2(new_n313_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT11), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n316_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT11), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(new_n319_), .A3(new_n314_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G71gat), .B(G78gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n317_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(KEYINPUT11), .B(new_n321_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n241_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n324_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n269_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(KEYINPUT12), .A3(new_n328_), .ZN(new_n329_));
  OR3_X1    g128(.A1(new_n327_), .A2(new_n269_), .A3(KEYINPUT12), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n311_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n310_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G120gat), .B(G148gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(G204gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(KEYINPUT5), .B(G176gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n333_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n333_), .A2(new_n337_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT13), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n338_), .A2(KEYINPUT13), .A3(new_n339_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G127gat), .B(G155gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G183gat), .B(G211gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT17), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G15gat), .B(G22gat), .ZN(new_n352_));
  INV_X1    g151(.A(G1gat), .ZN(new_n353_));
  INV_X1    g152(.A(G8gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT14), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G1gat), .B(G8gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT73), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G231gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n361_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n327_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n325_), .A3(new_n363_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n351_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n350_), .A2(KEYINPUT17), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(new_n368_), .A3(new_n366_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n365_), .A2(KEYINPUT75), .A3(new_n368_), .A4(new_n366_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n367_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AOI211_X1 g174(.A(KEYINPUT76), .B(new_n367_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n308_), .A2(new_n345_), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G169gat), .B(G197gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT80), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G113gat), .B(G141gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n380_), .B(new_n381_), .Z(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G229gat), .A2(G233gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n263_), .A2(new_n264_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT77), .B1(new_n387_), .B2(new_n358_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n358_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n389_), .A2(new_n263_), .A3(new_n390_), .A4(new_n264_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n387_), .A2(new_n358_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n386_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n389_), .B1(new_n264_), .B2(new_n263_), .ZN(new_n395_));
  AOI211_X1 g194(.A(KEYINPUT78), .B(new_n395_), .C1(new_n388_), .C2(new_n391_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n385_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT79), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT79), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n399_), .B(new_n385_), .C1(new_n394_), .C2(new_n396_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n280_), .A2(new_n358_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n392_), .A3(new_n384_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n383_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  AOI211_X1 g204(.A(new_n405_), .B(new_n382_), .C1(new_n398_), .C2(new_n400_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT81), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G141gat), .A2(G148gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT2), .ZN(new_n411_));
  INV_X1    g210(.A(G141gat), .ZN(new_n412_));
  INV_X1    g211(.A(G148gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(KEYINPUT3), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT3), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(G141gat), .B2(G148gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n411_), .A2(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(G155gat), .A2(G162gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(G155gat), .A2(G162gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n422_), .B1(new_n420_), .B2(KEYINPUT1), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT1), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n419_), .A2(KEYINPUT86), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT86), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(new_n422_), .B2(KEYINPUT1), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n423_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT85), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n430_), .A2(new_n431_), .B1(G141gat), .B2(G148gat), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n418_), .A2(new_n421_), .B1(new_n428_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G78gat), .B(G106gat), .Z(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G22gat), .B(G50gat), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n439_), .B(KEYINPUT28), .Z(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT87), .B(KEYINPUT29), .ZN(new_n443_));
  INV_X1    g242(.A(new_n417_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT2), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n410_), .B(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n421_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n428_), .A2(new_n432_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n443_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT21), .ZN(new_n450_));
  INV_X1    g249(.A(G211gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n451_), .A2(G218gat), .ZN(new_n452_));
  INV_X1    g251(.A(G218gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(G211gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n450_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G197gat), .B(G204gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(G211gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n451_), .A2(G218gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(KEYINPUT21), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n455_), .A2(new_n457_), .A3(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n456_), .A2(KEYINPUT21), .A3(new_n458_), .A4(new_n459_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n442_), .B1(new_n449_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT88), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT88), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n466_), .B(new_n442_), .C1(new_n449_), .C2(new_n463_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n434_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n469_), .A2(new_n463_), .A3(new_n442_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n441_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n472_));
  AOI211_X1 g271(.A(new_n470_), .B(new_n440_), .C1(new_n465_), .C2(new_n467_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n438_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n467_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n461_), .A2(new_n462_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n476_), .B1(new_n433_), .B2(new_n443_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n466_), .B1(new_n477_), .B2(new_n442_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n471_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n440_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n468_), .A2(new_n471_), .A3(new_n441_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n437_), .A3(new_n481_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n474_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G8gat), .B(G36gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT18), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(G64gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(G92gat), .ZN(new_n487_));
  INV_X1    g286(.A(G64gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n485_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G92gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n487_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G226gat), .A2(G233gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT19), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G183gat), .A2(G190gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT23), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT23), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(G183gat), .A3(G190gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT83), .ZN(new_n501_));
  INV_X1    g300(.A(G183gat), .ZN(new_n502_));
  INV_X1    g301(.A(G190gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT83), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G169gat), .A2(G176gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT22), .B(G169gat), .ZN(new_n512_));
  INV_X1    g311(.A(G176gat), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n505_), .A2(new_n509_), .A3(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(G169gat), .A2(G176gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(KEYINPUT24), .A3(new_n510_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT24), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n497_), .A2(new_n499_), .B1(new_n519_), .B2(new_n516_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT26), .B(G190gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT25), .B1(new_n502_), .B2(KEYINPUT82), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT25), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(G183gat), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n525_), .A2(KEYINPUT82), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n518_), .B(new_n520_), .C1(new_n523_), .C2(new_n526_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n515_), .A2(new_n527_), .B1(new_n462_), .B2(new_n461_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n512_), .A2(new_n513_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n510_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n500_), .A2(new_n504_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n500_), .A2(KEYINPUT90), .A3(new_n504_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n530_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n503_), .A2(KEYINPUT26), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT26), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(G190gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n502_), .A2(KEYINPUT25), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n536_), .A2(new_n538_), .A3(new_n539_), .A4(new_n525_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n520_), .A2(new_n540_), .A3(new_n518_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT20), .B1(new_n535_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n528_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  OAI211_X1 g344(.A(KEYINPUT95), .B(KEYINPUT20), .C1(new_n535_), .C2(new_n542_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n495_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT20), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n515_), .A2(new_n527_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n549_), .B2(new_n463_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT90), .B1(new_n500_), .B2(new_n504_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(G183gat), .A2(G190gat), .ZN(new_n552_));
  AOI211_X1 g351(.A(new_n532_), .B(new_n552_), .C1(new_n497_), .C2(new_n499_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n514_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT89), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n520_), .A2(new_n540_), .A3(new_n555_), .A4(new_n518_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n541_), .A2(KEYINPUT89), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n476_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n550_), .A2(new_n495_), .A3(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n492_), .B1(new_n547_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT96), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(KEYINPUT96), .B(new_n492_), .C1(new_n547_), .C2(new_n560_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT27), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n463_), .A2(new_n554_), .A3(new_n556_), .A4(new_n557_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n515_), .A2(new_n527_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n476_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(KEYINPUT20), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n495_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n550_), .A2(new_n494_), .A3(new_n559_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n492_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n565_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n563_), .A2(new_n564_), .A3(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G57gat), .B(G85gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G1gat), .B(G29gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G225gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT91), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n447_), .A2(new_n448_), .ZN(new_n584_));
  INV_X1    g383(.A(G134gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(G127gat), .ZN(new_n586_));
  INV_X1    g385(.A(G127gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(G134gat), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(G113gat), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(G120gat), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n590_), .A2(G120gat), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n589_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G113gat), .B(G120gat), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n584_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n433_), .A2(new_n596_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n583_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n599_), .A3(KEYINPUT4), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n596_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT4), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n583_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n581_), .B(new_n601_), .C1(new_n606_), .C2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n580_), .B1(new_n609_), .B2(new_n600_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(G71gat), .B(G99gat), .Z(new_n612_));
  XOR2_X1   g411(.A(G15gat), .B(G43gat), .Z(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  AND3_X1   g413(.A1(new_n515_), .A2(KEYINPUT30), .A3(new_n527_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT30), .B1(new_n515_), .B2(new_n527_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n614_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT30), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n567_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n515_), .A2(KEYINPUT30), .A3(new_n527_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n614_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n617_), .A2(new_n622_), .A3(new_n596_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n596_), .B1(new_n617_), .B2(new_n622_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G227gat), .A2(G233gat), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT84), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT31), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n623_), .A2(new_n624_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n617_), .A2(new_n622_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n597_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n617_), .A2(new_n622_), .A3(new_n596_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n627_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n611_), .A2(new_n629_), .A3(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n570_), .A2(new_n492_), .A3(new_n571_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n492_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n565_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n483_), .A2(new_n575_), .A3(new_n634_), .A4(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT97), .ZN(new_n639_));
  INV_X1    g438(.A(new_n636_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n570_), .A2(new_n571_), .A3(new_n492_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT27), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n564_), .A2(new_n574_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n643_), .B2(new_n563_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n644_), .A2(new_n645_), .A3(new_n483_), .A4(new_n634_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n639_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n629_), .A2(new_n633_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n611_), .B1(new_n474_), .B2(new_n482_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n650_), .A2(new_n575_), .A3(new_n637_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n474_), .A2(new_n482_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT93), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n447_), .A2(new_n448_), .A3(new_n596_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n654_), .A2(new_n603_), .A3(new_n607_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n653_), .B1(new_n655_), .B2(new_n580_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n598_), .A2(new_n599_), .A3(new_n583_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n581_), .A2(new_n657_), .A3(KEYINPUT93), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n602_), .A2(new_n607_), .A3(new_n605_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n656_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT94), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n656_), .A2(KEYINPUT94), .A3(new_n658_), .A4(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n610_), .A2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n635_), .A2(new_n636_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n610_), .A2(new_n665_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n664_), .A2(new_n666_), .A3(new_n667_), .A4(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n573_), .A2(KEYINPUT32), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n572_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n547_), .A2(new_n560_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n611_), .B(new_n671_), .C1(new_n670_), .C2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n652_), .B1(new_n669_), .B2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n649_), .B1(new_n651_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n647_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n378_), .A2(new_n409_), .A3(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n678_), .A2(new_n353_), .A3(new_n611_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT38), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n676_), .A2(new_n300_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n373_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n344_), .A2(new_n407_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n611_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G1gat), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n679_), .A2(new_n680_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n681_), .A2(new_n688_), .A3(new_n689_), .ZN(G1324gat));
  NOR2_X1   g489(.A1(new_n644_), .A2(G8gat), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n678_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G8gat), .B1(new_n686_), .B2(new_n644_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT98), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n692_), .B1(new_n695_), .B2(KEYINPUT39), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n693_), .A2(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(KEYINPUT39), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g500(.A(G15gat), .B1(new_n686_), .B2(new_n649_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT41), .Z(new_n703_));
  INV_X1    g502(.A(G15gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n678_), .A2(new_n704_), .A3(new_n648_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1326gat));
  NOR2_X1   g505(.A1(new_n483_), .A2(G22gat), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT100), .Z(new_n708_));
  NAND2_X1  g507(.A1(new_n678_), .A2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G22gat), .B1(new_n686_), .B2(new_n483_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n710_), .A2(KEYINPUT99), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(KEYINPUT99), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n711_), .A2(KEYINPUT42), .A3(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT42), .B1(new_n711_), .B2(new_n712_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n709_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT101), .Z(G1327gat));
  NOR2_X1   g515(.A1(new_n409_), .A2(new_n677_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n377_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n345_), .A2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n719_), .A2(new_n300_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n717_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G29gat), .B1(new_n721_), .B2(new_n611_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n303_), .A2(new_n676_), .A3(new_n307_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT43), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n303_), .A2(new_n676_), .A3(new_n307_), .A4(new_n725_), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n407_), .B(new_n719_), .C1(new_n724_), .C2(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(KEYINPUT102), .A2(KEYINPUT44), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n687_), .A2(new_n244_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n722_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT103), .ZN(G1328gat));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n733_));
  INV_X1    g532(.A(new_n644_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n242_), .B1(new_n729_), .B2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n644_), .A2(G36gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n717_), .A2(new_n720_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT104), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n717_), .A2(new_n720_), .A3(new_n739_), .A4(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n738_), .A2(KEYINPUT45), .A3(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n733_), .B1(new_n735_), .B2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT46), .ZN(G1329gat));
  AOI21_X1  g546(.A(G43gat), .B1(new_n721_), .B2(new_n648_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n649_), .A2(new_n246_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n729_), .B2(new_n749_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g550(.A(G50gat), .B1(new_n721_), .B2(new_n652_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n483_), .A2(new_n260_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n729_), .B2(new_n753_), .ZN(G1331gat));
  NAND2_X1  g553(.A1(new_n344_), .A2(new_n377_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n408_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n683_), .ZN(new_n757_));
  INV_X1    g556(.A(G57gat), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(new_n687_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n407_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n677_), .A2(new_n755_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n308_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT106), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT106), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n611_), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n759_), .B1(new_n765_), .B2(new_n758_), .ZN(G1332gat));
  OAI21_X1  g565(.A(G64gat), .B1(new_n757_), .B2(new_n644_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT48), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n734_), .A2(new_n488_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n762_), .B2(new_n769_), .ZN(G1333gat));
  OAI21_X1  g569(.A(G71gat), .B1(new_n757_), .B2(new_n649_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT49), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n649_), .A2(G71gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n762_), .B2(new_n773_), .ZN(G1334gat));
  OR3_X1    g573(.A1(new_n762_), .A2(G78gat), .A3(new_n483_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G78gat), .B1(new_n757_), .B2(new_n483_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(KEYINPUT50), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(KEYINPUT50), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n775_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT107), .Z(G1335gat));
  NAND3_X1  g579(.A1(new_n718_), .A2(new_n407_), .A3(new_n344_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n781_), .A2(new_n677_), .A3(new_n300_), .ZN(new_n782_));
  AOI21_X1  g581(.A(G85gat), .B1(new_n782_), .B2(new_n611_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n781_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n611_), .A2(G85gat), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT108), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n783_), .B1(new_n784_), .B2(new_n786_), .ZN(G1336gat));
  NAND3_X1  g586(.A1(new_n782_), .A2(new_n490_), .A3(new_n734_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n784_), .A2(new_n734_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(new_n490_), .ZN(G1337gat));
  NAND3_X1  g589(.A1(new_n782_), .A2(new_n648_), .A3(new_n234_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT109), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n216_), .B1(new_n784_), .B2(new_n648_), .ZN(new_n793_));
  OAI22_X1  g592(.A1(new_n792_), .A2(new_n793_), .B1(KEYINPUT110), .B2(KEYINPUT51), .ZN(new_n794_));
  NAND2_X1  g593(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n794_), .B(new_n795_), .ZN(G1338gat));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797_));
  INV_X1    g596(.A(new_n781_), .ZN(new_n798_));
  AOI221_X4 g597(.A(new_n290_), .B1(KEYINPUT72), .B2(KEYINPUT37), .C1(new_n305_), .C2(new_n298_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n305_), .A2(new_n298_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n301_), .B1(new_n800_), .B2(new_n291_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n725_), .B1(new_n802_), .B2(new_n676_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n726_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n652_), .B(new_n798_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT111), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n784_), .A2(new_n807_), .A3(new_n652_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n217_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n797_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n724_), .A2(new_n726_), .ZN(new_n812_));
  AND4_X1   g611(.A1(new_n807_), .A2(new_n812_), .A3(new_n652_), .A4(new_n798_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n807_), .B1(new_n784_), .B2(new_n652_), .ZN(new_n814_));
  OAI21_X1  g613(.A(G106gat), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n217_), .A2(KEYINPUT52), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(KEYINPUT112), .B(new_n817_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n811_), .A2(new_n816_), .A3(new_n820_), .A4(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n782_), .A2(new_n217_), .A3(new_n652_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT53), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n822_), .A2(new_n826_), .A3(new_n823_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1339gat));
  OAI21_X1  g627(.A(KEYINPUT54), .B1(new_n378_), .B2(new_n408_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n377_), .A2(new_n343_), .A3(new_n342_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n409_), .A2(new_n830_), .A3(new_n308_), .A4(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n829_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n392_), .A2(new_n393_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT78), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n392_), .A2(new_n386_), .A3(new_n393_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n399_), .B1(new_n839_), .B2(new_n385_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n400_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n403_), .B(new_n383_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n384_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n384_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n383_), .B1(new_n844_), .B2(new_n402_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n340_), .A2(new_n842_), .A3(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n329_), .A2(new_n311_), .A3(new_n330_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n331_), .B1(KEYINPUT55), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n850_), .B(new_n311_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n337_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT56), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(KEYINPUT114), .A3(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n854_), .B(new_n338_), .C1(new_n404_), .C2(new_n406_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n852_), .A2(new_n853_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT56), .B(new_n337_), .C1(new_n849_), .C2(new_n851_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n847_), .B1(new_n855_), .B2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n835_), .B1(new_n860_), .B2(new_n300_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n835_), .A3(new_n300_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n842_), .A2(new_n338_), .A3(new_n846_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT115), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n856_), .A2(new_n858_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n842_), .A2(new_n870_), .A3(new_n338_), .A4(new_n846_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n865_), .A2(new_n866_), .A3(new_n869_), .A4(new_n871_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n802_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n865_), .A2(new_n866_), .A3(new_n871_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n862_), .A2(new_n863_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n834_), .B1(new_n876_), .B2(new_n377_), .ZN(new_n877_));
  NOR4_X1   g676(.A1(new_n734_), .A2(new_n652_), .A3(new_n687_), .A4(new_n649_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(KEYINPUT59), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n877_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n875_), .A2(new_n802_), .A3(new_n872_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n863_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n861_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n884_), .A2(new_n684_), .B1(new_n829_), .B2(new_n833_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n879_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n881_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G113gat), .B1(new_n888_), .B2(new_n409_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n886_), .A2(new_n590_), .A3(new_n760_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1340gat));
  NAND2_X1  g690(.A1(new_n862_), .A2(new_n863_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n373_), .B1(new_n892_), .B2(new_n882_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n829_), .A2(new_n833_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n878_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n895_), .A2(KEYINPUT59), .B1(new_n877_), .B2(new_n880_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n345_), .A2(G120gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n886_), .B1(KEYINPUT60), .B2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n898_), .A3(new_n344_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G120gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(KEYINPUT60), .B2(new_n898_), .ZN(G1341gat));
  OAI21_X1  g700(.A(new_n587_), .B1(new_n895_), .B2(new_n718_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n902_), .A2(KEYINPUT117), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(KEYINPUT117), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n373_), .A2(G127gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT118), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n903_), .A2(new_n904_), .B1(new_n896_), .B2(new_n906_), .ZN(G1342gat));
  AOI21_X1  g706(.A(new_n585_), .B1(new_n896_), .B2(new_n802_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n895_), .A2(G134gat), .A3(new_n300_), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT119), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(G134gat), .B1(new_n888_), .B2(new_n308_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n912_));
  INV_X1    g711(.A(new_n909_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n911_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n914_), .ZN(G1343gat));
  NOR4_X1   g714(.A1(new_n734_), .A2(new_n483_), .A3(new_n687_), .A4(new_n648_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n884_), .A2(new_n684_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n834_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n760_), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT120), .B(G141gat), .Z(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1344gat));
  NAND2_X1  g721(.A1(new_n919_), .A2(new_n344_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT121), .B(G148gat), .Z(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1345gat));
  AOI21_X1  g724(.A(KEYINPUT122), .B1(new_n919_), .B2(new_n377_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n885_), .A2(new_n927_), .A3(new_n718_), .A4(new_n917_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT61), .B1(new_n926_), .B2(new_n928_), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n377_), .B(new_n916_), .C1(new_n893_), .C2(new_n894_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n927_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n919_), .A2(KEYINPUT122), .A3(new_n377_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n929_), .A2(G155gat), .A3(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(G155gat), .B1(new_n929_), .B2(new_n934_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1346gat));
  INV_X1    g736(.A(new_n919_), .ZN(new_n938_));
  OAI21_X1  g737(.A(G162gat), .B1(new_n938_), .B2(new_n308_), .ZN(new_n939_));
  OR2_X1    g738(.A1(new_n300_), .A2(G162gat), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n938_), .B2(new_n940_), .ZN(G1347gat));
  INV_X1    g740(.A(new_n877_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n734_), .A2(new_n483_), .A3(new_n634_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n760_), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n946_));
  AND3_X1   g745(.A1(new_n945_), .A2(new_n946_), .A3(G169gat), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n946_), .B1(new_n945_), .B2(G169gat), .ZN(new_n948_));
  INV_X1    g747(.A(new_n944_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n760_), .A2(new_n512_), .ZN(new_n950_));
  XOR2_X1   g749(.A(new_n950_), .B(KEYINPUT123), .Z(new_n951_));
  OAI22_X1  g750(.A1(new_n947_), .A2(new_n948_), .B1(new_n949_), .B2(new_n951_), .ZN(G1348gat));
  AOI21_X1  g751(.A(G176gat), .B1(new_n944_), .B2(new_n344_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n885_), .A2(new_n652_), .ZN(new_n954_));
  AND4_X1   g753(.A1(G176gat), .A2(new_n344_), .A3(new_n734_), .A4(new_n634_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n953_), .B1(new_n954_), .B2(new_n955_), .ZN(G1349gat));
  NAND4_X1  g755(.A1(new_n954_), .A2(new_n734_), .A3(new_n634_), .A4(new_n377_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n684_), .B1(new_n539_), .B2(new_n525_), .ZN(new_n958_));
  AOI22_X1  g757(.A1(new_n957_), .A2(new_n502_), .B1(new_n944_), .B2(new_n958_), .ZN(G1350gat));
  OAI21_X1  g758(.A(G190gat), .B1(new_n949_), .B2(new_n308_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n944_), .A2(new_n521_), .A3(new_n306_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1351gat));
  NAND2_X1  g761(.A1(new_n918_), .A2(new_n834_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n650_), .A2(new_n649_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n734_), .B1(new_n964_), .B2(KEYINPUT124), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n965_), .B1(KEYINPUT124), .B2(new_n964_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n963_), .A2(new_n966_), .ZN(new_n967_));
  INV_X1    g766(.A(new_n967_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(new_n760_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g769(.A1(new_n967_), .A2(new_n345_), .ZN(new_n971_));
  XOR2_X1   g770(.A(KEYINPUT125), .B(G204gat), .Z(new_n972_));
  XNOR2_X1  g771(.A(new_n971_), .B(new_n972_), .ZN(G1353gat));
  NAND2_X1  g772(.A1(new_n968_), .A2(new_n373_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(KEYINPUT63), .B(G211gat), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n974_), .A2(new_n975_), .ZN(new_n976_));
  INV_X1    g775(.A(KEYINPUT63), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n974_), .A2(new_n977_), .A3(new_n451_), .ZN(new_n978_));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n978_), .A2(new_n979_), .ZN(new_n980_));
  NAND4_X1  g779(.A1(new_n974_), .A2(KEYINPUT126), .A3(new_n977_), .A4(new_n451_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n976_), .B1(new_n980_), .B2(new_n981_), .ZN(G1354gat));
  NOR3_X1   g781(.A1(new_n967_), .A2(new_n453_), .A3(new_n308_), .ZN(new_n983_));
  AOI21_X1  g782(.A(KEYINPUT127), .B1(new_n968_), .B2(new_n306_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n984_), .A2(G218gat), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n968_), .A2(KEYINPUT127), .A3(new_n306_), .ZN(new_n986_));
  AOI21_X1  g785(.A(new_n983_), .B1(new_n985_), .B2(new_n986_), .ZN(G1355gat));
endmodule


