//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_, new_n958_;
  XNOR2_X1  g000(.A(G1gat), .B(G8gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT77), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT76), .B(G1gat), .ZN(new_n204_));
  INV_X1    g003(.A(G8gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n203_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n203_), .A2(new_n208_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G231gat), .A2(G233gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT70), .B(G71gat), .ZN(new_n214_));
  INV_X1    g013(.A(G78gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G57gat), .B(G64gat), .Z(new_n217_));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT71), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT71), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n216_), .A2(new_n222_), .A3(new_n219_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n217_), .A2(new_n218_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n221_), .A2(new_n225_), .A3(new_n223_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n213_), .B(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT72), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n221_), .A2(new_n225_), .A3(new_n223_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n225_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n213_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT72), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n238_));
  XNOR2_X1  g037(.A(G127gat), .B(G155gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G183gat), .B(G211gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n242_), .A2(KEYINPUT17), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n231_), .A2(new_n237_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n242_), .A2(KEYINPUT17), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n230_), .A2(new_n243_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G230gat), .A2(G233gat), .ZN(new_n254_));
  INV_X1    g053(.A(G106gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT10), .B(G99gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(G99gat), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n259_), .A2(KEYINPUT10), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(KEYINPUT10), .ZN(new_n261_));
  NOR3_X1   g060(.A1(new_n260_), .A2(new_n261_), .A3(KEYINPUT64), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n255_), .B1(new_n258_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(G85gat), .ZN(new_n264_));
  INV_X1    g063(.A(G92gat), .ZN(new_n265_));
  OR3_X1    g064(.A1(new_n264_), .A2(new_n265_), .A3(KEYINPUT9), .ZN(new_n266_));
  XOR2_X1   g065(.A(G85gat), .B(G92gat), .Z(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT9), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n263_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G99gat), .A2(G106gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(KEYINPUT6), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(KEYINPUT65), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n270_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(KEYINPUT65), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(KEYINPUT6), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(G99gat), .A4(G106gat), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n275_), .A2(KEYINPUT66), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT66), .B1(new_n275_), .B2(new_n278_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n269_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NOR3_X1   g084(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT68), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT7), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(new_n259_), .A3(new_n255_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n290_), .A3(new_n284_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n287_), .A2(new_n275_), .A3(new_n278_), .A4(new_n291_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n292_), .A2(KEYINPUT69), .A3(new_n267_), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT69), .B1(new_n292_), .B2(new_n267_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT8), .ZN(new_n295_));
  NOR3_X1   g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(KEYINPUT67), .B(KEYINPUT8), .Z(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n267_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n279_), .A2(new_n280_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n289_), .A2(new_n284_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n298_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n283_), .B1(new_n296_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT12), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n304_), .A2(KEYINPUT72), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n234_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n292_), .A2(new_n267_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n292_), .A2(KEYINPUT69), .A3(new_n267_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(KEYINPUT8), .A3(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n267_), .B(new_n297_), .C1(new_n281_), .C2(new_n300_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n282_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n305_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n229_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n304_), .ZN(new_n316_));
  AND4_X1   g115(.A1(new_n254_), .A2(new_n306_), .A3(new_n315_), .A4(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n229_), .B(new_n313_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n254_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT5), .B(G176gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G204gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G120gat), .B(G148gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n326_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n318_), .A2(new_n321_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT13), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n327_), .A2(KEYINPUT13), .A3(new_n329_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G29gat), .B(G36gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G50gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT73), .B(G43gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n211_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n211_), .A2(new_n339_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G229gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(KEYINPUT74), .B(KEYINPUT15), .Z(new_n346_));
  NAND3_X1  g145(.A1(new_n340_), .A2(new_n341_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n339_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n346_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n343_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n345_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G113gat), .B(G141gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G169gat), .B(G197gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT81), .B1(new_n352_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT81), .ZN(new_n358_));
  AOI211_X1 g157(.A(new_n358_), .B(new_n355_), .C1(new_n345_), .C2(new_n351_), .ZN(new_n359_));
  OAI22_X1  g158(.A1(new_n357_), .A2(new_n359_), .B1(new_n356_), .B2(new_n352_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n335_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT22), .B(G169gat), .ZN(new_n363_));
  INV_X1    g162(.A(G176gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT83), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367_));
  INV_X1    g166(.A(G183gat), .ZN(new_n368_));
  INV_X1    g167(.A(G190gat), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT23), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT23), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(G183gat), .A3(G190gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n369_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n363_), .A2(new_n376_), .A3(new_n364_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n366_), .A2(new_n367_), .A3(new_n375_), .A4(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n372_), .A2(KEYINPUT82), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n380_), .A2(new_n371_), .A3(G183gat), .A4(G190gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n370_), .A3(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT25), .B(G183gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT26), .B(G190gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n386_), .A2(KEYINPUT24), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(KEYINPUT24), .A3(new_n367_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n382_), .A2(new_n385_), .A3(new_n387_), .A4(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n378_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT30), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT84), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(KEYINPUT84), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(G15gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(G43gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G71gat), .B(G99gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  MUX2_X1   g198(.A(new_n392_), .B(new_n393_), .S(new_n399_), .Z(new_n400_));
  XNOR2_X1  g199(.A(G127gat), .B(G134gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G113gat), .B(G120gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n400_), .B(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(KEYINPUT99), .B(KEYINPUT0), .Z(new_n407_));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G57gat), .B(G85gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT100), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT86), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G155gat), .A2(G162gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT89), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT89), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n420_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT3), .ZN(new_n423_));
  NOR4_X1   g222(.A1(new_n423_), .A2(KEYINPUT87), .A3(G141gat), .A4(G148gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G141gat), .A2(G148gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT87), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT3), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n422_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT90), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n428_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(G141gat), .ZN(new_n434_));
  INV_X1    g233(.A(G148gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n426_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n423_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT3), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n437_), .A2(new_n438_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n429_), .B(KEYINPUT88), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT90), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n417_), .B1(new_n433_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n415_), .A2(KEYINPUT1), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n415_), .A2(KEYINPUT1), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n414_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n425_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G141gat), .A2(G148gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n442_), .A2(new_n403_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n403_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n432_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n439_), .A2(KEYINPUT90), .A3(new_n440_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n416_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n448_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n450_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT98), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n449_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n442_), .A2(new_n448_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(KEYINPUT98), .A3(new_n450_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G225gat), .A2(G233gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n412_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n461_), .ZN(new_n463_));
  AOI211_X1 g262(.A(KEYINPUT100), .B(new_n463_), .C1(new_n457_), .C2(new_n459_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(KEYINPUT4), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n455_), .A2(KEYINPUT4), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n468_));
  AOI211_X1 g267(.A(KEYINPUT105), .B(new_n411_), .C1(new_n465_), .C2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT105), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n457_), .A2(new_n459_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT100), .B1(new_n471_), .B2(new_n463_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n460_), .A2(new_n412_), .A3(new_n461_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n468_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n411_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n470_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n469_), .A2(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n468_), .A2(new_n472_), .A3(new_n411_), .A4(new_n473_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT104), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT104), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n465_), .A2(new_n480_), .A3(new_n411_), .A4(new_n468_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G197gat), .B(G204gat), .Z(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT21), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G197gat), .B(G204gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT21), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(G211gat), .A2(G218gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT93), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G211gat), .A2(G218gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n490_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT93), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n484_), .A2(new_n487_), .A3(new_n491_), .A4(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n491_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n489_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n496_));
  OAI211_X1 g295(.A(KEYINPUT21), .B(new_n483_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n365_), .A2(new_n367_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n499_), .B1(new_n382_), .B2(new_n374_), .ZN(new_n500_));
  AND4_X1   g299(.A1(new_n385_), .A2(new_n387_), .A3(new_n388_), .A4(new_n373_), .ZN(new_n501_));
  OR3_X1    g300(.A1(new_n498_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G226gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n390_), .A2(new_n498_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n502_), .A2(KEYINPUT20), .A3(new_n505_), .A4(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n498_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n378_), .A2(new_n389_), .A3(new_n494_), .A4(new_n497_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(KEYINPUT20), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n511_));
  INV_X1    g310(.A(new_n505_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n511_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n507_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G64gat), .B(G92gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(G8gat), .B(G36gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n515_), .A2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n520_), .B(new_n507_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(KEYINPUT97), .A3(new_n523_), .ZN(new_n524_));
  OR3_X1    g323(.A1(new_n515_), .A2(KEYINPUT97), .A3(new_n521_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT27), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n502_), .A2(new_n506_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT103), .B(KEYINPUT20), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n512_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n530_), .B1(new_n512_), .B2(new_n510_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n521_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(KEYINPUT27), .A3(new_n523_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n527_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n458_), .A2(KEYINPUT29), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT29), .B1(new_n453_), .B2(new_n454_), .ZN(new_n539_));
  INV_X1    g338(.A(G228gat), .ZN(new_n540_));
  INV_X1    g339(.A(G233gat), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n539_), .A2(new_n498_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n543_), .B1(new_n539_), .B2(new_n498_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n538_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n546_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(new_n544_), .A3(new_n537_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n536_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n549_), .A3(new_n536_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G78gat), .B(G106gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(G50gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT91), .B(G22gat), .Z(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n556_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n552_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n558_), .B1(new_n559_), .B2(new_n550_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n477_), .A2(new_n482_), .A3(new_n534_), .A4(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT106), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n479_), .A2(new_n481_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n565_), .A2(new_n469_), .A3(new_n476_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n566_), .A2(KEYINPUT106), .A3(new_n561_), .A4(new_n534_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n474_), .A2(new_n475_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT105), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n474_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n479_), .A4(new_n481_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n520_), .A2(KEYINPUT32), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n531_), .A2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n515_), .A2(new_n574_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n572_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n478_), .A2(KEYINPUT101), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT33), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n466_), .A2(new_n461_), .A3(new_n467_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n471_), .B(KEYINPUT102), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n475_), .B(new_n580_), .C1(new_n581_), .C2(new_n461_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT33), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n478_), .A2(KEYINPUT101), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n524_), .A2(new_n525_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n579_), .A2(new_n582_), .A3(new_n584_), .A4(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n561_), .B1(new_n577_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n406_), .B1(new_n568_), .B2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n561_), .A2(new_n406_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n534_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n590_), .A2(new_n572_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n588_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT34), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n303_), .A2(new_n339_), .A3(new_n346_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n348_), .B1(new_n313_), .B2(new_n349_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT75), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n602_), .A2(new_n603_), .A3(new_n598_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n605_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n607_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT75), .B1(new_n609_), .B2(new_n604_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G190gat), .B(G218gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n611_), .B(new_n612_), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT36), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n608_), .A2(new_n610_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT107), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n605_), .A2(new_n617_), .A3(new_n613_), .A4(new_n607_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n615_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n616_), .B1(new_n615_), .B2(new_n618_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n594_), .A2(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n622_), .A2(KEYINPUT108), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(KEYINPUT108), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n253_), .B(new_n362_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G1gat), .B1(new_n625_), .B2(new_n566_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT80), .B1(new_n248_), .B2(new_n251_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT80), .ZN(new_n628_));
  AOI211_X1 g427(.A(new_n628_), .B(new_n250_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n615_), .A2(new_n618_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n631_), .A2(KEYINPUT37), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n614_), .B1(new_n609_), .B2(new_n604_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n618_), .A2(KEYINPUT37), .A3(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n630_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(new_n361_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n594_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n572_), .A3(new_n204_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT38), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n626_), .A2(new_n641_), .ZN(G1324gat));
  NAND3_X1  g441(.A1(new_n639_), .A2(new_n205_), .A3(new_n591_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n644_), .B(G8gat), .C1(new_n625_), .C2(new_n534_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n622_), .B(KEYINPUT108), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n647_), .A2(new_n253_), .A3(new_n362_), .A4(new_n591_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n644_), .B1(new_n648_), .B2(G8gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n643_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT40), .B(new_n643_), .C1(new_n646_), .C2(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1325gat));
  INV_X1    g453(.A(new_n406_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n647_), .A2(new_n253_), .A3(new_n362_), .A4(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G15gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT109), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT109), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n656_), .A2(new_n659_), .A3(G15gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n639_), .A2(new_n395_), .A3(new_n655_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n658_), .A2(KEYINPUT41), .A3(new_n660_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n663_), .A2(new_n664_), .A3(new_n665_), .ZN(G1326gat));
  INV_X1    g465(.A(new_n561_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G22gat), .B1(new_n625_), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT42), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n667_), .A2(G22gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n638_), .B2(new_n670_), .ZN(G1327gat));
  AOI22_X1  g470(.A1(new_n477_), .A2(new_n482_), .B1(new_n531_), .B2(new_n574_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n579_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n673_));
  AOI22_X1  g472(.A1(new_n672_), .A2(new_n576_), .B1(new_n673_), .B2(new_n582_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n564_), .B(new_n567_), .C1(new_n674_), .C2(new_n561_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n592_), .B1(new_n675_), .B2(new_n406_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(new_n621_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n630_), .A2(new_n361_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(G29gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(new_n572_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT111), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n682_), .B(new_n683_), .C1(new_n676_), .C2(new_n635_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n635_), .B1(new_n588_), .B2(new_n593_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT43), .B1(new_n685_), .B2(KEYINPUT111), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n678_), .B(KEYINPUT110), .Z(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n684_), .A2(new_n686_), .A3(new_n687_), .A4(KEYINPUT44), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n572_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n693_), .A2(KEYINPUT112), .A3(G29gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT112), .B1(new_n693_), .B2(G29gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n681_), .B1(new_n694_), .B2(new_n695_), .ZN(G1328gat));
  INV_X1    g495(.A(G36gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n679_), .A2(new_n697_), .A3(new_n591_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT45), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n690_), .A2(new_n591_), .A3(new_n691_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G36gat), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n699_), .A2(KEYINPUT46), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  AOI21_X1  g505(.A(G43gat), .B1(new_n679_), .B2(new_n655_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT113), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n690_), .A2(G43gat), .A3(new_n655_), .A4(new_n691_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT47), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n713_), .A3(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1330gat));
  AOI21_X1  g514(.A(G50gat), .B1(new_n679_), .B2(new_n561_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n561_), .A2(G50gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n692_), .B2(new_n717_), .ZN(G1331gat));
  NOR2_X1   g517(.A1(new_n636_), .A2(new_n335_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT114), .ZN(new_n720_));
  INV_X1    g519(.A(new_n360_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(new_n594_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G57gat), .B1(new_n723_), .B2(new_n572_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n334_), .A2(new_n721_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n647_), .A2(new_n630_), .A3(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(G57gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n572_), .B2(KEYINPUT115), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(KEYINPUT115), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n724_), .B1(new_n730_), .B2(new_n731_), .ZN(G1332gat));
  INV_X1    g531(.A(G64gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n723_), .A2(new_n733_), .A3(new_n591_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n727_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n733_), .B1(new_n735_), .B2(new_n591_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n736_), .A2(new_n737_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n734_), .B1(new_n739_), .B2(new_n740_), .ZN(G1333gat));
  INV_X1    g540(.A(G71gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n723_), .A2(new_n742_), .A3(new_n655_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n735_), .B2(new_n655_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT49), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n744_), .A2(new_n745_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n743_), .B1(new_n747_), .B2(new_n748_), .ZN(G1334gat));
  OAI21_X1  g548(.A(G78gat), .B1(new_n727_), .B2(new_n667_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT50), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n723_), .A2(new_n215_), .A3(new_n561_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n630_), .A2(new_n725_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n677_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G85gat), .B1(new_n755_), .B2(new_n572_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n684_), .A2(new_n686_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n754_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n566_), .A2(new_n264_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(G1336gat));
  AOI21_X1  g560(.A(G92gat), .B1(new_n755_), .B2(new_n591_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n534_), .A2(new_n265_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n759_), .B2(new_n763_), .ZN(G1337gat));
  OAI21_X1  g563(.A(G99gat), .B1(new_n758_), .B2(new_n406_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n755_), .B(new_n655_), .C1(new_n258_), .C2(new_n262_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n684_), .A2(new_n686_), .A3(new_n561_), .A4(new_n754_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(new_n771_), .A3(G106gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(G106gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n770_), .A2(G106gat), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT117), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n770_), .A2(new_n771_), .A3(G106gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(KEYINPUT52), .A3(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n755_), .A2(new_n255_), .A3(new_n561_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n774_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT53), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n774_), .A2(new_n778_), .A3(new_n782_), .A4(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1339gat));
  INV_X1    g583(.A(KEYINPUT122), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n360_), .A2(new_n329_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n306_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n320_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n317_), .B1(KEYINPUT55), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n787_), .A2(new_n790_), .A3(new_n320_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n326_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT56), .B(new_n326_), .C1(new_n789_), .C2(new_n791_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n786_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n347_), .A2(new_n797_), .A3(new_n350_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n344_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  OR2_X1    g599(.A1(new_n342_), .A2(new_n344_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n355_), .A3(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n621_), .B1(new_n796_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n621_), .B(KEYINPUT119), .C1(new_n796_), .C2(new_n804_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT120), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n788_), .A2(KEYINPUT55), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n318_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n791_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n328_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n811_), .B1(new_n815_), .B2(KEYINPUT56), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n792_), .A2(KEYINPUT120), .A3(new_n793_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n795_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n803_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(new_n329_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n632_), .A2(new_n634_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n818_), .A2(KEYINPUT58), .A3(new_n820_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n823_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n809_), .A2(new_n810_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n805_), .A2(new_n810_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n818_), .A2(KEYINPUT58), .A3(new_n820_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT58), .B1(new_n818_), .B2(new_n820_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n635_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n830_), .B1(new_n833_), .B2(KEYINPUT121), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n253_), .B1(new_n828_), .B2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n630_), .A2(new_n635_), .A3(new_n721_), .A4(new_n335_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT54), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n785_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n807_), .A2(new_n810_), .A3(new_n808_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n833_), .B2(KEYINPUT121), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n829_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n252_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(KEYINPUT122), .A3(new_n837_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n590_), .A2(new_n566_), .A3(new_n591_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n839_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(new_n721_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(G113gat), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n807_), .A2(new_n810_), .A3(new_n808_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n833_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n826_), .A2(new_n840_), .A3(KEYINPUT123), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n829_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n630_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n838_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n845_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  AOI211_X1 g657(.A(new_n721_), .B(new_n858_), .C1(KEYINPUT59), .C2(new_n846_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n848_), .B1(new_n859_), .B2(G113gat), .ZN(G1340gat));
  AOI211_X1 g659(.A(new_n335_), .B(new_n858_), .C1(KEYINPUT59), .C2(new_n846_), .ZN(new_n861_));
  INV_X1    g660(.A(G120gat), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(KEYINPUT60), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n839_), .A2(new_n844_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n862_), .B1(new_n335_), .B2(KEYINPUT60), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n845_), .A3(new_n865_), .ZN(new_n866_));
  OAI22_X1  g665(.A1(new_n861_), .A2(new_n862_), .B1(new_n863_), .B2(new_n866_), .ZN(G1341gat));
  INV_X1    g666(.A(G127gat), .ZN(new_n868_));
  AOI211_X1 g667(.A(new_n868_), .B(new_n858_), .C1(KEYINPUT59), .C2(new_n846_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n864_), .A2(new_n630_), .A3(new_n845_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n869_), .A2(new_n253_), .B1(new_n868_), .B2(new_n870_), .ZN(G1342gat));
  NOR2_X1   g670(.A1(new_n846_), .A2(new_n621_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(G134gat), .ZN(new_n873_));
  AOI211_X1 g672(.A(new_n635_), .B(new_n858_), .C1(KEYINPUT59), .C2(new_n846_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(G134gat), .ZN(G1343gat));
  NAND4_X1  g674(.A1(new_n839_), .A2(new_n572_), .A3(new_n561_), .A4(new_n844_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n591_), .A2(new_n655_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G141gat), .B1(new_n879_), .B2(new_n721_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n876_), .A2(new_n878_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(new_n434_), .A3(new_n360_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1344gat));
  OAI21_X1  g682(.A(G148gat), .B1(new_n879_), .B2(new_n335_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n881_), .A2(new_n435_), .A3(new_n334_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1345gat));
  XNOR2_X1  g685(.A(KEYINPUT61), .B(G155gat), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n881_), .B2(new_n630_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n887_), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n876_), .A2(new_n854_), .A3(new_n878_), .A4(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1346gat));
  INV_X1    g690(.A(G162gat), .ZN(new_n892_));
  NOR4_X1   g691(.A1(new_n876_), .A2(new_n892_), .A3(new_n635_), .A4(new_n878_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n621_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n881_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n892_), .B2(new_n895_), .ZN(G1347gat));
  NAND2_X1  g695(.A1(new_n360_), .A2(new_n363_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT125), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n853_), .A2(new_n854_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n590_), .B1(new_n900_), .B2(new_n837_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n572_), .A2(new_n534_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n899_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n902_), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n855_), .A2(KEYINPUT124), .A3(new_n590_), .A4(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n898_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n901_), .A2(new_n360_), .A3(new_n902_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n907_), .A2(new_n908_), .A3(G169gat), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n908_), .B1(new_n907_), .B2(G169gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n906_), .B1(new_n910_), .B2(new_n911_), .ZN(G1348gat));
  OAI21_X1  g711(.A(new_n334_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n864_), .A2(new_n667_), .ZN(new_n914_));
  NOR4_X1   g713(.A1(new_n904_), .A2(new_n335_), .A3(new_n364_), .A4(new_n406_), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n913_), .A2(new_n364_), .B1(new_n914_), .B2(new_n915_), .ZN(G1349gat));
  NOR2_X1   g715(.A1(new_n252_), .A2(new_n383_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n854_), .A2(new_n406_), .A3(new_n904_), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n839_), .A2(new_n667_), .A3(new_n844_), .A4(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n368_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n918_), .A2(KEYINPUT126), .A3(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923_));
  INV_X1    g722(.A(new_n917_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n826_), .A2(new_n840_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n830_), .B1(new_n925_), .B2(new_n849_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n630_), .B1(new_n926_), .B2(new_n852_), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n589_), .B(new_n902_), .C1(new_n927_), .C2(new_n838_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(KEYINPUT124), .ZN(new_n929_));
  AND3_X1   g728(.A1(new_n826_), .A2(new_n840_), .A3(KEYINPUT123), .ZN(new_n930_));
  AOI21_X1  g729(.A(KEYINPUT123), .B1(new_n826_), .B2(new_n840_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n930_), .A2(new_n931_), .A3(new_n830_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n837_), .B1(new_n932_), .B2(new_n630_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n933_), .A2(new_n899_), .A3(new_n589_), .A4(new_n902_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n924_), .B1(new_n929_), .B2(new_n934_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n920_), .A2(new_n368_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n923_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n922_), .A2(new_n937_), .ZN(G1350gat));
  OAI211_X1 g737(.A(new_n894_), .B(new_n384_), .C1(new_n903_), .C2(new_n905_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n635_), .B1(new_n929_), .B2(new_n934_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n369_), .B2(new_n940_), .ZN(G1351gat));
  NAND4_X1  g740(.A1(new_n839_), .A2(new_n561_), .A3(new_n844_), .A4(new_n902_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n942_), .A2(new_n721_), .A3(new_n655_), .ZN(new_n943_));
  INV_X1    g742(.A(G197gat), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n943_), .B(new_n944_), .ZN(G1352gat));
  NOR3_X1   g744(.A1(new_n942_), .A2(new_n335_), .A3(new_n655_), .ZN(new_n946_));
  INV_X1    g745(.A(G204gat), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n946_), .B(new_n947_), .ZN(G1353gat));
  XNOR2_X1  g747(.A(KEYINPUT63), .B(G211gat), .ZN(new_n949_));
  NOR4_X1   g748(.A1(new_n942_), .A2(new_n252_), .A3(new_n655_), .A4(new_n949_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n942_), .A2(new_n655_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(new_n253_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n950_), .B1(new_n952_), .B2(new_n953_), .ZN(G1354gat));
  NAND2_X1  g753(.A1(new_n951_), .A2(new_n894_), .ZN(new_n955_));
  INV_X1    g754(.A(G218gat), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n824_), .A2(G218gat), .ZN(new_n957_));
  XOR2_X1   g756(.A(new_n957_), .B(KEYINPUT127), .Z(new_n958_));
  AOI22_X1  g757(.A1(new_n955_), .A2(new_n956_), .B1(new_n951_), .B2(new_n958_), .ZN(G1355gat));
endmodule


