//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT94), .ZN(new_n204_));
  OR3_X1    g003(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n205_));
  INV_X1    g004(.A(G183gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT78), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT78), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G183gat), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n207_), .A2(new_n209_), .A3(KEYINPUT25), .ZN(new_n210_));
  INV_X1    g009(.A(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT26), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT26), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G190gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT25), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(G183gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n205_), .B1(new_n210_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT80), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT23), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(KEYINPUT23), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT79), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n227_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G169gat), .ZN(new_n232_));
  INV_X1    g031(.A(G176gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n234_), .A2(KEYINPUT79), .A3(KEYINPUT24), .A4(new_n228_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n218_), .A2(new_n226_), .A3(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(new_n232_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n219_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n221_), .A2(new_n222_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n242_), .B1(new_n243_), .B2(KEYINPUT23), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT78), .B(G183gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(new_n211_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n239_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT81), .B1(new_n237_), .B2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G211gat), .B(G218gat), .Z(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT21), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT91), .ZN(new_n251_));
  INV_X1    g050(.A(G204gat), .ZN(new_n252_));
  INV_X1    g051(.A(G197gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT89), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT89), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G197gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n252_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(G197gat), .A2(G204gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n251_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n258_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT89), .B(G197gat), .ZN(new_n261_));
  OAI211_X1 g060(.A(KEYINPUT91), .B(new_n260_), .C1(new_n261_), .C2(new_n252_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n250_), .B1(new_n259_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n254_), .A2(new_n256_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n258_), .B1(new_n264_), .B2(G204gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT90), .B1(new_n265_), .B2(KEYINPUT21), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT90), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT21), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n267_), .B(new_n268_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n261_), .A2(new_n252_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n268_), .B1(G197gat), .B2(G204gat), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n249_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n263_), .B1(new_n270_), .B2(new_n273_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n231_), .A2(new_n235_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n245_), .A2(KEYINPUT25), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n212_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(KEYINPUT80), .A2(G183gat), .A3(G190gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT80), .B1(G183gat), .B2(G190gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n240_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n224_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n275_), .A2(new_n278_), .A3(new_n282_), .A4(new_n205_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n239_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n279_), .A2(new_n280_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n241_), .B1(new_n285_), .B2(new_n240_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n245_), .A2(new_n211_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n284_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT81), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n283_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n248_), .A2(new_n274_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT96), .ZN(new_n292_));
  NOR2_X1   g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n281_), .B2(new_n224_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n292_), .B1(new_n294_), .B2(new_n239_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n293_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n296_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n297_), .A2(KEYINPUT96), .A3(new_n284_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n212_), .A2(new_n214_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n206_), .A2(KEYINPUT25), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT95), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n216_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n301_), .B1(new_n216_), .B2(new_n300_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n299_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n205_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n286_), .A2(new_n305_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n295_), .A2(new_n298_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT20), .B1(new_n274_), .B2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n204_), .B1(new_n291_), .B2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G8gat), .B(G36gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(G64gat), .B(G92gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n269_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n260_), .B1(new_n261_), .B2(new_n252_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n267_), .B1(new_n317_), .B2(new_n268_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n273_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n263_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n283_), .A2(new_n289_), .A3(new_n288_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n289_), .B1(new_n283_), .B2(new_n288_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n274_), .A2(new_n307_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT20), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n203_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n309_), .A2(new_n315_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT27), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n314_), .B(KEYINPUT104), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n306_), .A2(new_n304_), .ZN(new_n333_));
  NOR3_X1   g132(.A1(new_n294_), .A2(new_n292_), .A3(new_n239_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT96), .B1(new_n297_), .B2(new_n284_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n326_), .B1(new_n321_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n204_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n248_), .A2(new_n274_), .A3(new_n290_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT101), .B(KEYINPUT20), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n306_), .A2(new_n304_), .B1(new_n297_), .B2(new_n284_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n341_), .B1(new_n274_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n324_), .A2(new_n343_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n340_), .A2(KEYINPUT102), .B1(new_n344_), .B2(new_n203_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT102), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n337_), .A2(new_n339_), .A3(new_n346_), .A4(new_n338_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n332_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT105), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n330_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n340_), .A2(KEYINPUT102), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n344_), .A2(new_n203_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n347_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n331_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT105), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n350_), .A2(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n324_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n338_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n357_), .A2(new_n358_), .A3(new_n314_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n315_), .B1(new_n309_), .B2(new_n328_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT106), .B(KEYINPUT27), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n356_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G71gat), .B(G99gat), .ZN(new_n366_));
  INV_X1    g165(.A(G43gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT30), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n370_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n372_), .B(G15gat), .Z(new_n373_));
  NAND3_X1  g172(.A1(new_n248_), .A2(new_n290_), .A3(new_n369_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(KEYINPUT85), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT84), .ZN(new_n378_));
  INV_X1    g177(.A(G134gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G127gat), .ZN(new_n380_));
  INV_X1    g179(.A(G127gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G134gat), .ZN(new_n382_));
  INV_X1    g181(.A(G113gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n383_), .A2(G120gat), .ZN(new_n384_));
  INV_X1    g183(.A(G120gat), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n385_), .A2(G113gat), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n380_), .B(new_n382_), .C1(new_n384_), .C2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n380_), .A2(new_n382_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G113gat), .B(G120gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n387_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n378_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n387_), .A2(new_n390_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n391_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n387_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(KEYINPUT84), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(KEYINPUT31), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(KEYINPUT31), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n375_), .A2(new_n377_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n377_), .B2(new_n375_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(G141gat), .A2(G148gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G141gat), .A2(G148gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(G155gat), .A2(G162gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT1), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n413_), .A2(KEYINPUT1), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n409_), .B(new_n410_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT2), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n410_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT86), .B1(new_n409_), .B2(KEYINPUT3), .ZN(new_n423_));
  OR4_X1    g222(.A1(KEYINPUT86), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n412_), .A2(new_n413_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n417_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n394_), .A2(new_n399_), .A3(new_n427_), .ZN(new_n428_));
  OAI221_X1 g227(.A(new_n417_), .B1(new_n425_), .B2(new_n426_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(KEYINPUT4), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n394_), .A2(new_n399_), .A3(new_n427_), .A4(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G225gat), .A2(G233gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT98), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n428_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G1gat), .B(G29gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT99), .B(G85gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT0), .B(G57gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n437_), .A2(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n428_), .A2(KEYINPUT4), .A3(new_n429_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n432_), .A2(new_n434_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n436_), .B(new_n442_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G78gat), .B(G106gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n427_), .A2(KEYINPUT29), .ZN(new_n451_));
  XOR2_X1   g250(.A(KEYINPUT87), .B(G228gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT88), .B(G233gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n321_), .A2(new_n451_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n455_), .B1(new_n321_), .B2(new_n451_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n450_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT93), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n321_), .A2(new_n451_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n454_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n450_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n456_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT92), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT93), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n466_), .B(new_n450_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT92), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n462_), .A2(new_n468_), .A3(new_n456_), .A4(new_n463_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n460_), .A2(new_n465_), .A3(new_n467_), .A4(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G22gat), .B(G50gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n427_), .A2(KEYINPUT29), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT28), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n473_), .A2(new_n474_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n472_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n477_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(new_n475_), .A3(new_n471_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n470_), .A2(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n459_), .A2(new_n464_), .A3(new_n480_), .A4(new_n478_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n407_), .A2(new_n449_), .A3(new_n482_), .A4(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n365_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT103), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n315_), .A2(KEYINPUT32), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n309_), .A2(new_n328_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n447_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n442_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n487_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n486_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT100), .B1(new_n447_), .B2(new_n494_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n428_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n432_), .A2(new_n434_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n430_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT100), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(KEYINPUT33), .A4(new_n442_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n430_), .A2(new_n433_), .A3(new_n432_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n428_), .A2(new_n429_), .A3(new_n434_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n503_), .A2(new_n443_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n447_), .A2(new_n494_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n361_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n487_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n353_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n508_), .A2(KEYINPUT103), .A3(new_n448_), .A4(new_n488_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n493_), .A2(new_n506_), .A3(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n482_), .A2(new_n483_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n448_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(new_n356_), .A3(new_n364_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n407_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n485_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518_));
  INV_X1    g317(.A(G1gat), .ZN(new_n519_));
  INV_X1    g318(.A(G8gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT14), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G1gat), .B(G8gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G29gat), .B(G36gat), .Z(new_n525_));
  XOR2_X1   g324(.A(G43gat), .B(G50gat), .Z(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G29gat), .B(G36gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G43gat), .B(G50gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n524_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT76), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(G229gat), .A3(G233gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(KEYINPUT68), .B(KEYINPUT15), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n531_), .B(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n524_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538_));
  INV_X1    g337(.A(new_n531_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n537_), .B(new_n538_), .C1(new_n524_), .C2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n534_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G113gat), .B(G141gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G169gat), .B(G197gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n534_), .A2(new_n540_), .A3(new_n544_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n548_), .B(KEYINPUT77), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n517_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G230gat), .A2(G233gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n552_), .B(KEYINPUT64), .Z(new_n553_));
  XNOR2_X1  g352(.A(G85gat), .B(G92gat), .ZN(new_n554_));
  INV_X1    g353(.A(G92gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n554_), .B1(KEYINPUT9), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT65), .ZN(new_n557_));
  AND2_X1   g356(.A1(G85gat), .A2(G92gat), .ZN(new_n558_));
  NOR2_X1   g357(.A1(G85gat), .A2(G92gat), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT9), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n557_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(G85gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n555_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G85gat), .A2(G92gat), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n565_), .A2(new_n566_), .B1(new_n561_), .B2(G92gat), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n558_), .A2(new_n559_), .A3(KEYINPUT9), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT65), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(KEYINPUT10), .B(G99gat), .Z(new_n570_));
  INV_X1    g369(.A(G106gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT6), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT6), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(G99gat), .A3(G106gat), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n570_), .A2(new_n571_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n563_), .A2(new_n569_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT7), .ZN(new_n578_));
  INV_X1    g377(.A(G99gat), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n579_), .A3(new_n571_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT66), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n580_), .A2(KEYINPUT66), .A3(new_n581_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n573_), .A2(new_n575_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT8), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n554_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n560_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n588_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n577_), .A2(new_n590_), .A3(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G57gat), .B(G64gat), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT11), .ZN(new_n596_));
  XOR2_X1   g395(.A(G71gat), .B(G78gat), .Z(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n595_), .A2(KEYINPUT11), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n596_), .A2(new_n597_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n594_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n601_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n604_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n605_), .A2(new_n577_), .A3(new_n590_), .A4(new_n593_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n603_), .A2(KEYINPUT12), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT12), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n594_), .A2(new_n608_), .A3(new_n602_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n553_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n553_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT5), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n615_), .B(new_n616_), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n613_), .B(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT13), .Z(new_n619_));
  XOR2_X1   g418(.A(G127gat), .B(G155gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT16), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(KEYINPUT74), .A3(KEYINPUT17), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n625_), .B1(KEYINPUT17), .B2(new_n624_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT17), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT75), .B1(new_n623_), .B2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(KEYINPUT74), .B2(new_n624_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n524_), .B(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(new_n602_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n626_), .B1(new_n629_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n628_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT37), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT35), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n639_));
  NAND2_X1  g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n536_), .A2(new_n594_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT69), .ZN(new_n643_));
  AOI211_X1 g442(.A(new_n638_), .B(new_n641_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n594_), .A2(new_n539_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n642_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n642_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n638_), .B2(new_n641_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n648_), .B2(new_n644_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G190gat), .B(G218gat), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT70), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(G134gat), .B(G162gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(KEYINPUT36), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n649_), .A2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT71), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n654_), .B(KEYINPUT36), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT72), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n661_), .B(new_n646_), .C1(new_n644_), .C2(new_n648_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT73), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n637_), .B1(new_n658_), .B2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n646_), .B(new_n659_), .C1(new_n648_), .C2(new_n644_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n657_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(KEYINPUT37), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n619_), .B(new_n636_), .C1(new_n665_), .C2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n551_), .A2(new_n670_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n671_), .A2(G1gat), .A3(new_n449_), .ZN(new_n672_));
  XOR2_X1   g471(.A(KEYINPUT107), .B(KEYINPUT38), .Z(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n667_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n517_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n619_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n548_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n636_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n676_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G1gat), .B1(new_n681_), .B2(new_n449_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n672_), .A2(new_n673_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n674_), .A2(new_n682_), .A3(new_n683_), .ZN(G1324gat));
  NAND3_X1  g483(.A1(new_n676_), .A2(new_n365_), .A3(new_n680_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n685_), .A2(KEYINPUT108), .A3(G8gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT108), .B1(new_n685_), .B2(G8gat), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT39), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n686_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n688_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n551_), .A2(new_n520_), .A3(new_n365_), .A4(new_n670_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT40), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n689_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(new_n689_), .B2(new_n692_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1325gat));
  NOR3_X1   g495(.A1(new_n671_), .A2(G15gat), .A3(new_n516_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT109), .Z(new_n698_));
  OAI21_X1  g497(.A(G15gat), .B1(new_n681_), .B2(new_n516_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT41), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n699_), .A2(KEYINPUT41), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n698_), .A2(new_n700_), .A3(new_n701_), .ZN(G1326gat));
  OAI21_X1  g501(.A(G22gat), .B1(new_n681_), .B2(new_n511_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT42), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n511_), .A2(G22gat), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT110), .Z(new_n706_));
  OAI21_X1  g505(.A(new_n704_), .B1(new_n671_), .B2(new_n706_), .ZN(G1327gat));
  NAND2_X1  g506(.A1(new_n658_), .A2(new_n664_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n668_), .B1(new_n708_), .B2(KEYINPUT37), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n517_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n407_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n712_), .B(new_n709_), .C1(new_n713_), .C2(new_n485_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n677_), .A2(new_n678_), .A3(new_n636_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT44), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n363_), .B1(new_n350_), .B2(new_n355_), .ZN(new_n718_));
  AOI22_X1  g517(.A1(new_n513_), .A2(new_n718_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n719_), .A2(new_n407_), .B1(new_n365_), .B2(new_n484_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n712_), .B1(new_n720_), .B2(new_n709_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n714_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT44), .B(new_n716_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n716_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n711_), .B2(new_n714_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(KEYINPUT111), .A3(KEYINPUT44), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n717_), .B1(new_n725_), .B2(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(new_n448_), .ZN(new_n730_));
  INV_X1    g529(.A(G29gat), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n675_), .A2(new_n679_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT112), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n677_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n551_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n448_), .A2(new_n731_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT113), .ZN(new_n737_));
  OAI22_X1  g536(.A1(new_n730_), .A2(new_n731_), .B1(new_n735_), .B2(new_n737_), .ZN(G1328gat));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739_));
  INV_X1    g538(.A(G36gat), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n725_), .A2(new_n728_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n365_), .B1(new_n727_), .B2(KEYINPUT44), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n740_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n551_), .A2(new_n734_), .A3(new_n740_), .A4(new_n365_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT45), .Z(new_n746_));
  OAI21_X1  g545(.A(new_n739_), .B1(new_n744_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n746_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n742_), .B1(new_n725_), .B2(new_n728_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n748_), .B(KEYINPUT46), .C1(new_n740_), .C2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(G1329gat));
  NOR2_X1   g550(.A1(new_n516_), .A2(new_n367_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n753_), .B(new_n717_), .C1(new_n725_), .C2(new_n728_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n735_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G43gat), .B1(new_n755_), .B2(new_n407_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT47), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n729_), .A2(new_n752_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n759_));
  INV_X1    g558(.A(new_n756_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n757_), .A2(new_n761_), .ZN(G1330gat));
  INV_X1    g561(.A(new_n511_), .ZN(new_n763_));
  AOI21_X1  g562(.A(G50gat), .B1(new_n755_), .B2(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n763_), .A2(G50gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n729_), .B2(new_n765_), .ZN(G1331gat));
  NAND4_X1  g565(.A1(new_n676_), .A2(new_n550_), .A3(new_n677_), .A4(new_n636_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G57gat), .B1(new_n767_), .B2(new_n449_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n517_), .A2(new_n548_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n709_), .A2(new_n679_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n677_), .A3(new_n770_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n449_), .A2(G57gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(G1332gat));
  OAI21_X1  g572(.A(G64gat), .B1(new_n767_), .B2(new_n718_), .ZN(new_n774_));
  XOR2_X1   g573(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n775_));
  XNOR2_X1  g574(.A(new_n774_), .B(new_n775_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n718_), .A2(G64gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n771_), .B2(new_n777_), .ZN(G1333gat));
  OAI21_X1  g577(.A(G71gat), .B1(new_n767_), .B2(new_n516_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n516_), .A2(G71gat), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT116), .Z(new_n783_));
  OAI21_X1  g582(.A(new_n781_), .B1(new_n771_), .B2(new_n783_), .ZN(G1334gat));
  OAI21_X1  g583(.A(G78gat), .B1(new_n767_), .B2(new_n511_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT50), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n511_), .A2(G78gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n771_), .B2(new_n787_), .ZN(G1335gat));
  NAND3_X1  g587(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n715_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791_), .B2(new_n449_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n733_), .A2(new_n619_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n769_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(new_n564_), .A3(new_n448_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n792_), .A2(new_n796_), .ZN(G1336gat));
  OAI21_X1  g596(.A(G92gat), .B1(new_n791_), .B2(new_n718_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n555_), .A3(new_n365_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(G1337gat));
  NAND3_X1  g599(.A1(new_n795_), .A2(new_n407_), .A3(new_n570_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n791_), .A2(new_n516_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n579_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n803_), .B(new_n804_), .Z(G1338gat));
  OAI211_X1 g604(.A(new_n763_), .B(new_n790_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n715_), .A2(KEYINPUT119), .A3(new_n763_), .A4(new_n790_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n808_), .A2(KEYINPUT52), .A3(G106gat), .A4(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n763_), .A2(new_n571_), .ZN(new_n811_));
  OR3_X1    g610(.A1(new_n794_), .A2(KEYINPUT118), .A3(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT118), .B1(new_n794_), .B2(new_n811_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n810_), .A2(new_n814_), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n511_), .B(new_n789_), .C1(new_n711_), .C2(new_n714_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n571_), .B1(new_n816_), .B2(KEYINPUT119), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(new_n817_), .B2(new_n808_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT53), .B1(new_n815_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820_));
  INV_X1    g619(.A(new_n808_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n809_), .A2(G106gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n820_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n810_), .A4(new_n814_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n819_), .A2(new_n825_), .ZN(G1339gat));
  INV_X1    g625(.A(new_n617_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n613_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n548_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n607_), .A2(new_n609_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n611_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n607_), .A2(new_n553_), .A3(new_n609_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(KEYINPUT55), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n830_), .A2(new_n835_), .A3(new_n611_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n833_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n834_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n617_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n832_), .A2(KEYINPUT55), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n610_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n836_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT120), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n833_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(KEYINPUT56), .A3(new_n617_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n829_), .B1(new_n841_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n533_), .A2(new_n538_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n524_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n538_), .B1(new_n851_), .B2(new_n531_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n544_), .B1(new_n537_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n547_), .A2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n618_), .A2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n667_), .B1(new_n849_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT57), .B(new_n667_), .C1(new_n849_), .C2(new_n856_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n855_), .B1(new_n613_), .B2(new_n827_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT56), .B1(new_n847_), .B2(new_n617_), .ZN(new_n862_));
  AOI211_X1 g661(.A(new_n840_), .B(new_n827_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n861_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT58), .B(new_n861_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n709_), .A3(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n859_), .A2(new_n860_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n679_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n670_), .A2(new_n871_), .A3(new_n550_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT54), .B1(new_n669_), .B2(new_n549_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n763_), .B1(new_n870_), .B2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n718_), .A2(new_n448_), .A3(new_n407_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n875_), .A2(new_n383_), .A3(new_n548_), .A4(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n870_), .A2(new_n874_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n879_), .A2(KEYINPUT121), .A3(new_n511_), .A4(new_n877_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n875_), .A2(KEYINPUT121), .A3(KEYINPUT59), .A4(new_n877_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n550_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n878_), .B1(new_n884_), .B2(new_n383_), .ZN(G1340gat));
  INV_X1    g684(.A(KEYINPUT60), .ZN(new_n886_));
  AOI21_X1  g685(.A(G120gat), .B1(new_n677_), .B2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n886_), .B2(G120gat), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n879_), .A2(new_n511_), .A3(new_n877_), .A4(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n619_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n385_), .ZN(G1341gat));
  NAND4_X1  g692(.A1(new_n875_), .A2(new_n381_), .A3(new_n636_), .A4(new_n877_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n679_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n381_), .ZN(G1342gat));
  NAND4_X1  g695(.A1(new_n875_), .A2(new_n379_), .A3(new_n675_), .A4(new_n877_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n710_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n379_), .ZN(G1343gat));
  NOR4_X1   g698(.A1(new_n365_), .A2(new_n449_), .A3(new_n511_), .A4(new_n407_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n879_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n548_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n677_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g705(.A1(new_n901_), .A2(new_n679_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT61), .B(G155gat), .Z(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1346gat));
  OR3_X1    g708(.A1(new_n901_), .A2(G162gat), .A3(new_n667_), .ZN(new_n910_));
  OAI21_X1  g709(.A(G162gat), .B1(new_n901_), .B2(new_n710_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1347gat));
  NOR2_X1   g711(.A1(new_n516_), .A2(new_n448_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n365_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n875_), .A2(new_n548_), .A3(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917_));
  AND3_X1   g716(.A1(new_n916_), .A2(new_n917_), .A3(G169gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n916_), .B2(G169gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n875_), .A2(new_n915_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT22), .B(G169gat), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n548_), .A2(new_n921_), .ZN(new_n922_));
  XOR2_X1   g721(.A(new_n922_), .B(KEYINPUT123), .Z(new_n923_));
  OAI22_X1  g722(.A1(new_n918_), .A2(new_n919_), .B1(new_n920_), .B2(new_n923_), .ZN(G1348gat));
  AND2_X1   g723(.A1(new_n870_), .A2(new_n874_), .ZN(new_n925_));
  OAI21_X1  g724(.A(KEYINPUT124), .B1(new_n925_), .B2(new_n763_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n875_), .A2(new_n927_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n926_), .A2(new_n928_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n914_), .A2(new_n619_), .A3(new_n233_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n875_), .A2(new_n677_), .A3(new_n915_), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n929_), .A2(new_n930_), .B1(new_n233_), .B2(new_n931_), .ZN(G1349gat));
  NOR4_X1   g731(.A1(new_n920_), .A2(new_n302_), .A3(new_n303_), .A4(new_n679_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n926_), .A2(new_n636_), .A3(new_n915_), .A4(new_n928_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n934_), .B2(new_n245_), .ZN(G1350gat));
  OAI21_X1  g734(.A(G190gat), .B1(new_n920_), .B2(new_n710_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n675_), .A2(new_n299_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n920_), .B2(new_n937_), .ZN(G1351gat));
  NAND3_X1  g737(.A1(new_n365_), .A2(new_n513_), .A3(new_n516_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n925_), .A2(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n548_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n677_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  XOR2_X1   g744(.A(new_n945_), .B(KEYINPUT125), .Z(new_n946_));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n948_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n940_), .A2(new_n636_), .A3(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n946_), .A2(new_n947_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(KEYINPUT127), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n950_), .B(new_n952_), .ZN(G1354gat));
  INV_X1    g752(.A(G218gat), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n940_), .A2(new_n954_), .A3(new_n675_), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n925_), .A2(new_n710_), .A3(new_n939_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n956_), .B2(new_n954_), .ZN(G1355gat));
endmodule


