//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G155gat), .B(G162gat), .Z(new_n207_));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT83), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT83), .B1(G141gat), .B2(G148gat), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n209_), .A2(new_n216_), .B1(new_n217_), .B2(new_n207_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT82), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G127gat), .B(G134gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G113gat), .B(G120gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n211_), .B(new_n212_), .C1(new_n225_), .C2(KEYINPUT84), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT84), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(KEYINPUT3), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n225_), .A2(new_n211_), .A3(new_n212_), .A4(KEYINPUT84), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n228_), .B(new_n229_), .C1(new_n217_), .C2(new_n219_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n207_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n221_), .A2(new_n224_), .A3(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n224_), .B(KEYINPUT81), .Z(new_n233_));
  NOR2_X1   g032(.A1(new_n218_), .A2(new_n220_), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n230_), .A2(new_n207_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n232_), .B1(new_n233_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n232_), .B(KEYINPUT4), .C1(new_n233_), .C2(new_n236_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n221_), .A2(new_n231_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n224_), .B(KEYINPUT81), .ZN(new_n242_));
  XOR2_X1   g041(.A(KEYINPUT90), .B(KEYINPUT4), .Z(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n206_), .B(new_n239_), .C1(new_n245_), .C2(new_n238_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n238_), .B1(new_n240_), .B2(new_n244_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n237_), .A2(new_n238_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n205_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G226gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT19), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT23), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT23), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(G183gat), .A3(G190gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(G169gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n262_), .A2(KEYINPUT88), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(KEYINPUT88), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n256_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n254_), .A2(new_n256_), .A3(new_n265_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(G190gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT25), .B(G183gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  OR2_X1    g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(KEYINPUT24), .A3(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n272_), .A2(KEYINPUT24), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n271_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n263_), .A2(new_n264_), .B1(new_n268_), .B2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G211gat), .B(G218gat), .Z(new_n278_));
  INV_X1    g077(.A(KEYINPUT21), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G197gat), .B(G204gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT21), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n278_), .A3(KEYINPUT21), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT20), .B1(new_n277_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n261_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n266_), .A2(new_n267_), .A3(new_n258_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT80), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(new_n290_), .B2(new_n289_), .ZN(new_n292_));
  INV_X1    g091(.A(G190gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT78), .B1(new_n293_), .B2(KEYINPUT26), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n294_), .B(new_n270_), .C1(new_n269_), .C2(KEYINPUT78), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n295_), .A2(new_n257_), .A3(new_n274_), .A4(new_n275_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n296_), .A3(new_n286_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n252_), .B1(new_n287_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n292_), .A2(new_n296_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n284_), .A2(new_n285_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n277_), .A2(new_n286_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT20), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n252_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n302_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G8gat), .B(G36gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G64gat), .B(G92gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT32), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n299_), .A2(new_n306_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT93), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT93), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n299_), .A2(new_n316_), .A3(new_n306_), .A4(new_n313_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n263_), .A2(new_n264_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n276_), .A2(new_n268_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n304_), .B1(new_n321_), .B2(new_n301_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n252_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n297_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n286_), .A2(new_n320_), .A3(new_n262_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT20), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n286_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n252_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(KEYINPUT32), .A3(new_n312_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n250_), .A2(new_n318_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT33), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n249_), .B(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n323_), .B1(new_n322_), .B2(new_n297_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n302_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n311_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n299_), .A2(new_n312_), .A3(new_n306_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n237_), .A2(KEYINPUT91), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n238_), .B1(new_n237_), .B2(KEYINPUT91), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n205_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n240_), .A2(new_n238_), .A3(new_n244_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT92), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n342_), .A2(new_n343_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n341_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n338_), .A2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n331_), .B1(new_n333_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n241_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT29), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n351_), .B1(new_n236_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G22gat), .B(G50gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n350_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT28), .B1(new_n241_), .B2(KEYINPUT29), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n236_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n354_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n349_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G228gat), .A2(G233gat), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n301_), .B(new_n361_), .C1(new_n236_), .C2(new_n352_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(KEYINPUT86), .B(KEYINPUT29), .Z(new_n365_));
  AOI21_X1  g164(.A(new_n286_), .B1(new_n241_), .B2(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n362_), .B(new_n364_), .C1(new_n366_), .C2(new_n361_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n361_), .B1(new_n368_), .B2(new_n301_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n301_), .A2(new_n361_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n241_), .B2(KEYINPUT29), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n363_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n355_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n357_), .A2(new_n358_), .A3(new_n354_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(KEYINPUT85), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n360_), .A2(new_n373_), .A3(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n356_), .A2(new_n359_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n369_), .A2(new_n371_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT87), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n364_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n367_), .A2(KEYINPUT87), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n378_), .A2(new_n381_), .A3(new_n382_), .A4(new_n372_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n377_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n348_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT27), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n336_), .A2(new_n337_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT94), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n337_), .A2(new_n389_), .B1(new_n329_), .B2(new_n311_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n299_), .A2(KEYINPUT94), .A3(new_n312_), .A4(new_n306_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n388_), .B1(new_n392_), .B2(KEYINPUT27), .ZN(new_n393_));
  INV_X1    g192(.A(new_n250_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n384_), .A2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT95), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n250_), .B1(new_n377_), .B2(new_n383_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT95), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n387_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n397_), .B(new_n398_), .C1(new_n388_), .C2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n386_), .A2(new_n396_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G15gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT30), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n300_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(new_n233_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G71gat), .B(G99gat), .ZN(new_n407_));
  INV_X1    g206(.A(G43gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT31), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n406_), .A2(new_n410_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT96), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n393_), .B2(new_n384_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n385_), .B(KEYINPUT96), .C1(new_n388_), .C2(new_n399_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n394_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n401_), .A2(new_n414_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G229gat), .A2(G233gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G43gat), .B(G50gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G29gat), .B(G36gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT70), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n426_), .A2(new_n427_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n425_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n430_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(new_n428_), .A3(new_n424_), .ZN(new_n433_));
  OR2_X1    g232(.A1(G1gat), .A2(G8gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G1gat), .A2(G8gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT74), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT74), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n434_), .A2(new_n438_), .A3(new_n435_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G15gat), .B(G22gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(KEYINPUT14), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n437_), .A2(new_n442_), .A3(new_n441_), .A4(new_n439_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n431_), .A2(new_n433_), .A3(new_n444_), .A4(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n433_), .A2(new_n431_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n423_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n445_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n431_), .A2(new_n433_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT15), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT15), .B1(new_n431_), .B2(new_n433_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n450_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n446_), .A2(new_n422_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n449_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G113gat), .B(G141gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G169gat), .B(G197gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n459_), .B(new_n460_), .Z(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n449_), .B(new_n461_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n421_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G190gat), .B(G218gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G134gat), .B(G162gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT36), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT64), .ZN(new_n473_));
  AND2_X1   g272(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G106gat), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n473_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NOR4_X1   g277(.A1(new_n474_), .A2(new_n475_), .A3(KEYINPUT64), .A4(G106gat), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G99gat), .A2(G106gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT6), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(G99gat), .A3(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(G85gat), .A2(G92gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(G85gat), .A2(G92gat), .ZN(new_n487_));
  OAI22_X1  g286(.A1(new_n486_), .A2(new_n487_), .B1(KEYINPUT9), .B2(G92gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n485_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(KEYINPUT9), .A2(G92gat), .ZN(new_n491_));
  INV_X1    g290(.A(G85gat), .ZN(new_n492_));
  INV_X1    g291(.A(G92gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G85gat), .A2(G92gat), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n491_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT9), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT65), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT65), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT9), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n496_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n490_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n486_), .A2(new_n487_), .ZN(new_n504_));
  INV_X1    g303(.A(G99gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n477_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT66), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n509_), .B1(new_n510_), .B2(new_n506_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n485_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n504_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT8), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n480_), .A2(new_n503_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n509_), .B(KEYINPUT67), .C1(new_n510_), .C2(new_n506_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n485_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n504_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(new_n514_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n515_), .A2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n515_), .A2(new_n522_), .A3(new_n433_), .A4(new_n431_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G232gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT34), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT35), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n525_), .A3(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n528_), .A2(new_n529_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n532_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n524_), .A2(new_n525_), .A3(new_n534_), .A4(new_n530_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n472_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n471_), .A2(KEYINPUT36), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(new_n537_), .A3(new_n535_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n538_), .A2(KEYINPUT73), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(KEYINPUT73), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n536_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(KEYINPUT37), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT37), .ZN(new_n543_));
  AOI211_X1 g342(.A(new_n543_), .B(new_n536_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n546_));
  XOR2_X1   g345(.A(G71gat), .B(G78gat), .Z(new_n547_));
  AND2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n546_), .A2(new_n547_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(new_n450_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G127gat), .B(G155gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G183gat), .B(G211gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n557_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT76), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n557_), .A2(KEYINPUT76), .A3(new_n564_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n562_), .B(KEYINPUT17), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n556_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT77), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n542_), .A2(new_n544_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n505_), .A2(new_n477_), .B1(new_n507_), .B2(KEYINPUT66), .ZN(new_n577_));
  INV_X1    g376(.A(new_n506_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT66), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT7), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n508_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n577_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n520_), .B1(new_n582_), .B2(new_n485_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n496_), .A2(new_n501_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n488_), .A2(new_n489_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n485_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n478_), .A2(new_n479_), .ZN(new_n587_));
  OAI22_X1  g386(.A1(new_n583_), .A2(KEYINPUT8), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n521_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n512_), .B1(new_n511_), .B2(new_n516_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n590_), .B2(new_n518_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n551_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n588_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n553_), .B1(new_n515_), .B2(new_n522_), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT12), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT12), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n588_), .A2(new_n591_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n597_), .B1(new_n598_), .B2(new_n553_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n595_), .A2(new_n596_), .A3(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n592_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n515_), .A2(new_n553_), .A3(new_n522_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n596_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(G120gat), .B(G148gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(G176gat), .B(G204gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT69), .B1(new_n606_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n600_), .A2(new_n605_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT69), .ZN(new_n614_));
  INV_X1    g413(.A(new_n611_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  OAI22_X1  g415(.A1(new_n612_), .A2(new_n616_), .B1(new_n606_), .B2(new_n611_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT13), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n606_), .A2(KEYINPUT69), .A3(new_n611_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n614_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n620_), .A2(new_n621_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(KEYINPUT13), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n619_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n576_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n466_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(G1gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n250_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n421_), .A2(new_n541_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n625_), .A2(new_n465_), .A3(new_n574_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G1gat), .B1(new_n634_), .B2(new_n394_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n629_), .A2(new_n630_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n631_), .A2(new_n635_), .A3(new_n636_), .ZN(G1324gat));
  INV_X1    g436(.A(new_n393_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G8gat), .B1(new_n634_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI211_X1 g440(.A(KEYINPUT39), .B(G8gat), .C1(new_n634_), .C2(new_n638_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n638_), .A2(G8gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n466_), .A2(new_n626_), .A3(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT97), .Z(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n643_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n643_), .B2(new_n646_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1325gat));
  OAI21_X1  g449(.A(G15gat), .B1(new_n634_), .B2(new_n414_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT41), .Z(new_n652_));
  INV_X1    g451(.A(G15gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n627_), .A2(new_n653_), .A3(new_n413_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(G1326gat));
  INV_X1    g454(.A(G22gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n384_), .B(KEYINPUT99), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n627_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n659_));
  INV_X1    g458(.A(new_n634_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n657_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n659_), .B1(new_n661_), .B2(G22gat), .ZN(new_n662_));
  AOI211_X1 g461(.A(KEYINPUT42), .B(new_n656_), .C1(new_n660_), .C2(new_n657_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n658_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT100), .ZN(G1327gat));
  INV_X1    g464(.A(new_n574_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n541_), .ZN(new_n667_));
  NOR4_X1   g466(.A1(new_n623_), .A2(new_n619_), .A3(new_n666_), .A4(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n466_), .A2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G29gat), .B1(new_n669_), .B2(new_n250_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n465_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n624_), .A2(new_n671_), .A3(new_n574_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT101), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n401_), .A2(new_n414_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n418_), .A2(new_n420_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n542_), .A2(new_n544_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n674_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n421_), .A2(KEYINPUT43), .A3(new_n678_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n673_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT44), .B(new_n673_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n250_), .A2(G29gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n670_), .B1(new_n686_), .B2(new_n687_), .ZN(G1328gat));
  NAND3_X1  g487(.A1(new_n684_), .A2(new_n393_), .A3(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G36gat), .ZN(new_n690_));
  NOR2_X1   g489(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n691_));
  XOR2_X1   g490(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n638_), .A2(G36gat), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n677_), .A2(new_n671_), .A3(new_n668_), .A4(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(KEYINPUT103), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(KEYINPUT103), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n695_), .A2(KEYINPUT103), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n695_), .A2(KEYINPUT103), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n692_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n691_), .B1(new_n698_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n690_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n690_), .B2(new_n702_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  NAND4_X1  g505(.A1(new_n684_), .A2(G43gat), .A3(new_n413_), .A4(new_n685_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n669_), .A2(new_n413_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n408_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(G1330gat));
  INV_X1    g511(.A(G50gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n669_), .A2(new_n713_), .A3(new_n657_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n686_), .B2(new_n384_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n684_), .A2(new_n715_), .A3(new_n384_), .A4(new_n685_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G50gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n716_), .B2(new_n718_), .ZN(G1331gat));
  NOR3_X1   g518(.A1(new_n624_), .A2(new_n671_), .A3(new_n574_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n632_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(G57gat), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n394_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT109), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n421_), .A2(new_n671_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n625_), .A2(KEYINPUT107), .A3(new_n575_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n727_), .B1(new_n576_), .B2(new_n624_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n725_), .A2(new_n726_), .A3(new_n728_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n729_), .A2(KEYINPUT108), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(KEYINPUT108), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n250_), .A3(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n724_), .B1(new_n722_), .B2(new_n732_), .ZN(G1332gat));
  OAI21_X1  g532(.A(G64gat), .B1(new_n721_), .B2(new_n638_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT48), .ZN(new_n735_));
  INV_X1    g534(.A(G64gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n729_), .A2(new_n736_), .A3(new_n393_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1333gat));
  INV_X1    g537(.A(G71gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n729_), .A2(new_n739_), .A3(new_n413_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n632_), .A2(new_n413_), .A3(new_n720_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G71gat), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(KEYINPUT49), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(KEYINPUT49), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT110), .Z(G1334gat));
  INV_X1    g545(.A(G78gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n729_), .A2(new_n747_), .A3(new_n657_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n657_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G78gat), .B1(new_n721_), .B2(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(KEYINPUT50), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(KEYINPUT50), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT111), .ZN(G1335gat));
  NOR3_X1   g553(.A1(new_n624_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n725_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G85gat), .B1(new_n756_), .B2(new_n250_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT112), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n680_), .A2(new_n681_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n625_), .A2(new_n465_), .A3(new_n574_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n394_), .A2(new_n492_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(G1336gat));
  NAND3_X1  g562(.A1(new_n756_), .A2(new_n493_), .A3(new_n393_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n759_), .A2(new_n638_), .A3(new_n760_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n493_), .ZN(G1337gat));
  NAND4_X1  g565(.A1(new_n725_), .A2(new_n413_), .A3(new_n476_), .A4(new_n755_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT113), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n761_), .A2(new_n413_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(G99gat), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n756_), .A2(new_n477_), .A3(new_n384_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n760_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n384_), .B(new_n774_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(G106gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n775_), .B2(G106gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n773_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g579(.A1(new_n418_), .A2(new_n413_), .A3(new_n250_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT120), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT12), .B1(new_n523_), .B2(new_n592_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(KEYINPUT12), .B2(new_n603_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n785_), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(new_n596_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n595_), .A2(KEYINPUT55), .A3(new_n599_), .A4(new_n596_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n595_), .A2(new_n599_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n604_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n600_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n786_), .B(new_n789_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n615_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n615_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n795_), .A2(new_n796_), .A3(KEYINPUT117), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n615_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(KEYINPUT117), .A3(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n422_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n462_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n455_), .A2(new_n446_), .A3(new_n423_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n451_), .A2(new_n450_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n423_), .B1(new_n805_), .B2(new_n446_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT115), .B1(new_n806_), .B2(new_n461_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n803_), .A2(new_n804_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n464_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(KEYINPUT116), .A3(new_n464_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n620_), .A2(new_n621_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n800_), .A2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n783_), .B1(new_n797_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n798_), .A2(new_n799_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n615_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n816_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n819_), .A2(KEYINPUT58), .A3(new_n800_), .A4(new_n813_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n815_), .A2(new_n679_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n465_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n811_), .A2(new_n812_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n617_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n824_), .B1(new_n829_), .B2(new_n667_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n824_), .A2(new_n831_), .ZN(new_n832_));
  AOI211_X1 g631(.A(new_n541_), .B(new_n832_), .C1(new_n826_), .C2(new_n828_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n815_), .A2(new_n679_), .A3(new_n820_), .A4(KEYINPUT118), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n823_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n574_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n575_), .A2(new_n624_), .A3(new_n465_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n782_), .B1(new_n837_), .B2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(G113gat), .B1(new_n842_), .B2(new_n671_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n782_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n666_), .B1(new_n834_), .B2(new_n821_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n844_), .B(new_n845_), .C1(new_n846_), .C2(new_n840_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n840_), .B1(new_n836_), .B2(new_n574_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT59), .B1(new_n851_), .B2(new_n782_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(KEYINPUT121), .A3(new_n847_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n671_), .A2(G113gat), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n855_), .B(KEYINPUT122), .Z(new_n856_));
  AOI21_X1  g655(.A(new_n843_), .B1(new_n854_), .B2(new_n856_), .ZN(G1340gat));
  NAND3_X1  g656(.A1(new_n852_), .A2(new_n625_), .A3(new_n847_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT123), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n852_), .A2(new_n860_), .A3(new_n625_), .A4(new_n847_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(G120gat), .A3(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n624_), .A2(KEYINPUT60), .ZN(new_n863_));
  MUX2_X1   g662(.A(new_n863_), .B(KEYINPUT60), .S(G120gat), .Z(new_n864_));
  NAND2_X1  g663(.A1(new_n842_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(G1341gat));
  AOI21_X1  g665(.A(G127gat), .B1(new_n842_), .B2(new_n666_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n666_), .A2(G127gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n854_), .B2(new_n868_), .ZN(G1342gat));
  INV_X1    g668(.A(G134gat), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n678_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n851_), .A2(new_n667_), .A3(new_n782_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(G134gat), .ZN(new_n874_));
  INV_X1    g673(.A(new_n873_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(KEYINPUT124), .A3(new_n870_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n854_), .A2(new_n871_), .B1(new_n874_), .B2(new_n876_), .ZN(G1343gat));
  INV_X1    g676(.A(new_n851_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n413_), .A2(new_n385_), .A3(new_n394_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n638_), .A3(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n465_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(new_n211_), .ZN(G1344gat));
  NOR2_X1   g681(.A1(new_n880_), .A2(new_n624_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n212_), .ZN(G1345gat));
  NOR2_X1   g683(.A1(new_n880_), .A2(new_n574_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT61), .B(G155gat), .Z(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1346gat));
  OAI21_X1  g686(.A(G162gat), .B1(new_n880_), .B2(new_n678_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n667_), .A2(G162gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n880_), .B2(new_n889_), .ZN(G1347gat));
  OR2_X1    g689(.A1(new_n846_), .A2(new_n840_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n638_), .A2(new_n419_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n657_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n891_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT22), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n897_), .A3(new_n671_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n898_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n895_), .A2(new_n465_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n897_), .ZN(new_n902_));
  INV_X1    g701(.A(G169gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n901_), .B2(new_n900_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n899_), .B1(new_n902_), .B2(new_n904_), .ZN(G1348gat));
  AOI21_X1  g704(.A(G176gat), .B1(new_n896_), .B2(new_n625_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n851_), .A2(new_n384_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n625_), .A2(G176gat), .A3(new_n892_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n906_), .B1(new_n907_), .B2(new_n909_), .ZN(G1349gat));
  NOR2_X1   g709(.A1(new_n574_), .A2(new_n270_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n896_), .A2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n893_), .A2(new_n574_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n907_), .A2(new_n913_), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n912_), .B(KEYINPUT125), .C1(new_n914_), .C2(G183gat), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n895_), .A2(new_n270_), .A3(new_n574_), .ZN(new_n917_));
  AOI21_X1  g716(.A(G183gat), .B1(new_n907_), .B2(new_n913_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n916_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n915_), .A2(new_n919_), .ZN(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n895_), .B2(new_n678_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n541_), .A2(new_n269_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n895_), .B2(new_n922_), .ZN(G1351gat));
  NOR4_X1   g722(.A1(new_n851_), .A2(new_n413_), .A3(new_n638_), .A4(new_n395_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n671_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n625_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g727(.A(new_n574_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n924_), .A2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  XOR2_X1   g730(.A(new_n931_), .B(KEYINPUT126), .Z(new_n932_));
  XNOR2_X1  g731(.A(new_n930_), .B(new_n932_), .ZN(G1354gat));
  NAND2_X1  g732(.A1(new_n924_), .A2(new_n541_), .ZN(new_n934_));
  XOR2_X1   g733(.A(KEYINPUT127), .B(G218gat), .Z(new_n935_));
  NOR2_X1   g734(.A1(new_n678_), .A2(new_n935_), .ZN(new_n936_));
  AOI22_X1  g735(.A1(new_n934_), .A2(new_n935_), .B1(new_n924_), .B2(new_n936_), .ZN(G1355gat));
endmodule


