//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_;
  INV_X1    g000(.A(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT26), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT26), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(G183gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT25), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT25), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G183gat), .ZN(new_n209_));
  AND4_X1   g008(.A1(new_n203_), .A2(new_n205_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT78), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT24), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(new_n210_), .A2(new_n216_), .A3(new_n221_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n214_), .A2(KEYINPUT24), .A3(new_n215_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT79), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT79), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G169gat), .A3(G176gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT80), .B1(new_n223_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n214_), .A2(KEYINPUT24), .A3(new_n215_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT80), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n231_), .A2(new_n228_), .A3(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n222_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n206_), .A2(new_n202_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n219_), .A2(new_n220_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT82), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT81), .B(G176gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT22), .B(G169gat), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n228_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(new_n237_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n234_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G71gat), .B(G99gat), .ZN(new_n245_));
  INV_X1    g044(.A(G43gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n244_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G127gat), .B(G134gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G113gat), .B(G120gat), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n249_), .A2(new_n250_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n248_), .B(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G227gat), .A2(G233gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n255_), .B(G15gat), .Z(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT30), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT31), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n254_), .A2(new_n259_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G141gat), .B(G148gat), .Z(new_n264_));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT1), .ZN(new_n266_));
  INV_X1    g065(.A(G155gat), .ZN(new_n267_));
  INV_X1    g066(.A(G162gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n265_), .A2(KEYINPUT1), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n264_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G141gat), .A2(G148gat), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT2), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT3), .ZN(new_n276_));
  INV_X1    g075(.A(G141gat), .ZN(new_n277_));
  INV_X1    g076(.A(G148gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n281_));
  AND4_X1   g080(.A1(new_n275_), .A2(new_n279_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT83), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT83), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n269_), .A2(new_n286_), .A3(new_n265_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n272_), .B1(new_n282_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT29), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G197gat), .B(G204gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT21), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G197gat), .A2(G204gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(KEYINPUT21), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G218gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G211gat), .ZN(new_n298_));
  INV_X1    g097(.A(G211gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G218gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT85), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n298_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n301_), .B1(new_n298_), .B2(new_n300_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n293_), .B(new_n296_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n296_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n298_), .A2(new_n300_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT85), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n298_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n304_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n290_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G228gat), .ZN(new_n312_));
  INV_X1    g111(.A(G233gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n290_), .B(new_n310_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G78gat), .B(G106gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n318_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n315_), .A2(new_n316_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT84), .ZN(new_n323_));
  OR3_X1    g122(.A1(new_n289_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT28), .B1(new_n289_), .B2(KEYINPUT29), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G22gat), .B(G50gat), .Z(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n328_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n329_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n331_), .B1(new_n332_), .B2(new_n326_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n322_), .A2(new_n330_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n319_), .A2(KEYINPUT86), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT87), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n321_), .A2(new_n336_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n315_), .A2(KEYINPUT87), .A3(new_n316_), .A4(new_n320_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT86), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n317_), .A2(new_n339_), .A3(new_n318_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n335_), .A2(new_n337_), .A3(new_n338_), .A4(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n333_), .A2(new_n330_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n334_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G1gat), .B(G29gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G57gat), .B(G85gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n289_), .A2(KEYINPUT94), .A3(new_n253_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n279_), .A2(new_n275_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n353_), .B(new_n272_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(KEYINPUT4), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT4), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n289_), .A2(KEYINPUT94), .A3(new_n253_), .A4(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n350_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n289_), .A2(new_n253_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n354_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n360_), .A2(new_n350_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n349_), .B1(new_n358_), .B2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(KEYINPUT33), .B1(new_n362_), .B2(KEYINPUT96), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT96), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n364_), .B(new_n349_), .C1(new_n358_), .C2(new_n361_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n363_), .A2(KEYINPUT97), .A3(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(KEYINPUT33), .B(new_n349_), .C1(new_n358_), .C2(new_n361_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n355_), .A2(new_n350_), .A3(new_n357_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n349_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n368_), .B(new_n369_), .C1(new_n350_), .C2(new_n360_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT89), .ZN(new_n373_));
  XOR2_X1   g172(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n304_), .A2(new_n309_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n207_), .A2(new_n209_), .A3(KEYINPUT90), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT90), .B1(new_n207_), .B2(new_n209_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n203_), .A2(new_n205_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n214_), .A2(new_n215_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT91), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n224_), .A2(new_n383_), .A3(KEYINPUT24), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n224_), .B2(KEYINPUT24), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n382_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT92), .B1(new_n381_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n379_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n380_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n207_), .A2(new_n209_), .A3(KEYINPUT90), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT92), .ZN(new_n393_));
  INV_X1    g192(.A(new_n386_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n394_), .A2(new_n384_), .A3(new_n215_), .A4(new_n214_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n392_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n217_), .B(new_n218_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n388_), .A2(new_n396_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n241_), .A2(new_n236_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n377_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n234_), .A2(new_n377_), .A3(new_n243_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT20), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n376_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n406_), .B1(new_n244_), .B2(new_n310_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n400_), .A2(new_n377_), .A3(new_n401_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n375_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G8gat), .B(G36gat), .Z(new_n411_));
  XNOR2_X1  g210(.A(G64gat), .B(G92gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n410_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n415_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n405_), .A2(new_n417_), .A3(new_n409_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n371_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT97), .B1(new_n363_), .B2(new_n365_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n366_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n402_), .A2(new_n404_), .A3(new_n376_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n375_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT32), .B(new_n417_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n424_));
  OR3_X1    g223(.A1(new_n358_), .A2(new_n361_), .A3(new_n349_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n362_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n417_), .A2(KEYINPUT32), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n405_), .A2(new_n427_), .A3(new_n409_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n344_), .B1(new_n421_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n426_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433_));
  INV_X1    g232(.A(new_n418_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n417_), .B1(new_n405_), .B2(new_n409_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n415_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(KEYINPUT27), .A3(new_n418_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n343_), .A2(new_n432_), .A3(new_n436_), .A4(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n263_), .B1(new_n431_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n260_), .A2(new_n432_), .A3(new_n261_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(new_n438_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT98), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT98), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n436_), .A2(new_n444_), .A3(new_n438_), .ZN(new_n445_));
  AOI211_X1 g244(.A(new_n343_), .B(new_n441_), .C1(new_n443_), .C2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n440_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT14), .ZN(new_n448_));
  XOR2_X1   g247(.A(KEYINPUT72), .B(G1gat), .Z(new_n449_));
  XOR2_X1   g248(.A(KEYINPUT73), .B(G8gat), .Z(new_n450_));
  AOI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G15gat), .B(G22gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(G1gat), .B(G8gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OR3_X1    g253(.A1(new_n451_), .A2(new_n452_), .A3(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n454_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G29gat), .B(G36gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G43gat), .B(G50gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT77), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(G229gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n457_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n460_), .B(KEYINPUT15), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n462_), .B1(new_n465_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n468_), .B1(new_n470_), .B2(new_n464_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G113gat), .B(G141gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G169gat), .B(G197gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n472_), .B(new_n473_), .Z(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n474_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n468_), .B(new_n476_), .C1(new_n470_), .C2(new_n464_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n447_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G85gat), .B(G92gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT9), .ZN(new_n483_));
  INV_X1    g282(.A(G85gat), .ZN(new_n484_));
  INV_X1    g283(.A(G92gat), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n484_), .A2(new_n485_), .A3(KEYINPUT9), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT6), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(G99gat), .A3(G106gat), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n486_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G106gat), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT65), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT65), .ZN(new_n497_));
  NOR4_X1   g296(.A1(new_n492_), .A2(new_n493_), .A3(new_n497_), .A4(G106gat), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n483_), .B(new_n491_), .C1(new_n496_), .C2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n488_), .A2(new_n490_), .ZN(new_n504_));
  AOI211_X1 g303(.A(KEYINPUT8), .B(new_n481_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT8), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n507_));
  INV_X1    g306(.A(G99gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n508_), .A3(new_n495_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n504_), .A2(new_n500_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n506_), .B1(new_n510_), .B2(new_n482_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n499_), .B1(new_n505_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT66), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n499_), .B(KEYINPUT66), .C1(new_n505_), .C2(new_n511_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G57gat), .B(G64gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT11), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G71gat), .B(G78gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n517_), .A2(KEYINPUT11), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(new_n519_), .A3(KEYINPUT11), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n516_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n525_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n514_), .A2(new_n527_), .A3(new_n515_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(KEYINPUT67), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G230gat), .A2(G233gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT64), .Z(new_n531_));
  OAI211_X1 g330(.A(new_n529_), .B(new_n531_), .C1(KEYINPUT67), .C2(new_n526_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n531_), .B1(new_n516_), .B2(new_n525_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT12), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n528_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT69), .ZN(new_n536_));
  INV_X1    g335(.A(new_n499_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT68), .B1(new_n505_), .B2(new_n511_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n488_), .A2(new_n490_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n509_), .A2(new_n500_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n482_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT8), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT68), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n510_), .A2(new_n506_), .A3(new_n482_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n537_), .B1(new_n538_), .B2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n523_), .A2(KEYINPUT12), .A3(new_n524_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n536_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n505_), .A2(new_n511_), .A3(KEYINPUT68), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n543_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n499_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n547_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(KEYINPUT69), .A3(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n533_), .A2(new_n535_), .A3(new_n548_), .A4(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n532_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G120gat), .B(G148gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT5), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G176gat), .B(G204gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n532_), .A2(new_n554_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n560_), .A2(KEYINPUT13), .A3(new_n562_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n516_), .A2(new_n460_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT70), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT34), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT35), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n551_), .A2(new_n469_), .B1(new_n574_), .B2(new_n573_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n570_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n569_), .A2(KEYINPUT70), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT70), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n580_), .B1(new_n516_), .B2(new_n460_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n577_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n575_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G190gat), .B(G218gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT71), .ZN(new_n585_));
  XOR2_X1   g384(.A(G134gat), .B(G162gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n578_), .A2(new_n583_), .A3(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n587_), .B(new_n588_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT37), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n578_), .A2(new_n583_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n578_), .A2(new_n583_), .A3(new_n590_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n594_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G127gat), .B(G155gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G183gat), .B(G211gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n457_), .B(new_n525_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT74), .Z(new_n610_));
  XNOR2_X1  g409(.A(new_n608_), .B(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n607_), .B1(new_n611_), .B2(KEYINPUT76), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT17), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT17), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n611_), .B2(new_n607_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n613_), .B1(new_n612_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n601_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n568_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n432_), .A2(new_n449_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n480_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n620_), .A2(KEYINPUT99), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(KEYINPUT99), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(KEYINPUT38), .A3(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n567_), .A2(new_n478_), .A3(new_n616_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n597_), .A2(new_n599_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n447_), .A2(new_n628_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n626_), .A2(KEYINPUT101), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT101), .B1(new_n626_), .B2(new_n629_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n426_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(G1gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT38), .B1(new_n621_), .B2(new_n622_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n634_), .A2(KEYINPUT102), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(KEYINPUT102), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n623_), .B(new_n633_), .C1(new_n635_), .C2(new_n636_), .ZN(G1324gat));
  NAND2_X1  g436(.A1(new_n480_), .A2(new_n618_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n443_), .A2(new_n445_), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n638_), .A2(new_n450_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n639_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n626_), .A2(new_n641_), .A3(new_n629_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n642_), .A2(new_n643_), .A3(G8gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n642_), .B2(G8gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n640_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n263_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(G15gat), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n638_), .A2(G15gat), .A3(new_n262_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT103), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n650_), .B1(new_n649_), .B2(G15gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n648_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n655_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n657_), .A2(KEYINPUT104), .A3(new_n651_), .A4(new_n653_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(G1326gat));
  OR3_X1    g458(.A1(new_n638_), .A2(G22gat), .A3(new_n344_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n343_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n661_), .A2(new_n662_), .A3(G22gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n661_), .B2(G22gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n660_), .B1(new_n663_), .B2(new_n664_), .ZN(G1327gat));
  INV_X1    g464(.A(new_n616_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n628_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n568_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n480_), .A2(new_n668_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n669_), .A2(G29gat), .A3(new_n432_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n568_), .A2(new_n479_), .A3(new_n616_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n601_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n672_), .B1(new_n440_), .B2(new_n446_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT43), .B1(new_n673_), .B2(KEYINPUT105), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n362_), .A2(KEYINPUT96), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT33), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(new_n676_), .A3(new_n365_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT97), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n363_), .A2(KEYINPUT97), .A3(new_n365_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n434_), .A2(new_n435_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .A4(new_n371_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n343_), .B1(new_n682_), .B2(new_n429_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n439_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n262_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n441_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n639_), .A2(new_n344_), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n601_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n671_), .B1(new_n674_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n673_), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n690_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT44), .B1(new_n697_), .B2(new_n671_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n694_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n426_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n670_), .B1(new_n700_), .B2(G29gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT106), .ZN(G1328gat));
  OR2_X1    g501(.A1(new_n641_), .A2(KEYINPUT108), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n641_), .A2(KEYINPUT108), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n669_), .A2(G36gat), .A3(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT45), .Z(new_n708_));
  NAND2_X1  g507(.A1(new_n692_), .A2(new_n693_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n697_), .A2(KEYINPUT44), .A3(new_n671_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n641_), .A3(new_n710_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n711_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT107), .B1(new_n711_), .B2(G36gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n708_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT46), .B(new_n708_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1329gat));
  NOR4_X1   g517(.A1(new_n694_), .A2(new_n698_), .A3(new_n246_), .A4(new_n262_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT109), .B(G43gat), .ZN(new_n720_));
  INV_X1    g519(.A(new_n669_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(new_n263_), .ZN(new_n722_));
  OR3_X1    g521(.A1(new_n719_), .A2(KEYINPUT47), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT47), .B1(new_n719_), .B2(new_n722_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1330gat));
  NAND3_X1  g524(.A1(new_n699_), .A2(KEYINPUT110), .A3(new_n343_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G50gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT110), .B1(new_n699_), .B2(new_n343_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n344_), .A2(G50gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT111), .ZN(new_n730_));
  OAI22_X1  g529(.A1(new_n727_), .A2(new_n728_), .B1(new_n669_), .B2(new_n730_), .ZN(G1331gat));
  NOR2_X1   g530(.A1(new_n447_), .A2(new_n478_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n617_), .A2(new_n567_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G57gat), .B1(new_n735_), .B2(new_n426_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n666_), .A2(new_n478_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n629_), .A2(new_n568_), .A3(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(G57gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n426_), .B2(KEYINPUT112), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(KEYINPUT112), .B2(new_n739_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n736_), .B1(new_n738_), .B2(new_n741_), .ZN(G1332gat));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n735_), .A2(new_n743_), .A3(new_n705_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n738_), .B2(new_n705_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n746_), .ZN(new_n748_));
  XOR2_X1   g547(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n749_));
  AND3_X1   g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n744_), .B1(new_n750_), .B2(new_n751_), .ZN(G1333gat));
  INV_X1    g551(.A(G71gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n738_), .B2(new_n263_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT49), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n735_), .A2(new_n753_), .A3(new_n263_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1334gat));
  NAND2_X1  g556(.A1(new_n738_), .A2(new_n343_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G78gat), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT50), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n344_), .A2(G78gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n734_), .B2(new_n761_), .ZN(G1335gat));
  NOR3_X1   g561(.A1(new_n567_), .A2(new_n478_), .A3(new_n616_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n697_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n432_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n667_), .A2(new_n567_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n732_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n732_), .B2(new_n768_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n484_), .A3(new_n426_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n766_), .A2(new_n773_), .ZN(G1336gat));
  OAI21_X1  g573(.A(G92gat), .B1(new_n765_), .B2(new_n706_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(new_n485_), .A3(new_n641_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1337gat));
  NOR4_X1   g576(.A1(new_n771_), .A2(new_n262_), .A3(new_n493_), .A4(new_n492_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n508_), .B1(new_n764_), .B2(new_n263_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g580(.A1(new_n772_), .A2(new_n495_), .A3(new_n343_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n763_), .B(new_n343_), .C1(new_n674_), .C2(new_n691_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n697_), .A2(KEYINPUT116), .A3(new_n343_), .A4(new_n763_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n495_), .B1(KEYINPUT117), .B2(KEYINPUT52), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n787_), .A2(new_n788_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n790_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n788_), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n792_), .B(new_n793_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n782_), .B1(new_n791_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT53), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n782_), .B(new_n797_), .C1(new_n791_), .C2(new_n794_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1339gat));
  NAND2_X1  g598(.A1(new_n478_), .A2(new_n562_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n554_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n554_), .A2(KEYINPUT119), .A3(new_n801_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n535_), .A2(new_n553_), .A3(new_n526_), .A4(new_n548_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n531_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(new_n805_), .A3(new_n807_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n535_), .A2(new_n548_), .A3(new_n553_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n809_), .A2(KEYINPUT120), .A3(KEYINPUT55), .A4(new_n533_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT120), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n554_), .B2(new_n801_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n559_), .B1(new_n808_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n802_), .A2(new_n803_), .B1(new_n531_), .B2(new_n806_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n810_), .A2(new_n812_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n805_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(KEYINPUT56), .A3(new_n559_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n800_), .B1(new_n816_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n470_), .A2(new_n464_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n462_), .B1(new_n466_), .B2(new_n465_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n822_), .B(new_n476_), .C1(new_n464_), .C2(new_n823_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n563_), .A2(new_n475_), .A3(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n627_), .B1(new_n821_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT57), .B(new_n627_), .C1(new_n821_), .C2(new_n825_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n824_), .A2(new_n475_), .A3(new_n562_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n819_), .A2(KEYINPUT56), .A3(new_n559_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT56), .B1(new_n819_), .B2(new_n559_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n830_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n830_), .B(KEYINPUT58), .C1(new_n831_), .C2(new_n832_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n672_), .A3(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n828_), .A2(new_n829_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n666_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n737_), .A2(new_n567_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT118), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n737_), .A2(new_n567_), .A3(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n841_), .A2(new_n601_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT54), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n841_), .A2(new_n846_), .A3(new_n601_), .A4(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n839_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NOR4_X1   g649(.A1(new_n641_), .A2(new_n432_), .A3(new_n343_), .A4(new_n262_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(G113gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n478_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n849_), .A2(KEYINPUT59), .A3(new_n851_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n479_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n855_), .B1(new_n859_), .B2(new_n854_), .ZN(G1340gat));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n861_));
  AOI21_X1  g660(.A(G120gat), .B1(new_n568_), .B2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(new_n861_), .B2(G120gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT121), .B1(new_n853_), .B2(new_n863_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n853_), .A2(KEYINPUT121), .A3(new_n863_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n567_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n866_));
  INV_X1    g665(.A(G120gat), .ZN(new_n867_));
  OAI22_X1  g666(.A1(new_n864_), .A2(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(G1341gat));
  INV_X1    g667(.A(G127gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n853_), .A2(new_n869_), .A3(new_n616_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n666_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n869_), .ZN(G1342gat));
  INV_X1    g671(.A(G134gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n853_), .A2(new_n873_), .A3(new_n628_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n601_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n873_), .ZN(G1343gat));
  NAND4_X1  g675(.A1(new_n706_), .A2(new_n426_), .A3(new_n343_), .A4(new_n262_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT122), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n850_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n478_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n568_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n616_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT61), .B(G155gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1346gat));
  NAND3_X1  g685(.A1(new_n879_), .A2(new_n268_), .A3(new_n628_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n850_), .A2(new_n878_), .A3(new_n601_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n268_), .ZN(G1347gat));
  NAND3_X1  g688(.A1(new_n705_), .A2(new_n344_), .A3(new_n686_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n850_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  OAI211_X1 g691(.A(KEYINPUT62), .B(G169gat), .C1(new_n892_), .C2(new_n479_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n850_), .A2(new_n479_), .A3(new_n890_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n212_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n240_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n893_), .A2(new_n896_), .A3(new_n897_), .ZN(G1348gat));
  NAND4_X1  g697(.A1(new_n891_), .A2(KEYINPUT123), .A3(G176gat), .A4(new_n568_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n891_), .A2(G176gat), .A3(new_n568_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n239_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n891_), .B2(new_n568_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n899_), .B1(new_n902_), .B2(new_n904_), .ZN(G1349gat));
  AOI21_X1  g704(.A(G183gat), .B1(new_n891_), .B2(new_n616_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n892_), .A2(new_n666_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n389_), .A2(new_n391_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n892_), .B2(new_n601_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n628_), .A2(new_n390_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT124), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n892_), .B2(new_n912_), .ZN(G1351gat));
  NOR2_X1   g712(.A1(new_n344_), .A2(new_n426_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n705_), .A2(new_n914_), .A3(new_n262_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n915_), .B1(new_n839_), .B2(new_n848_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n478_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n568_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g719(.A(new_n666_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n916_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(KEYINPUT125), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n922_), .A2(KEYINPUT125), .ZN(new_n925_));
  OAI22_X1  g724(.A1(new_n924_), .A2(new_n925_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n926_));
  INV_X1    g725(.A(new_n925_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n927_), .A2(new_n928_), .A3(new_n923_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n926_), .A2(new_n929_), .ZN(G1354gat));
  NAND3_X1  g729(.A1(new_n916_), .A2(G218gat), .A3(new_n672_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932_));
  INV_X1    g731(.A(new_n915_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n849_), .A2(new_n932_), .A3(new_n628_), .A4(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n297_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n932_), .B1(new_n916_), .B2(new_n628_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n931_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(KEYINPUT127), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n939_), .B(new_n931_), .C1(new_n935_), .C2(new_n936_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1355gat));
endmodule


