//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G43gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT84), .B(G176gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G169gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT85), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(KEYINPUT85), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT23), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n210_), .B(new_n211_), .C1(new_n212_), .C2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT25), .B(G183gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(KEYINPUT82), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n214_), .A2(KEYINPUT26), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n214_), .A2(KEYINPUT26), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT82), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n225_), .B1(KEYINPUT25), .B2(new_n213_), .ZN(new_n226_));
  NOR3_X1   g025(.A1(new_n221_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G169gat), .ZN(new_n228_));
  INV_X1    g027(.A(G176gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(KEYINPUT24), .A3(new_n208_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n231_), .B1(KEYINPUT24), .B2(new_n230_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n227_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT83), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n217_), .B(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n215_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n219_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G227gat), .A2(G233gat), .ZN(new_n239_));
  INV_X1    g038(.A(G15gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT30), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G113gat), .B(G120gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n246_), .A2(KEYINPUT31), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(KEYINPUT31), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(KEYINPUT86), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n219_), .A2(new_n237_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n242_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n243_), .A2(new_n249_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n249_), .B1(new_n243_), .B2(new_n252_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n204_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n255_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(new_n203_), .A3(new_n253_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT88), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266_));
  INV_X1    g065(.A(G141gat), .ZN(new_n267_));
  INV_X1    g066(.A(G148gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT2), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n269_), .B(new_n270_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n262_), .B1(new_n265_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT89), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  OAI211_X1 g075(.A(KEYINPUT89), .B(new_n262_), .C1(new_n265_), .C2(new_n273_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OR3_X1    g077(.A1(new_n261_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT87), .B1(new_n261_), .B2(KEYINPUT1), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n261_), .A2(KEYINPUT1), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n279_), .A2(new_n260_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n267_), .A2(new_n268_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n272_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n278_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n246_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n284_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n246_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(KEYINPUT4), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G225gat), .A2(G233gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OR3_X1    g092(.A1(new_n288_), .A2(KEYINPUT4), .A3(new_n289_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n291_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n286_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G1gat), .B(G29gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(G85gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT0), .B(G57gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n295_), .A2(new_n296_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n301_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT104), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n304_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT104), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(new_n302_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n259_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G8gat), .B(G36gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT18), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G64gat), .B(G92gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n312_), .B(new_n313_), .Z(new_n314_));
  INV_X1    g113(.A(G204gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G197gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT91), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT21), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G197gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(G204gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n319_), .B(KEYINPUT92), .C1(KEYINPUT91), .C2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT92), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n322_), .A2(KEYINPUT91), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n324_), .B1(new_n325_), .B2(new_n318_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G211gat), .B(G218gat), .Z(new_n328_));
  OR3_X1    g127(.A1(new_n322_), .A2(KEYINPUT93), .A3(KEYINPUT21), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT93), .B1(new_n322_), .B2(KEYINPUT21), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n322_), .A2(KEYINPUT21), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n328_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT94), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n327_), .A2(new_n331_), .B1(new_n328_), .B2(new_n333_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT94), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n250_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT20), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G226gat), .A2(G233gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n220_), .A2(new_n223_), .A3(new_n222_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n345_), .A2(new_n232_), .A3(new_n218_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n236_), .B1(G183gat), .B2(G190gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n208_), .B(KEYINPUT98), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n207_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n346_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  AOI211_X1 g149(.A(new_n341_), .B(new_n344_), .C1(new_n350_), .C2(new_n337_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n340_), .A2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT20), .B1(new_n350_), .B2(new_n337_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n336_), .A2(new_n339_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n354_), .B2(new_n238_), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n344_), .B(KEYINPUT97), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n314_), .B(new_n352_), .C1(new_n355_), .C2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT99), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n250_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n356_), .B1(new_n361_), .B2(new_n353_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n362_), .A2(KEYINPUT99), .A3(new_n314_), .A4(new_n352_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n352_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n314_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n360_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT27), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n350_), .A2(new_n337_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT20), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT103), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT103), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n373_), .A3(KEYINPUT20), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n340_), .A3(new_n374_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n375_), .A2(new_n344_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n376_));
  OAI211_X1 g175(.A(KEYINPUT27), .B(new_n358_), .C1(new_n376_), .C2(new_n314_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n369_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n285_), .A2(KEYINPUT29), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G228gat), .A2(G233gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT90), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n379_), .A2(new_n336_), .A3(new_n339_), .A4(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n335_), .B1(new_n288_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(G228gat), .A3(G233gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G78gat), .B(G106gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n382_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT95), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n288_), .A2(new_n383_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G22gat), .B(G50gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT28), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n390_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n382_), .A2(new_n385_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n386_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n388_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n394_), .B(new_n397_), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n310_), .A2(new_n378_), .A3(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n305_), .A2(new_n308_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n400_), .A2(new_n398_), .A3(new_n369_), .A4(new_n377_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n314_), .A2(KEYINPUT32), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  OAI22_X1  g202(.A1(new_n303_), .A2(new_n304_), .B1(new_n364_), .B2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n376_), .A2(new_n402_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n286_), .A2(new_n290_), .A3(new_n293_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n300_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n291_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT102), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n291_), .A2(KEYINPUT102), .A3(new_n294_), .A4(new_n292_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n295_), .A2(KEYINPUT33), .A3(new_n296_), .A4(new_n301_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n367_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n302_), .A2(KEYINPUT100), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT100), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n295_), .A2(new_n418_), .A3(new_n296_), .A4(new_n301_), .ZN(new_n419_));
  XOR2_X1   g218(.A(KEYINPUT101), .B(KEYINPUT33), .Z(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n406_), .B1(new_n416_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n401_), .B1(new_n422_), .B2(new_n398_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n259_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n399_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G29gat), .B(G36gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G43gat), .B(G50gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G15gat), .B(G22gat), .ZN(new_n429_));
  INV_X1    g228(.A(G1gat), .ZN(new_n430_));
  INV_X1    g229(.A(G8gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT14), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G8gat), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n434_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n428_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT78), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n428_), .B1(new_n436_), .B2(new_n435_), .ZN(new_n439_));
  OR2_X1    g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(G229gat), .A3(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n438_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n428_), .B(KEYINPUT15), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n435_), .A2(new_n436_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G229gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT79), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n442_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n441_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT80), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G113gat), .B(G141gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G169gat), .B(G197gat), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n451_), .B(new_n452_), .Z(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OR3_X1    g253(.A1(new_n449_), .A2(new_n450_), .A3(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n454_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT81), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n425_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G57gat), .B(G64gat), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n460_), .A2(KEYINPUT11), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(KEYINPUT11), .ZN(new_n462_));
  XOR2_X1   g261(.A(G71gat), .B(G78gat), .Z(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n462_), .A2(new_n463_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G99gat), .A2(G106gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G106gat), .ZN(new_n470_));
  XOR2_X1   g269(.A(KEYINPUT10), .B(G99gat), .Z(new_n471_));
  AOI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT9), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT65), .B(G92gat), .ZN(new_n474_));
  INV_X1    g273(.A(G85gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(G85gat), .A2(G92gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G85gat), .A2(G92gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n479_), .B1(new_n481_), .B2(KEYINPUT9), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n482_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n472_), .B1(new_n478_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT8), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT67), .B1(G99gat), .B2(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT7), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NOR3_X1   g287(.A1(KEYINPUT67), .A2(G99gat), .A3(G106gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT68), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  OR3_X1    g289(.A1(KEYINPUT67), .A2(G99gat), .A3(G106gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT68), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n487_), .A4(new_n486_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT70), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n468_), .A2(KEYINPUT69), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT69), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT6), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n496_), .A2(new_n498_), .A3(new_n467_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n467_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n495_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n467_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n497_), .A2(KEYINPUT6), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n468_), .A2(KEYINPUT69), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n496_), .A2(new_n498_), .A3(new_n467_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(KEYINPUT70), .A3(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n494_), .A2(new_n501_), .A3(new_n507_), .A4(new_n508_), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n481_), .A2(new_n479_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n485_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n508_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n469_), .A2(new_n513_), .ZN(new_n514_));
  AOI211_X1 g313(.A(KEYINPUT8), .B(new_n510_), .C1(new_n494_), .C2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n466_), .B(new_n484_), .C1(new_n512_), .C2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G230gat), .A2(G233gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n517_), .B(KEYINPUT64), .Z(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n484_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT12), .ZN(new_n522_));
  INV_X1    g321(.A(new_n466_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n522_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n520_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n521_), .A2(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n516_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n518_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G120gat), .B(G148gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n530_), .A2(new_n536_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(KEYINPUT13), .A3(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n521_), .A2(new_n443_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT73), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n428_), .B(new_n484_), .C1(new_n512_), .C2(new_n515_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G232gat), .A2(G233gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT34), .Z(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .A4(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n549_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n544_), .A2(new_n546_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n550_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n546_), .B2(KEYINPUT73), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n551_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT75), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n560_), .B(KEYINPUT36), .Z(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT74), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT75), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n564_), .B(new_n551_), .C1(new_n553_), .C2(new_n555_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n557_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n560_), .A2(KEYINPUT36), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n556_), .A2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT76), .B(KEYINPUT37), .Z(new_n569_));
  NAND3_X1  g368(.A1(new_n566_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n568_), .B1(new_n556_), .B2(new_n562_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT37), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n444_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(new_n523_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G127gat), .B(G155gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT16), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT17), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n576_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT77), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n580_), .A2(new_n581_), .ZN(new_n585_));
  OR3_X1    g384(.A1(new_n576_), .A2(new_n582_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n543_), .A2(new_n573_), .A3(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n459_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n400_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n430_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n566_), .A2(new_n568_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n425_), .A2(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n543_), .A2(new_n457_), .A3(new_n587_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G1gat), .B1(new_n598_), .B2(new_n400_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n591_), .A2(new_n592_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n593_), .A2(new_n599_), .A3(new_n600_), .ZN(G1324gat));
  NAND3_X1  g400(.A1(new_n589_), .A2(new_n431_), .A3(new_n378_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n603_));
  INV_X1    g402(.A(new_n598_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n378_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n603_), .B1(new_n605_), .B2(G8gat), .ZN(new_n606_));
  AOI211_X1 g405(.A(KEYINPUT39), .B(new_n431_), .C1(new_n604_), .C2(new_n378_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n602_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT40), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  OAI211_X1 g409(.A(KEYINPUT40), .B(new_n602_), .C1(new_n606_), .C2(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(G1325gat));
  NAND2_X1  g411(.A1(new_n604_), .A2(new_n259_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(G15gat), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT105), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT105), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n616_), .A3(G15gat), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT41), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n615_), .A2(KEYINPUT41), .A3(new_n617_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n589_), .A2(new_n240_), .A3(new_n259_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(G1326gat));
  INV_X1    g422(.A(new_n398_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G22gat), .B1(new_n598_), .B2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT42), .ZN(new_n626_));
  INV_X1    g425(.A(G22gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n589_), .A2(new_n627_), .A3(new_n398_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1327gat));
  NAND2_X1  g428(.A1(new_n570_), .A2(new_n572_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT43), .B1(new_n425_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n360_), .A2(new_n366_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n413_), .A2(new_n414_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n633_), .A2(new_n634_), .A3(new_n421_), .A4(new_n363_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n406_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n624_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n259_), .B1(new_n638_), .B2(new_n401_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n632_), .B(new_n573_), .C1(new_n639_), .C2(new_n399_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n631_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n457_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n541_), .A2(new_n642_), .A3(new_n542_), .A4(new_n587_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT106), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT44), .B1(new_n641_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n647_), .B(new_n644_), .C1(new_n631_), .C2(new_n640_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(new_n590_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G29gat), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n595_), .A2(new_n587_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n543_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n459_), .A2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n400_), .A2(G29gat), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT107), .Z(new_n656_));
  OAI21_X1  g455(.A(new_n651_), .B1(new_n654_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(KEYINPUT46), .ZN(new_n658_));
  INV_X1    g457(.A(G36gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n649_), .B2(new_n378_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n459_), .A2(new_n659_), .A3(new_n378_), .A4(new_n653_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n658_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n641_), .A2(new_n645_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n647_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n641_), .A2(KEYINPUT44), .A3(new_n645_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n378_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G36gat), .ZN(new_n669_));
  INV_X1    g468(.A(new_n663_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(KEYINPUT46), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n664_), .A2(new_n671_), .ZN(G1329gat));
  INV_X1    g471(.A(G43gat), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n424_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n666_), .A2(new_n667_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n654_), .B2(new_n424_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g477(.A(new_n654_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G50gat), .B1(new_n679_), .B2(new_n398_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n398_), .A2(G50gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n649_), .B2(new_n681_), .ZN(G1331gat));
  INV_X1    g481(.A(new_n458_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n543_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n683_), .A2(new_n684_), .A3(new_n587_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n596_), .A2(new_n685_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n686_), .A2(KEYINPUT111), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(KEYINPUT111), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT112), .B(G57gat), .Z(new_n689_));
  AND4_X1   g488(.A1(new_n590_), .A2(new_n687_), .A3(new_n688_), .A4(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n425_), .A2(new_n642_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n684_), .A2(new_n587_), .A3(new_n573_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n400_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n695_), .B1(new_n694_), .B2(new_n693_), .ZN(new_n696_));
  INV_X1    g495(.A(G57gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n696_), .A2(KEYINPUT110), .A3(new_n697_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n690_), .B1(new_n700_), .B2(new_n701_), .ZN(G1332gat));
  NAND3_X1  g501(.A1(new_n687_), .A2(new_n378_), .A3(new_n688_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT48), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(new_n704_), .A3(G64gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n703_), .B2(G64gat), .ZN(new_n706_));
  INV_X1    g505(.A(G64gat), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n378_), .A2(new_n707_), .ZN(new_n708_));
  OAI22_X1  g507(.A1(new_n705_), .A2(new_n706_), .B1(new_n693_), .B2(new_n708_), .ZN(G1333gat));
  OR3_X1    g508(.A1(new_n693_), .A2(G71gat), .A3(new_n424_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n687_), .A2(new_n259_), .A3(new_n688_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT49), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n711_), .A2(new_n712_), .A3(G71gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n711_), .B2(G71gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(G1334gat));
  OR3_X1    g514(.A1(new_n693_), .A2(G78gat), .A3(new_n624_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n687_), .A2(new_n398_), .A3(new_n688_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT50), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n717_), .A2(new_n718_), .A3(G78gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n717_), .B2(G78gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(G1335gat));
  NOR2_X1   g520(.A1(new_n684_), .A2(new_n652_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n691_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n475_), .B1(new_n723_), .B2(new_n400_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT113), .Z(new_n725_));
  NAND3_X1  g524(.A1(new_n543_), .A2(new_n457_), .A3(new_n587_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n631_), .B2(new_n640_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n728_), .A2(new_n475_), .A3(new_n400_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n725_), .A2(new_n729_), .ZN(G1336gat));
  INV_X1    g529(.A(new_n723_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G92gat), .B1(new_n731_), .B2(new_n378_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n474_), .B1(new_n369_), .B2(new_n377_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n727_), .B2(new_n733_), .ZN(G1337gat));
  NAND2_X1  g533(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n735_));
  OR2_X1    g534(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n259_), .A2(new_n471_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n723_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(G99gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n727_), .B2(new_n259_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n741_), .B2(KEYINPUT114), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n743_));
  AOI211_X1 g542(.A(new_n743_), .B(new_n740_), .C1(new_n727_), .C2(new_n259_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n735_), .B(new_n736_), .C1(new_n742_), .C2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n726_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n423_), .A2(new_n424_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n399_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n632_), .B1(new_n749_), .B2(new_n573_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n425_), .A2(KEYINPUT43), .A3(new_n630_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n259_), .B(new_n746_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G99gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n738_), .B1(new_n753_), .B2(new_n743_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n741_), .A2(KEYINPUT114), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n754_), .A2(KEYINPUT115), .A3(KEYINPUT51), .A4(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n745_), .A2(new_n756_), .ZN(G1338gat));
  NAND3_X1  g556(.A1(new_n731_), .A2(new_n470_), .A3(new_n398_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n727_), .A2(new_n398_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(G106gat), .ZN(new_n761_));
  AOI211_X1 g560(.A(KEYINPUT52), .B(new_n470_), .C1(new_n727_), .C2(new_n398_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT53), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n758_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  INV_X1    g566(.A(new_n587_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n684_), .A2(new_n458_), .A3(new_n768_), .A4(new_n630_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n769_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n588_), .A2(new_n458_), .A3(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n454_), .B1(new_n441_), .B2(new_n448_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n440_), .A2(new_n447_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n447_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n442_), .A2(new_n445_), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n453_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n777_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n538_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n516_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n518_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n526_), .A2(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(KEYINPUT55), .B(new_n520_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n535_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n535_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n784_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n573_), .B1(new_n795_), .B2(KEYINPUT58), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n782_), .B1(new_n530_), .B2(new_n536_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n535_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n535_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT58), .B(new_n799_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n573_), .B(KEYINPUT118), .C1(new_n795_), .C2(KEYINPUT58), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n798_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n455_), .A2(new_n456_), .A3(new_n538_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n794_), .B1(new_n801_), .B2(KEYINPUT117), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n787_), .A2(new_n526_), .B1(new_n785_), .B2(new_n518_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n536_), .B1(new_n807_), .B2(new_n789_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n808_), .A2(new_n809_), .A3(KEYINPUT56), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n805_), .B1(new_n806_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n539_), .A2(new_n783_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(KEYINPUT57), .A3(new_n594_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n809_), .B1(new_n808_), .B2(KEYINPUT56), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n801_), .A2(KEYINPUT117), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n794_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n818_), .A2(new_n805_), .B1(new_n539_), .B2(new_n783_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n815_), .B1(new_n819_), .B2(new_n595_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n804_), .A2(new_n814_), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n776_), .B1(new_n821_), .B2(new_n587_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n378_), .A2(new_n398_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n400_), .A2(new_n424_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT59), .B1(new_n822_), .B2(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n825_), .B(KEYINPUT120), .ZN(new_n828_));
  XOR2_X1   g627(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n813_), .A2(new_n594_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n802_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n630_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n832_), .B1(new_n835_), .B2(KEYINPUT118), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n815_), .A2(new_n831_), .B1(new_n836_), .B2(new_n798_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n768_), .B1(new_n837_), .B2(new_n814_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n830_), .B1(new_n838_), .B2(new_n776_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n827_), .A2(new_n839_), .A3(new_n683_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G113gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n821_), .A2(new_n587_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n776_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n825_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n457_), .A2(G113gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n841_), .B1(new_n845_), .B2(new_n846_), .ZN(G1340gat));
  NOR2_X1   g646(.A1(new_n822_), .A2(new_n826_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT121), .B(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n684_), .B2(KEYINPUT60), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n848_), .B(new_n850_), .C1(KEYINPUT60), .C2(new_n849_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n684_), .B1(new_n844_), .B2(new_n830_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(KEYINPUT122), .A3(new_n827_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n849_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT122), .B1(new_n852_), .B2(new_n827_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n851_), .B1(new_n855_), .B2(new_n856_), .ZN(G1341gat));
  NAND3_X1  g656(.A1(new_n827_), .A2(new_n839_), .A3(new_n768_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G127gat), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n587_), .A2(G127gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n845_), .B2(new_n860_), .ZN(G1342gat));
  INV_X1    g660(.A(G134gat), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n630_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n827_), .A2(new_n839_), .A3(new_n863_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n595_), .B(new_n825_), .C1(new_n838_), .C2(new_n776_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n862_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n864_), .A2(new_n866_), .A3(KEYINPUT123), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1343gat));
  NAND3_X1  g670(.A1(new_n590_), .A2(new_n398_), .A3(new_n424_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n378_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n642_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n543_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n875_), .A2(new_n768_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT124), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n875_), .A2(new_n883_), .A3(new_n768_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n880_), .B1(new_n882_), .B2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n875_), .B2(new_n768_), .ZN(new_n886_));
  NOR4_X1   g685(.A1(new_n822_), .A2(KEYINPUT124), .A3(new_n587_), .A4(new_n874_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n880_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n886_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n885_), .A2(new_n889_), .ZN(G1346gat));
  INV_X1    g689(.A(new_n875_), .ZN(new_n891_));
  INV_X1    g690(.A(G162gat), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n630_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n891_), .B2(new_n594_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT125), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n896_), .B(new_n892_), .C1(new_n891_), .C2(new_n594_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n893_), .B1(new_n895_), .B2(new_n897_), .ZN(G1347gat));
  AOI21_X1  g697(.A(new_n822_), .B1(new_n369_), .B2(new_n377_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n310_), .A2(new_n398_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n642_), .A3(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n901_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  AND4_X1   g702(.A1(new_n378_), .A2(new_n844_), .A3(new_n642_), .A4(new_n900_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n228_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n206_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n902_), .A2(new_n905_), .A3(new_n906_), .ZN(G1348gat));
  NAND4_X1  g706(.A1(new_n844_), .A2(new_n378_), .A3(new_n543_), .A4(new_n900_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n229_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n909_), .B1(new_n205_), .B2(new_n908_), .ZN(G1349gat));
  NAND4_X1  g709(.A1(new_n844_), .A2(new_n378_), .A3(new_n768_), .A4(new_n900_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n220_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n213_), .B2(new_n911_), .ZN(G1350gat));
  NAND2_X1  g712(.A1(new_n899_), .A2(new_n900_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G190gat), .B1(new_n914_), .B2(new_n630_), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n594_), .A2(new_n224_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n914_), .B2(new_n916_), .ZN(G1351gat));
  NOR3_X1   g716(.A1(new_n590_), .A2(new_n624_), .A3(new_n259_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n899_), .A2(new_n642_), .A3(new_n918_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g719(.A1(new_n899_), .A2(new_n918_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G204gat), .B1(new_n921_), .B2(new_n684_), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n844_), .A2(new_n378_), .A3(new_n918_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n923_), .A2(new_n315_), .A3(new_n543_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1353gat));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n926_));
  INV_X1    g725(.A(G211gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n768_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n930_));
  OR3_X1    g729(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n923_), .A2(new_n929_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n921_), .A2(new_n928_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(new_n931_), .ZN(G1354gat));
  OAI21_X1  g733(.A(G218gat), .B1(new_n921_), .B2(new_n630_), .ZN(new_n935_));
  OR2_X1    g734(.A1(new_n594_), .A2(G218gat), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n921_), .B2(new_n936_), .ZN(G1355gat));
endmodule


