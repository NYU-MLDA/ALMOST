//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  AND2_X1   g002(.A1(G228gat), .A2(G233gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT92), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n208_));
  OR2_X1    g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  OR3_X1    g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI211_X1 g016(.A(KEYINPUT87), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT86), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n212_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT86), .B1(G141gat), .B2(G148gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  AND3_X1   g023(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n219_), .A2(new_n224_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT89), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n209_), .A2(new_n207_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT88), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n209_), .A2(KEYINPUT88), .A3(new_n207_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n228_), .A2(new_n229_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n229_), .B1(new_n228_), .B2(new_n234_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n214_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT29), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G197gat), .B(G204gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT21), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G211gat), .B(G218gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT91), .ZN(new_n245_));
  INV_X1    g044(.A(G197gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(G204gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT21), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n248_), .B1(KEYINPUT91), .B2(new_n239_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G197gat), .B(G204gat), .Z(new_n250_));
  OAI21_X1  g049(.A(new_n242_), .B1(new_n250_), .B2(KEYINPUT21), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n244_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n204_), .A2(KEYINPUT92), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n206_), .B1(new_n238_), .B2(new_n255_), .ZN(new_n256_));
  AOI211_X1 g055(.A(new_n254_), .B(new_n205_), .C1(new_n237_), .C2(KEYINPUT29), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n203_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT93), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n228_), .A2(new_n234_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT89), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n228_), .A2(new_n234_), .A3(new_n229_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n261_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT29), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n255_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n205_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n238_), .A2(new_n255_), .A3(new_n206_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(new_n202_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT94), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n268_), .A2(KEYINPUT94), .A3(new_n269_), .A4(new_n202_), .ZN(new_n273_));
  OAI211_X1 g072(.A(KEYINPUT93), .B(new_n203_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n260_), .A2(new_n272_), .A3(new_n273_), .A4(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G22gat), .B(G50gat), .Z(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n266_), .B(new_n214_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n281_), .A2(new_n278_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n277_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n265_), .A2(new_n266_), .A3(new_n279_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n278_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n285_), .A3(new_n276_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n275_), .A2(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n287_), .A2(new_n258_), .A3(new_n270_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT95), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT95), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n289_), .A2(new_n294_), .A3(new_n291_), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT104), .B(KEYINPUT27), .Z(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR3_X1   g096(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT25), .B(G183gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G190gat), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT24), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n309_), .A2(KEYINPUT96), .ZN(new_n310_));
  INV_X1    g109(.A(G169gat), .ZN(new_n311_));
  INV_X1    g110(.A(G176gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n312_), .A3(KEYINPUT82), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT82), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(G169gat), .B2(G176gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT96), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(new_n308_), .B2(KEYINPUT24), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n310_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n307_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT22), .B(G169gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n312_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n308_), .B(KEYINPUT97), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT98), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n306_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n304_), .A2(new_n305_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT98), .B1(new_n329_), .B2(new_n326_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n324_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n252_), .B1(new_n320_), .B2(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT81), .B(G190gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n306_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT84), .ZN(new_n338_));
  AOI21_X1  g137(.A(G176gat), .B1(new_n338_), .B2(KEYINPUT22), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(G169gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT83), .B1(new_n316_), .B2(new_n309_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n309_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT83), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(new_n313_), .A4(new_n315_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT24), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n329_), .B1(new_n348_), .B2(new_n316_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT25), .B1(new_n333_), .B2(new_n334_), .ZN(new_n350_));
  OR2_X1    g149(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n353_), .B1(new_n336_), .B2(KEYINPUT26), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n349_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n341_), .B1(new_n347_), .B2(new_n355_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n332_), .B(KEYINPUT20), .C1(new_n252_), .C2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT19), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT99), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n336_), .A2(KEYINPUT26), .ZN(new_n362_));
  INV_X1    g161(.A(new_n353_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n362_), .A2(new_n363_), .B1(new_n351_), .B2(new_n350_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n313_), .A2(new_n315_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n306_), .B1(new_n365_), .B2(KEYINPUT24), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n367_), .A2(new_n346_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n243_), .B1(new_n240_), .B2(new_n239_), .ZN(new_n369_));
  OAI211_X1 g168(.A(KEYINPUT21), .B(new_n247_), .C1(new_n250_), .C2(new_n245_), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n369_), .A2(new_n370_), .B1(new_n243_), .B2(new_n241_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n361_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n356_), .A2(KEYINPUT99), .A3(new_n252_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(KEYINPUT20), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n328_), .A2(new_n330_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n324_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n316_), .A2(new_n318_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n306_), .B(new_n301_), .C1(new_n378_), .C2(new_n310_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n371_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT100), .ZN(new_n381_));
  INV_X1    g180(.A(new_n359_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT100), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n377_), .A2(new_n371_), .A3(new_n383_), .A4(new_n379_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n360_), .B1(new_n374_), .B2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G8gat), .B(G36gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT18), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT20), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n346_), .B(new_n349_), .C1(new_n354_), .C2(new_n352_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n371_), .B1(new_n394_), .B2(new_n341_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n393_), .B1(new_n395_), .B2(KEYINPUT99), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n384_), .A2(new_n382_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n372_), .A4(new_n381_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n390_), .B1(new_n398_), .B2(new_n360_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n297_), .B1(new_n392_), .B2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n360_), .A3(new_n390_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n357_), .A2(new_n359_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT102), .B1(new_n320_), .B2(new_n331_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT102), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n377_), .A2(new_n404_), .A3(new_n379_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n405_), .A3(new_n371_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n396_), .A2(new_n372_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n402_), .B1(new_n407_), .B2(new_n359_), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n390_), .B(KEYINPUT103), .Z(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT27), .B(new_n401_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n400_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G127gat), .B(G134gat), .Z(new_n412_));
  XOR2_X1   g211(.A(G113gat), .B(G120gat), .Z(new_n413_));
  XOR2_X1   g212(.A(new_n412_), .B(new_n413_), .Z(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G71gat), .B(G99gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(G43gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n356_), .B(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419_));
  INV_X1    g218(.A(G15gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT30), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT31), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n418_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n368_), .A2(new_n417_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n368_), .A2(new_n417_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT85), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n424_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n429_), .B1(new_n424_), .B2(new_n428_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n415_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n432_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(new_n414_), .A3(new_n430_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G1gat), .B(G29gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(G85gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT0), .B(G57gat), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n438_), .B(new_n439_), .Z(new_n440_));
  NAND2_X1  g239(.A1(G225gat), .A2(G233gat), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n237_), .A2(KEYINPUT101), .A3(new_n415_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT101), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n414_), .B1(new_n265_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT4), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n265_), .A2(KEYINPUT4), .A3(new_n415_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n441_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n415_), .B1(new_n237_), .B2(KEYINPUT101), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n265_), .A2(new_n443_), .A3(new_n414_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n441_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n440_), .B1(new_n448_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n440_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n450_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n446_), .B1(new_n455_), .B2(KEYINPUT4), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n451_), .B(new_n454_), .C1(new_n456_), .C2(new_n441_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n436_), .A2(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n293_), .A2(new_n295_), .A3(new_n411_), .A4(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n436_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n293_), .A2(new_n295_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n458_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n411_), .A2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n462_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n390_), .A2(KEYINPUT32), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n398_), .A2(new_n360_), .A3(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n408_), .B2(new_n467_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(new_n453_), .B2(new_n457_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n451_), .B1(new_n456_), .B2(new_n441_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT33), .B1(new_n471_), .B2(new_n440_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n386_), .A2(new_n391_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n441_), .ZN(new_n474_));
  AOI211_X1 g273(.A(new_n474_), .B(new_n446_), .C1(new_n455_), .C2(KEYINPUT4), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n455_), .A2(new_n474_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n454_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n473_), .B(new_n401_), .C1(new_n475_), .C2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n472_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n471_), .A2(KEYINPUT33), .A3(new_n440_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n470_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n461_), .B1(new_n466_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT75), .B(G15gat), .ZN(new_n486_));
  INV_X1    g285(.A(G22gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(KEYINPUT75), .A2(G15gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(KEYINPUT75), .A2(G15gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(G22gat), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(G1gat), .ZN(new_n493_));
  INV_X1    g292(.A(G8gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT14), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G1gat), .B(G8gat), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n497_), .A2(KEYINPUT76), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(KEYINPUT76), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n492_), .A2(new_n498_), .A3(new_n495_), .A4(new_n499_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G29gat), .B(G36gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT77), .ZN(new_n510_));
  AOI211_X1 g309(.A(new_n510_), .B(new_n508_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT77), .B1(new_n503_), .B2(new_n507_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n485_), .B(new_n509_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n502_), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n492_), .A2(new_n495_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n507_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n510_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n503_), .A2(KEYINPUT77), .A3(new_n507_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n507_), .B(new_n519_), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n517_), .A2(new_n518_), .B1(new_n504_), .B2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n513_), .B1(new_n521_), .B2(new_n485_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G113gat), .B(G141gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G169gat), .B(G197gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  NOR2_X1   g324(.A1(new_n525_), .A2(KEYINPUT78), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n522_), .B(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n527_), .B(KEYINPUT79), .Z(new_n528_));
  NOR2_X1   g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(G85gat), .A2(G92gat), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(new_n529_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT9), .B1(new_n532_), .B2(KEYINPUT65), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT65), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535_));
  NOR4_X1   g334(.A1(new_n531_), .A2(new_n529_), .A3(new_n534_), .A4(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n530_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT66), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT66), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n539_), .B(new_n530_), .C1(new_n533_), .C2(new_n536_), .ZN(new_n540_));
  OR2_X1    g339(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT64), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT64), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n545_), .A3(new_n542_), .ZN(new_n546_));
  AOI21_X1  g345(.A(G106gat), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G99gat), .A2(G106gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT6), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT6), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(G99gat), .A3(G106gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT67), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n549_), .A2(new_n551_), .A3(KEYINPUT67), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n547_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n538_), .A2(new_n540_), .A3(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n531_), .A2(new_n529_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n559_), .B1(new_n563_), .B2(new_n552_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT8), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT69), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n549_), .A2(new_n551_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT7), .ZN(new_n568_));
  INV_X1    g367(.A(G99gat), .ZN(new_n569_));
  INV_X1    g368(.A(G106gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n560_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n532_), .B1(new_n567_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT69), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n574_), .A3(KEYINPUT8), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n554_), .A2(new_n555_), .A3(new_n563_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT68), .B(KEYINPUT8), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n559_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n566_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G57gat), .B(G64gat), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n581_), .A2(KEYINPUT11), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(KEYINPUT11), .ZN(new_n583_));
  XOR2_X1   g382(.A(G71gat), .B(G78gat), .Z(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n583_), .A2(new_n584_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n558_), .A2(new_n580_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n587_), .B1(new_n558_), .B2(new_n580_), .ZN(new_n590_));
  OAI211_X1 g389(.A(G230gat), .B(G233gat), .C1(new_n589_), .C2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT5), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G176gat), .B(G204gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n593_), .B(new_n594_), .Z(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT70), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G230gat), .A2(G233gat), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n588_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n558_), .A2(new_n580_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n587_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n600_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  AOI211_X1 g402(.A(KEYINPUT12), .B(new_n587_), .C1(new_n558_), .C2(new_n580_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n599_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n597_), .B1(new_n588_), .B2(new_n598_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n591_), .B(new_n596_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT71), .ZN(new_n608_));
  INV_X1    g407(.A(new_n606_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n609_), .B(new_n599_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT71), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n610_), .A2(new_n611_), .A3(new_n591_), .A4(new_n596_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n610_), .A2(new_n591_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n595_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n613_), .A2(new_n615_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n620_));
  OAI21_X1  g419(.A(new_n617_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n587_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(new_n504_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT17), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G127gat), .B(G155gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT16), .ZN(new_n628_));
  XOR2_X1   g427(.A(G183gat), .B(G211gat), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  OR3_X1    g429(.A1(new_n625_), .A2(new_n626_), .A3(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(KEYINPUT17), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n625_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT74), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n601_), .A2(new_n520_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(G232gat), .A2(G233gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT34), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n638_), .A2(KEYINPUT35), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n558_), .A2(new_n580_), .A3(new_n507_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(KEYINPUT35), .A3(new_n638_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n638_), .A2(KEYINPUT35), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n636_), .A2(new_n643_), .A3(new_n639_), .A4(new_n640_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n635_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(G190gat), .B(G218gat), .Z(new_n646_));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT36), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n649_), .A2(KEYINPUT36), .ZN(new_n652_));
  OR3_X1    g451(.A1(new_n645_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n645_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(KEYINPUT37), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT37), .ZN(new_n656_));
  INV_X1    g455(.A(new_n654_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n645_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n656_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n634_), .B1(new_n655_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR4_X1   g460(.A1(new_n483_), .A2(new_n528_), .A3(new_n622_), .A4(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n493_), .A3(new_n458_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n664_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n294_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n667_));
  AOI211_X1 g466(.A(KEYINPUT95), .B(new_n290_), .C1(new_n275_), .C2(new_n288_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n465_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n482_), .A2(new_n436_), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n460_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n622_), .A2(new_n527_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n634_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n657_), .A2(new_n658_), .ZN(new_n674_));
  AND4_X1   g473(.A1(new_n671_), .A2(new_n672_), .A3(new_n673_), .A4(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(new_n458_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n665_), .B(new_n666_), .C1(new_n493_), .C2(new_n676_), .ZN(G1324gat));
  INV_X1    g476(.A(new_n411_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n662_), .A2(new_n494_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n675_), .A2(new_n678_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G8gat), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n681_), .A2(KEYINPUT39), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(KEYINPUT39), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n679_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT40), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT40), .B(new_n679_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1325gat));
  INV_X1    g487(.A(new_n675_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G15gat), .B1(new_n689_), .B2(new_n436_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT106), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n690_), .A2(KEYINPUT106), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n690_), .A2(KEYINPUT106), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(KEYINPUT41), .A3(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n662_), .A2(new_n420_), .A3(new_n462_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n693_), .A2(new_n696_), .A3(new_n697_), .ZN(G1326gat));
  NAND3_X1  g497(.A1(new_n662_), .A2(new_n487_), .A3(new_n463_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n675_), .A2(new_n463_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G22gat), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT42), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(KEYINPUT42), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT107), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n706_), .B(new_n699_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1327gat));
  INV_X1    g507(.A(new_n674_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n621_), .A2(new_n634_), .A3(new_n709_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n483_), .A2(new_n528_), .A3(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G29gat), .B1(new_n711_), .B2(new_n458_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n672_), .A2(new_n634_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n655_), .A2(new_n659_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n718_), .B1(new_n671_), .B2(new_n720_), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n719_), .B(new_n716_), .C1(new_n670_), .C2(new_n460_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT44), .B(new_n714_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n671_), .A2(new_n720_), .A3(new_n715_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n719_), .B1(new_n670_), .B2(new_n460_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(new_n718_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n728_), .A2(KEYINPUT109), .A3(KEYINPUT44), .A4(new_n714_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n725_), .A2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n714_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n458_), .A2(G29gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n712_), .B1(new_n735_), .B2(new_n736_), .ZN(G1328gat));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738_));
  INV_X1    g537(.A(G36gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n411_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n730_), .B2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n711_), .A2(new_n739_), .A3(new_n678_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n742_), .A2(KEYINPUT45), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(KEYINPUT45), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n738_), .B1(new_n741_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n744_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n718_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(new_n483_), .B2(new_n719_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n713_), .B1(new_n749_), .B2(new_n726_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n678_), .B1(new_n750_), .B2(KEYINPUT44), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n725_), .B2(new_n729_), .ZN(new_n752_));
  OAI211_X1 g551(.A(KEYINPUT46), .B(new_n747_), .C1(new_n752_), .C2(new_n739_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n746_), .A2(new_n753_), .ZN(G1329gat));
  NAND2_X1  g553(.A1(new_n462_), .A2(G43gat), .ZN(new_n755_));
  AOI221_X4 g554(.A(new_n755_), .B1(new_n732_), .B2(new_n731_), .C1(new_n725_), .C2(new_n729_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n711_), .A2(new_n462_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(G43gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT47), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760_));
  INV_X1    g559(.A(new_n758_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n760_), .B(new_n761_), .C1(new_n734_), .C2(new_n755_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n762_), .ZN(G1330gat));
  INV_X1    g562(.A(new_n463_), .ZN(new_n764_));
  OAI21_X1  g563(.A(G50gat), .B1(new_n734_), .B2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(G50gat), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT110), .Z(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n711_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n765_), .A2(new_n768_), .ZN(G1331gat));
  XOR2_X1   g568(.A(new_n522_), .B(new_n526_), .Z(new_n770_));
  NOR4_X1   g569(.A1(new_n483_), .A2(new_n770_), .A3(new_n621_), .A4(new_n661_), .ZN(new_n771_));
  AOI21_X1  g570(.A(G57gat), .B1(new_n771_), .B2(new_n458_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n671_), .A2(new_n674_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n528_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n621_), .A2(new_n775_), .A3(new_n634_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n464_), .A2(KEYINPUT111), .ZN(new_n779_));
  MUX2_X1   g578(.A(KEYINPUT111), .B(new_n779_), .S(G57gat), .Z(new_n780_));
  AOI21_X1  g579(.A(new_n772_), .B1(new_n778_), .B2(new_n780_), .ZN(G1332gat));
  OAI21_X1  g580(.A(G64gat), .B1(new_n777_), .B2(new_n411_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT48), .ZN(new_n783_));
  INV_X1    g582(.A(G64gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n771_), .A2(new_n784_), .A3(new_n678_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1333gat));
  OAI21_X1  g585(.A(G71gat), .B1(new_n777_), .B2(new_n436_), .ZN(new_n787_));
  XOR2_X1   g586(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(G71gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n771_), .A2(new_n790_), .A3(new_n462_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1334gat));
  INV_X1    g591(.A(G78gat), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n771_), .A2(new_n793_), .A3(new_n463_), .ZN(new_n794_));
  OAI21_X1  g593(.A(G78gat), .B1(new_n777_), .B2(new_n764_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n795_), .A2(KEYINPUT50), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(KEYINPUT50), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n794_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT113), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n800_), .B(new_n794_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1335gat));
  NAND2_X1  g601(.A1(new_n622_), .A2(new_n634_), .ZN(new_n803_));
  NOR4_X1   g602(.A1(new_n483_), .A2(new_n803_), .A3(new_n770_), .A4(new_n674_), .ZN(new_n804_));
  INV_X1    g603(.A(G85gat), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n458_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n803_), .A2(new_n770_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n728_), .A2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT114), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n809_), .A2(new_n458_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n806_), .B1(new_n810_), .B2(new_n805_), .ZN(G1336gat));
  INV_X1    g610(.A(G92gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n804_), .A2(new_n812_), .A3(new_n678_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n809_), .A2(new_n678_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n812_), .ZN(G1337gat));
  NAND3_X1  g614(.A1(new_n728_), .A2(new_n462_), .A3(new_n807_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n436_), .B1(new_n546_), .B2(new_n544_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n816_), .A2(G99gat), .B1(new_n804_), .B2(new_n817_), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g618(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n463_), .B(new_n807_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(G106gat), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(new_n821_), .A3(G106gat), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n804_), .A2(new_n570_), .A3(new_n463_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n820_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n825_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n827_), .B(new_n820_), .C1(new_n829_), .C2(new_n823_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n828_), .A2(new_n831_), .ZN(G1339gat));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n590_), .B(new_n600_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n836_), .A2(KEYINPUT55), .A3(new_n609_), .A4(new_n599_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n588_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(G230gat), .A3(G233gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n835_), .A2(new_n837_), .A3(new_n839_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n840_), .A2(KEYINPUT56), .A3(new_n595_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT56), .B1(new_n840_), .B2(new_n595_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n841_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n840_), .A2(new_n595_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT56), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n843_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n504_), .A2(new_n520_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n485_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n484_), .B(new_n509_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n525_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n525_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n484_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n513_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT117), .B1(new_n852_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n850_), .A2(new_n851_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n853_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n522_), .A2(new_n525_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n856_), .A2(new_n861_), .B1(new_n608_), .B2(new_n612_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n847_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n833_), .B1(new_n844_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n845_), .A2(new_n846_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n840_), .A2(KEYINPUT56), .A3(new_n595_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(KEYINPUT118), .A3(new_n866_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n867_), .A2(KEYINPUT58), .A3(new_n847_), .A4(new_n862_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n864_), .A2(new_n720_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n613_), .A2(new_n615_), .B1(new_n856_), .B2(new_n861_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n613_), .A2(new_n770_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n840_), .A2(new_n595_), .B1(new_n873_), .B2(new_n846_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n840_), .A2(new_n873_), .A3(new_n846_), .A4(new_n595_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n871_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n870_), .B1(new_n877_), .B2(new_n709_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n845_), .B1(KEYINPUT116), .B2(KEYINPUT56), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n879_), .A2(new_n770_), .A3(new_n613_), .A4(new_n876_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n871_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(KEYINPUT57), .A3(new_n674_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n869_), .A2(new_n878_), .A3(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n634_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n660_), .A2(new_n621_), .A3(new_n528_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT54), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  NOR4_X1   g687(.A1(new_n463_), .A2(new_n678_), .A3(new_n464_), .A4(new_n436_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT59), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n884_), .A2(new_n892_), .A3(new_n634_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(new_n884_), .B2(new_n634_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n887_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n889_), .A2(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n891_), .B1(new_n897_), .B2(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G113gat), .B1(new_n900_), .B2(new_n528_), .ZN(new_n901_));
  OR3_X1    g700(.A1(new_n890_), .A2(G113gat), .A3(new_n527_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1340gat));
  OAI21_X1  g702(.A(G120gat), .B1(new_n900_), .B2(new_n621_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n890_), .ZN(new_n905_));
  INV_X1    g704(.A(G120gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(new_n621_), .B2(KEYINPUT60), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n905_), .B(new_n907_), .C1(KEYINPUT60), .C2(new_n906_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n904_), .A2(new_n908_), .ZN(G1341gat));
  OAI21_X1  g708(.A(G127gat), .B1(new_n900_), .B2(new_n634_), .ZN(new_n910_));
  OR3_X1    g709(.A1(new_n890_), .A2(G127gat), .A3(new_n634_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1342gat));
  OAI21_X1  g711(.A(G134gat), .B1(new_n900_), .B2(new_n719_), .ZN(new_n913_));
  OR3_X1    g712(.A1(new_n890_), .A2(G134gat), .A3(new_n674_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1343gat));
  NOR4_X1   g714(.A1(new_n764_), .A2(new_n678_), .A3(new_n464_), .A4(new_n462_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n888_), .A2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n770_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n622_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g721(.A1(new_n917_), .A2(new_n634_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT61), .B(G155gat), .Z(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1346gat));
  OAI21_X1  g724(.A(G162gat), .B1(new_n917_), .B2(new_n719_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n674_), .A2(G162gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n917_), .B2(new_n927_), .ZN(G1347gat));
  NAND2_X1  g727(.A1(new_n678_), .A2(new_n459_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n463_), .A2(new_n929_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n896_), .A2(new_n770_), .A3(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(G169gat), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n930_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n885_), .A2(KEYINPUT119), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n893_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n935_), .B1(new_n937_), .B2(new_n887_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n938_), .A2(new_n321_), .A3(new_n770_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n931_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n934_), .A2(new_n939_), .A3(new_n940_), .ZN(G1348gat));
  AOI21_X1  g740(.A(G176gat), .B1(new_n938_), .B2(new_n622_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n463_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n929_), .A2(new_n312_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n943_), .A2(new_n622_), .A3(new_n944_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  OAI21_X1  g745(.A(KEYINPUT120), .B1(new_n942_), .B2(new_n946_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n896_), .A2(new_n622_), .A3(new_n930_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(new_n312_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT120), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n949_), .A2(new_n950_), .A3(new_n945_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n947_), .A2(new_n951_), .ZN(G1349gat));
  NOR2_X1   g751(.A1(new_n929_), .A2(new_n634_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n335_), .B1(new_n943_), .B2(new_n953_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n634_), .A2(new_n299_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n954_), .B1(new_n938_), .B2(new_n955_), .ZN(G1350gat));
  NAND2_X1  g755(.A1(new_n938_), .A2(new_n720_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(G190gat), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n938_), .A2(new_n300_), .A3(new_n709_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1351gat));
  NAND4_X1  g759(.A1(new_n463_), .A2(new_n678_), .A3(new_n464_), .A4(new_n436_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n961_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(new_n770_), .ZN(new_n963_));
  XOR2_X1   g762(.A(KEYINPUT121), .B(G197gat), .Z(new_n964_));
  XNOR2_X1  g763(.A(new_n963_), .B(new_n964_), .ZN(G1352gat));
  NAND2_X1  g764(.A1(new_n962_), .A2(new_n622_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g766(.A(new_n961_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n888_), .A2(new_n968_), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n634_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n970_), .B(KEYINPUT122), .ZN(new_n971_));
  OR3_X1    g770(.A1(new_n969_), .A2(KEYINPUT123), .A3(new_n971_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n973_));
  OAI21_X1  g772(.A(KEYINPUT123), .B1(new_n969_), .B2(new_n971_), .ZN(new_n974_));
  AND3_X1   g773(.A1(new_n972_), .A2(new_n973_), .A3(new_n974_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n973_), .B1(new_n972_), .B2(new_n974_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n975_), .A2(new_n976_), .ZN(G1354gat));
  XOR2_X1   g776(.A(KEYINPUT125), .B(G218gat), .Z(new_n978_));
  AND3_X1   g777(.A1(new_n962_), .A2(KEYINPUT124), .A3(new_n709_), .ZN(new_n979_));
  AOI21_X1  g778(.A(KEYINPUT124), .B1(new_n962_), .B2(new_n709_), .ZN(new_n980_));
  OAI21_X1  g779(.A(new_n978_), .B1(new_n979_), .B2(new_n980_), .ZN(new_n981_));
  INV_X1    g780(.A(new_n978_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n720_), .A2(new_n982_), .ZN(new_n983_));
  OAI211_X1 g782(.A(new_n981_), .B(KEYINPUT126), .C1(new_n969_), .C2(new_n983_), .ZN(new_n984_));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n888_), .A2(new_n709_), .A3(new_n968_), .ZN(new_n986_));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n986_), .A2(new_n987_), .ZN(new_n988_));
  NAND3_X1  g787(.A1(new_n962_), .A2(KEYINPUT124), .A3(new_n709_), .ZN(new_n989_));
  AOI21_X1  g788(.A(new_n982_), .B1(new_n988_), .B2(new_n989_), .ZN(new_n990_));
  NOR2_X1   g789(.A1(new_n969_), .A2(new_n983_), .ZN(new_n991_));
  OAI21_X1  g790(.A(new_n985_), .B1(new_n990_), .B2(new_n991_), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n984_), .A2(new_n992_), .ZN(G1355gat));
endmodule


