//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G8gat), .B(G36gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G64gat), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n206_), .A2(G92gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(G92gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT93), .ZN(new_n211_));
  INV_X1    g010(.A(G197gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT88), .B1(new_n212_), .B2(G204gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT88), .ZN(new_n214_));
  INV_X1    g013(.A(G204gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(G197gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(G204gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT21), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT89), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(new_n212_), .B2(G204gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n215_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT21), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .A4(new_n217_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G211gat), .B(G218gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n219_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n223_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n221_), .A2(new_n217_), .A3(new_n222_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT76), .ZN(new_n230_));
  INV_X1    g029(.A(G183gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(KEYINPUT25), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT25), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(G183gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n230_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT26), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT26), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G190gat), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT76), .B1(new_n231_), .B2(KEYINPUT25), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n235_), .A2(KEYINPUT77), .A3(new_n240_), .A4(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT77), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n233_), .A2(G183gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n231_), .A2(KEYINPUT25), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT76), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n243_), .B1(new_n244_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT23), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT23), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(G183gat), .A3(G190gat), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT24), .ZN(new_n254_));
  INV_X1    g053(.A(G169gat), .ZN(new_n255_));
  INV_X1    g054(.A(G176gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT24), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n257_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n253_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n242_), .A2(new_n248_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n231_), .A2(new_n236_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT80), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n265_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT80), .B1(new_n249_), .B2(KEYINPUT23), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n264_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT22), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G169gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(G176gat), .B1(new_n270_), .B2(KEYINPUT79), .ZN(new_n271_));
  OR3_X1    g070(.A1(new_n255_), .A2(KEYINPUT79), .A3(KEYINPUT22), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT78), .B(G169gat), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n271_), .B(new_n272_), .C1(new_n269_), .C2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n268_), .A2(new_n258_), .A3(new_n274_), .ZN(new_n275_));
  AOI221_X4 g074(.A(KEYINPUT91), .B1(new_n226_), .B2(new_n229_), .C1(new_n263_), .C2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT91), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n263_), .A2(new_n275_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n226_), .A2(new_n229_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT20), .B1(new_n276_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT92), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n255_), .A2(KEYINPUT22), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n270_), .A2(new_n283_), .A3(new_n256_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n284_), .A2(new_n258_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n250_), .A2(new_n252_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n264_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n245_), .A2(new_n246_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n237_), .A2(new_n239_), .ZN(new_n290_));
  OAI221_X1 g089(.A(new_n257_), .B1(new_n260_), .B2(new_n259_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n266_), .A2(new_n267_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n288_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n282_), .B1(new_n293_), .B2(new_n279_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n289_), .A2(new_n290_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(new_n261_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n266_), .A2(new_n267_), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n296_), .A2(new_n297_), .B1(new_n287_), .B2(new_n285_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n224_), .A2(new_n225_), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n299_), .A2(new_n219_), .B1(new_n228_), .B2(new_n227_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n300_), .A3(KEYINPUT92), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n294_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G226gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT19), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n211_), .B1(new_n281_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n278_), .A2(new_n279_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT91), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n278_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n304_), .B1(new_n294_), .B2(new_n301_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n311_), .A2(KEYINPUT93), .A3(KEYINPUT20), .A4(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n307_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT20), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n315_), .B1(new_n293_), .B2(new_n279_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n300_), .A2(new_n275_), .A3(new_n263_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n304_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n210_), .B1(new_n314_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n319_), .ZN(new_n321_));
  AOI211_X1 g120(.A(new_n321_), .B(new_n209_), .C1(new_n307_), .C2(new_n313_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n203_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n314_), .A2(new_n319_), .A3(new_n210_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT95), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n298_), .A2(new_n300_), .ZN(new_n326_));
  OAI211_X1 g125(.A(KEYINPUT20), .B(new_n326_), .C1(new_n276_), .C2(new_n280_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n304_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n318_), .A2(new_n304_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n325_), .B1(new_n331_), .B2(new_n209_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n329_), .B1(new_n327_), .B2(new_n304_), .ZN(new_n333_));
  NOR3_X1   g132(.A1(new_n333_), .A2(KEYINPUT95), .A3(new_n210_), .ZN(new_n334_));
  OAI211_X1 g133(.A(KEYINPUT27), .B(new_n324_), .C1(new_n332_), .C2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G225gat), .A2(G233gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G155gat), .B(G162gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n340_));
  INV_X1    g139(.A(G141gat), .ZN(new_n341_));
  INV_X1    g140(.A(G148gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT85), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n343_), .B(new_n344_), .C1(new_n346_), .C2(KEYINPUT3), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n346_), .A2(KEYINPUT3), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n339_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G141gat), .B(G148gat), .Z(new_n350_));
  NAND3_X1  g149(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n350_), .B(new_n351_), .C1(KEYINPUT1), .C2(new_n338_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT86), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT86), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n349_), .A2(new_n355_), .A3(new_n352_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G127gat), .B(G134gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G113gat), .B(G120gat), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT82), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n358_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n357_), .A2(new_n358_), .A3(KEYINPUT82), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n354_), .A2(new_n356_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n359_), .A2(new_n361_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n349_), .A3(new_n352_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n349_), .A2(new_n355_), .A3(new_n352_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n355_), .B1(new_n349_), .B2(new_n352_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n370_), .B1(new_n373_), .B2(new_n364_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n337_), .B(new_n367_), .C1(new_n374_), .C2(new_n366_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n365_), .A2(new_n369_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n336_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT0), .ZN(new_n380_));
  INV_X1    g179(.A(G57gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G85gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n378_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n375_), .A2(new_n384_), .A3(new_n377_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n323_), .A2(new_n335_), .A3(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n373_), .A2(KEYINPUT87), .A3(KEYINPUT29), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n354_), .A2(KEYINPUT29), .A3(new_n356_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G228gat), .A2(G233gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n279_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n353_), .A2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n396_), .B1(new_n401_), .B2(new_n279_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G22gat), .B(G50gat), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n404_), .B(KEYINPUT28), .Z(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n399_), .A2(new_n403_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n397_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n405_), .B1(new_n408_), .B2(new_n402_), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n373_), .A2(KEYINPUT29), .ZN(new_n410_));
  XOR2_X1   g209(.A(G78gat), .B(G106gat), .Z(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n407_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n412_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n364_), .B(KEYINPUT31), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n263_), .A2(new_n275_), .A3(KEYINPUT30), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT30), .B1(new_n263_), .B2(new_n275_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G15gat), .B(G43gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G71gat), .B(G99gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n418_), .A2(new_n419_), .A3(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n422_), .A2(new_n423_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n422_), .A2(new_n423_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT30), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n278_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n263_), .A2(new_n275_), .A3(KEYINPUT30), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n428_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n417_), .A2(new_n425_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT81), .B1(new_n425_), .B2(new_n432_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n424_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n430_), .A2(new_n431_), .A3(new_n428_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n416_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT83), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n434_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AOI211_X1 g241(.A(KEYINPUT83), .B(new_n416_), .C1(new_n435_), .C2(new_n439_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n442_), .A2(KEYINPUT84), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n438_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n417_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n433_), .B1(new_n448_), .B2(KEYINPUT83), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n440_), .A2(new_n441_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n445_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n415_), .B1(new_n444_), .B2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT84), .B1(new_n442_), .B2(new_n443_), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n410_), .B(new_n411_), .Z(new_n454_));
  AOI21_X1  g253(.A(new_n406_), .B1(new_n399_), .B2(new_n403_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n408_), .A2(new_n402_), .A3(new_n405_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n407_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n449_), .A2(new_n445_), .A3(new_n450_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n453_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n390_), .B1(new_n452_), .B2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n366_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT4), .B1(new_n373_), .B2(new_n364_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n336_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n465_), .B(new_n384_), .C1(new_n376_), .C2(new_n336_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n384_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(KEYINPUT33), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT33), .ZN(new_n469_));
  AOI211_X1 g268(.A(new_n469_), .B(new_n384_), .C1(new_n375_), .C2(new_n377_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n320_), .A2(new_n322_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n207_), .A2(KEYINPUT32), .A3(new_n208_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT94), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(new_n319_), .A3(new_n314_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n386_), .A2(new_n387_), .B1(new_n331_), .B2(new_n473_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n471_), .A2(new_n472_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n415_), .A2(new_n453_), .A3(new_n460_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n462_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT7), .ZN(new_n481_));
  INV_X1    g280(.A(G99gat), .ZN(new_n482_));
  INV_X1    g281(.A(G106gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G99gat), .A2(G106gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n484_), .A2(new_n487_), .A3(new_n488_), .A4(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G85gat), .B(G92gat), .Z(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT8), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT8), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n490_), .A2(new_n494_), .A3(new_n491_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT64), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G85gat), .A2(G92gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT9), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n500_), .B1(new_n491_), .B2(new_n499_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT10), .B(G99gat), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n483_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n497_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n487_), .A2(new_n488_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n501_), .A2(new_n503_), .A3(new_n504_), .A4(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n496_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G43gat), .B(G50gat), .Z(new_n509_));
  XNOR2_X1  g308(.A(G29gat), .B(G36gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT35), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G232gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT34), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n508_), .A2(new_n513_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n513_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT67), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n493_), .A2(new_n521_), .A3(new_n495_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n506_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n518_), .B1(new_n520_), .B2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n517_), .A2(new_n514_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G190gat), .B(G218gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G134gat), .B(G162gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(KEYINPUT36), .ZN(new_n532_));
  INV_X1    g331(.A(new_n527_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n533_), .B(new_n518_), .C1(new_n520_), .C2(new_n525_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n528_), .A2(new_n532_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n531_), .B(KEYINPUT36), .Z(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n538_), .B1(new_n528_), .B2(new_n534_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n540_), .A2(KEYINPUT96), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(KEYINPUT96), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n480_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT97), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT66), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT11), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n381_), .A2(G64gat), .ZN(new_n548_));
  INV_X1    g347(.A(G64gat), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(G57gat), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n547_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G71gat), .B(G78gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT65), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n549_), .A2(G57gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n381_), .A2(G64gat), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT11), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT65), .B1(new_n558_), .B2(new_n552_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n556_), .A2(new_n557_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(new_n547_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n555_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n546_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n554_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n558_), .A2(KEYINPUT65), .A3(new_n552_), .ZN(new_n566_));
  OAI22_X1  g365(.A1(new_n565_), .A2(new_n566_), .B1(new_n547_), .B2(new_n560_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n555_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(KEYINPUT66), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n508_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n564_), .A2(new_n569_), .A3(new_n507_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(G230gat), .A3(G233gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT68), .B(KEYINPUT12), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G230gat), .A2(G233gat), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n567_), .A2(KEYINPUT12), .A3(new_n568_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n524_), .A2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n576_), .A2(new_n571_), .A3(new_n577_), .A4(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n574_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(new_n215_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT5), .B(G176gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n574_), .A2(new_n580_), .A3(new_n585_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n589_), .B1(new_n592_), .B2(new_n590_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT17), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G127gat), .B(G155gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT16), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(G183gat), .ZN(new_n599_));
  INV_X1    g398(.A(G211gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G15gat), .B(G22gat), .ZN(new_n602_));
  INV_X1    g401(.A(G8gat), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G1gat), .B(G8gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT72), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n607_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT73), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n562_), .A2(new_n563_), .ZN(new_n612_));
  AOI211_X1 g411(.A(new_n596_), .B(new_n601_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n613_), .B1(new_n612_), .B2(new_n611_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n601_), .B(KEYINPUT17), .ZN(new_n615_));
  INV_X1    g414(.A(new_n570_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n610_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(new_n610_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n614_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n513_), .B(KEYINPUT15), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(new_n607_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G229gat), .A2(G233gat), .ZN(new_n623_));
  INV_X1    g422(.A(new_n607_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n513_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n622_), .A2(new_n623_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n513_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n607_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(KEYINPUT74), .A3(new_n625_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n623_), .ZN(new_n630_));
  OR3_X1    g429(.A1(new_n513_), .A2(KEYINPUT74), .A3(new_n624_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n629_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n626_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G169gat), .B(G197gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT75), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G113gat), .B(G141gat), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n635_), .B(new_n636_), .Z(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n633_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n626_), .A2(new_n632_), .A3(new_n637_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n595_), .A2(new_n620_), .A3(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n545_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n202_), .B1(new_n644_), .B2(new_n388_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT98), .Z(new_n646_));
  AND3_X1   g445(.A1(new_n323_), .A2(new_n335_), .A3(new_n389_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n453_), .A2(new_n460_), .A3(new_n459_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n459_), .B1(new_n453_), .B2(new_n460_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n647_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n468_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n314_), .A2(new_n319_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n209_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n470_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n651_), .A2(new_n653_), .A3(new_n324_), .A4(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n476_), .A2(new_n475_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n444_), .A2(new_n451_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(new_n658_), .A3(new_n415_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n650_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n540_), .A2(KEYINPUT37), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT37), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n662_), .B1(new_n536_), .B2(new_n539_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n643_), .A2(new_n660_), .A3(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(new_n202_), .A3(new_n388_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT38), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n646_), .A2(new_n668_), .ZN(G1324gat));
  NAND2_X1  g468(.A1(new_n323_), .A2(new_n335_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n666_), .A2(new_n603_), .A3(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n544_), .A2(KEYINPUT97), .ZN(new_n672_));
  INV_X1    g471(.A(new_n543_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n660_), .A2(KEYINPUT97), .A3(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n643_), .B(new_n670_), .C1(new_n672_), .C2(new_n674_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n675_), .A2(KEYINPUT99), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT39), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n603_), .B1(new_n675_), .B2(KEYINPUT99), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n676_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n677_), .B1(new_n676_), .B2(new_n678_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n671_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT101), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n671_), .B(new_n683_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1325gat));
  INV_X1    g486(.A(KEYINPUT41), .ZN(new_n688_));
  INV_X1    g487(.A(new_n658_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n644_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n691_), .A3(G15gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n691_), .B1(new_n690_), .B2(G15gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n688_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n694_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(KEYINPUT41), .A3(new_n692_), .ZN(new_n697_));
  INV_X1    g496(.A(G15gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n666_), .A2(new_n698_), .A3(new_n689_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n695_), .A2(new_n697_), .A3(new_n699_), .ZN(G1326gat));
  INV_X1    g499(.A(G22gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n459_), .B(KEYINPUT103), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n644_), .B2(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT42), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n666_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1327gat));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n707_), .B(new_n664_), .C1(new_n462_), .C2(new_n479_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n660_), .A2(KEYINPUT104), .A3(new_n707_), .A4(new_n664_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n664_), .B1(new_n462_), .B2(new_n479_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT43), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n710_), .A2(new_n711_), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n620_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n595_), .A2(new_n715_), .A3(new_n642_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n714_), .A2(KEYINPUT44), .A3(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(G29gat), .A3(new_n388_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT44), .B1(new_n714_), .B2(new_n716_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n540_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n480_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n716_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n722_), .A2(new_n389_), .ZN(new_n723_));
  OAI22_X1  g522(.A1(new_n718_), .A2(new_n719_), .B1(G29gat), .B2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT105), .Z(G1328gat));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n717_), .A2(new_n670_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G36gat), .B1(new_n727_), .B2(new_n719_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n729_));
  INV_X1    g528(.A(new_n670_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n730_), .A2(G36gat), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n722_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n728_), .A2(new_n729_), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n729_), .B1(new_n728_), .B2(new_n734_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n726_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n728_), .A2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT106), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n728_), .A2(new_n729_), .A3(new_n734_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(KEYINPUT46), .A3(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n737_), .A2(new_n741_), .ZN(G1329gat));
  XNOR2_X1  g541(.A(KEYINPUT107), .B(G43gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n743_), .B1(new_n722_), .B2(new_n658_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n717_), .A2(G43gat), .A3(new_n689_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(new_n719_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g546(.A(new_n722_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G50gat), .B1(new_n748_), .B2(new_n702_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n717_), .A2(G50gat), .A3(new_n459_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n719_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(G1331gat));
  NAND2_X1  g551(.A1(new_n642_), .A2(new_n715_), .ZN(new_n753_));
  NOR4_X1   g552(.A1(new_n480_), .A2(new_n594_), .A3(new_n664_), .A4(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT108), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n381_), .A3(new_n388_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n594_), .A2(new_n753_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n545_), .A2(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(new_n388_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n759_), .B2(new_n381_), .ZN(G1332gat));
  AOI21_X1  g559(.A(new_n549_), .B1(new_n758_), .B2(new_n670_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT48), .Z(new_n762_));
  NAND3_X1  g561(.A1(new_n755_), .A2(new_n549_), .A3(new_n670_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1333gat));
  INV_X1    g563(.A(G71gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n758_), .B2(new_n689_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT49), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n755_), .A2(new_n765_), .A3(new_n689_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1334gat));
  INV_X1    g568(.A(G78gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n758_), .B2(new_n702_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT50), .Z(new_n772_));
  NAND3_X1  g571(.A1(new_n755_), .A2(new_n770_), .A3(new_n702_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1335gat));
  NOR3_X1   g573(.A1(new_n594_), .A2(new_n715_), .A3(new_n641_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n714_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n389_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n721_), .A2(new_n775_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n388_), .A2(new_n383_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n777_), .B1(new_n778_), .B2(new_n779_), .ZN(G1336gat));
  INV_X1    g579(.A(G92gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n778_), .B2(new_n730_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT109), .Z(new_n783_));
  NOR3_X1   g582(.A1(new_n776_), .A2(new_n781_), .A3(new_n730_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1337gat));
  NAND4_X1  g584(.A1(new_n721_), .A2(new_n502_), .A3(new_n689_), .A4(new_n775_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT110), .Z(new_n787_));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n788_));
  OAI21_X1  g587(.A(G99gat), .B1(new_n776_), .B2(new_n658_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n787_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g590(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n776_), .B2(new_n415_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n714_), .A2(KEYINPUT112), .A3(new_n459_), .A4(new_n775_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(G106gat), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT52), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n794_), .A2(new_n798_), .A3(G106gat), .A4(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n778_), .A2(G106gat), .A3(new_n415_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n792_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n792_), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n804_), .B(new_n801_), .C1(new_n797_), .C2(new_n799_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1339gat));
  INV_X1    g605(.A(G113gat), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n670_), .A2(new_n389_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n649_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n641_), .A2(new_n588_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n576_), .A2(new_n571_), .A3(new_n579_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(G230gat), .A3(G233gat), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n580_), .A2(new_n815_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n570_), .A2(new_n508_), .B1(new_n524_), .B2(new_n578_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n817_), .A2(KEYINPUT55), .A3(new_n577_), .A4(new_n576_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n814_), .A2(new_n816_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n585_), .B1(new_n819_), .B2(KEYINPUT115), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n814_), .A2(new_n816_), .A3(new_n821_), .A4(new_n818_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n820_), .A2(KEYINPUT56), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT56), .B1(new_n820_), .B2(new_n822_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n812_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n622_), .A2(new_n630_), .A3(new_n625_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n629_), .A2(new_n623_), .A3(new_n631_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n638_), .A3(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n828_), .A2(new_n640_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n589_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n540_), .B1(new_n825_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n810_), .B1(new_n831_), .B2(KEYINPUT57), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n819_), .A2(KEYINPUT115), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n586_), .A3(new_n822_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n820_), .A2(KEYINPUT56), .A3(new_n822_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n811_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n830_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT116), .B(new_n833_), .C1(new_n841_), .C2(new_n540_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n832_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n837_), .A2(new_n844_), .A3(new_n838_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n829_), .A2(new_n588_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n824_), .B2(KEYINPUT117), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT118), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n665_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n845_), .A2(new_n847_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT58), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n850_), .A2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(KEYINPUT57), .B(new_n720_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n825_), .A2(new_n830_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n859_), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n720_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n843_), .A2(new_n855_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n620_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n595_), .A2(new_n664_), .A3(new_n753_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n866_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n865_), .A2(new_n864_), .A3(new_n866_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n809_), .B1(new_n863_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n807_), .B1(new_n874_), .B2(new_n642_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT120), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n877_), .B(new_n807_), .C1(new_n874_), .C2(new_n642_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n871_), .B1(new_n620_), .B2(new_n862_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT59), .B1(new_n879_), .B2(new_n809_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n809_), .A2(KEYINPUT59), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n831_), .A2(KEYINPUT57), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n850_), .B2(new_n854_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n715_), .B1(new_n883_), .B2(new_n861_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n881_), .B1(new_n884_), .B2(new_n871_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n880_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n642_), .A2(new_n807_), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n876_), .A2(new_n878_), .B1(new_n887_), .B2(new_n888_), .ZN(G1340gat));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n595_), .B(new_n885_), .C1(new_n873_), .C2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n880_), .A2(KEYINPUT122), .A3(new_n595_), .A4(new_n885_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(G120gat), .A3(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(G120gat), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(KEYINPUT60), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n594_), .B2(KEYINPUT60), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(KEYINPUT121), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n873_), .B(new_n899_), .C1(KEYINPUT121), .C2(new_n898_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n895_), .A2(new_n900_), .ZN(G1341gat));
  OAI21_X1  g700(.A(G127gat), .B1(new_n886_), .B2(new_n620_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n620_), .A2(G127gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n874_), .B2(new_n903_), .ZN(G1342gat));
  OAI21_X1  g703(.A(G134gat), .B1(new_n886_), .B2(new_n665_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n673_), .A2(G134gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n874_), .B2(new_n906_), .ZN(G1343gat));
  NOR2_X1   g706(.A1(new_n879_), .A2(new_n461_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n908_), .A2(new_n641_), .A3(new_n808_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g709(.A1(new_n908_), .A2(new_n595_), .A3(new_n808_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g711(.A1(new_n908_), .A2(new_n715_), .A3(new_n808_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT61), .B(G155gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1346gat));
  NAND2_X1  g714(.A1(new_n908_), .A2(new_n808_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G162gat), .B1(new_n916_), .B2(new_n665_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n673_), .A2(G162gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n916_), .B2(new_n918_), .ZN(G1347gat));
  OR2_X1    g718(.A1(new_n884_), .A2(new_n871_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n730_), .A2(new_n388_), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n921_), .A2(KEYINPUT123), .A3(new_n689_), .ZN(new_n922_));
  AOI21_X1  g721(.A(KEYINPUT123), .B1(new_n921_), .B2(new_n689_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n702_), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n920_), .A2(new_n925_), .A3(KEYINPUT124), .A4(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n884_), .A2(new_n871_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n926_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n928_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n270_), .A2(new_n283_), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n927_), .A2(new_n931_), .A3(new_n641_), .A4(new_n932_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n920_), .A2(new_n925_), .A3(new_n641_), .A4(new_n926_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n934_), .A2(new_n935_), .A3(G169gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n934_), .B2(G169gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n933_), .B1(new_n936_), .B2(new_n937_), .ZN(G1348gat));
  NAND3_X1  g737(.A1(new_n927_), .A2(new_n595_), .A3(new_n931_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n879_), .A2(new_n459_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n924_), .A2(new_n256_), .A3(new_n594_), .ZN(new_n941_));
  AOI22_X1  g740(.A1(new_n939_), .A2(new_n256_), .B1(new_n940_), .B2(new_n941_), .ZN(G1349gat));
  NAND4_X1  g741(.A1(new_n927_), .A2(new_n931_), .A3(new_n715_), .A4(new_n289_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n940_), .A2(new_n715_), .A3(new_n925_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n231_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n943_), .A2(new_n945_), .ZN(G1350gat));
  NAND4_X1  g745(.A1(new_n927_), .A2(new_n931_), .A3(new_n543_), .A4(new_n240_), .ZN(new_n947_));
  AND3_X1   g746(.A1(new_n927_), .A2(new_n664_), .A3(new_n931_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n948_), .B2(new_n236_), .ZN(G1351gat));
  NAND2_X1  g748(.A1(new_n863_), .A2(new_n872_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n950_), .A2(new_n648_), .A3(new_n921_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n951_), .A2(new_n642_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(new_n212_), .ZN(G1352gat));
  NOR2_X1   g752(.A1(new_n951_), .A2(new_n594_), .ZN(new_n954_));
  OR2_X1    g753(.A1(new_n215_), .A2(KEYINPUT125), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n954_), .B(new_n955_), .ZN(G1353gat));
  AOI21_X1  g755(.A(new_n620_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n957_));
  XOR2_X1   g756(.A(new_n957_), .B(KEYINPUT126), .Z(new_n958_));
  NOR2_X1   g757(.A1(new_n951_), .A2(new_n958_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n959_), .B(new_n960_), .ZN(G1354gat));
  NAND4_X1  g760(.A1(new_n950_), .A2(new_n543_), .A3(new_n648_), .A4(new_n921_), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n963_));
  OR2_X1    g762(.A1(new_n962_), .A2(new_n963_), .ZN(new_n964_));
  AOI21_X1  g763(.A(G218gat), .B1(new_n962_), .B2(new_n963_), .ZN(new_n965_));
  INV_X1    g764(.A(new_n951_), .ZN(new_n966_));
  AND2_X1   g765(.A1(new_n664_), .A2(G218gat), .ZN(new_n967_));
  AOI22_X1  g766(.A1(new_n964_), .A2(new_n965_), .B1(new_n966_), .B2(new_n967_), .ZN(G1355gat));
endmodule


