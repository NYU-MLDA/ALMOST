//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_, new_n958_, new_n959_,
    new_n960_, new_n962_, new_n963_, new_n965_, new_n967_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_, new_n978_;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT81), .B(KEYINPUT37), .Z(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT78), .ZN(new_n205_));
  XOR2_X1   g004(.A(G85gat), .B(G92gat), .Z(new_n206_));
  INV_X1    g005(.A(KEYINPUT8), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NOR3_X1   g009(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT6), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n208_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT67), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT6), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n219_), .A3(new_n213_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n211_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(new_n209_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n213_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n206_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n207_), .B1(new_n224_), .B2(KEYINPUT68), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n226_), .B(new_n206_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n215_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n214_), .ZN(new_n229_));
  XOR2_X1   g028(.A(KEYINPUT10), .B(G99gat), .Z(new_n230_));
  INV_X1    g029(.A(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n229_), .B1(new_n232_), .B2(KEYINPUT65), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n232_), .A2(KEYINPUT65), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT66), .B(G85gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G92gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n233_), .A2(new_n234_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT69), .B1(new_n228_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n244_));
  INV_X1    g043(.A(new_n227_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n213_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n218_), .A2(KEYINPUT6), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n216_), .A2(KEYINPUT67), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(new_n212_), .A3(new_n220_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n226_), .B1(new_n250_), .B2(new_n206_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n245_), .A2(new_n251_), .A3(new_n207_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n244_), .B(new_n241_), .C1(new_n252_), .C2(new_n215_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT15), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G29gat), .B(G36gat), .ZN(new_n255_));
  INV_X1    g054(.A(G43gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G29gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(G36gat), .ZN(new_n259_));
  INV_X1    g058(.A(G36gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(G29gat), .ZN(new_n261_));
  NOR3_X1   g060(.A1(new_n259_), .A2(new_n261_), .A3(G43gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT76), .B1(new_n257_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n255_), .A2(new_n256_), .ZN(new_n264_));
  OAI21_X1  g063(.A(G43gat), .B1(new_n259_), .B2(new_n261_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT76), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(G50gat), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(G50gat), .B1(new_n263_), .B2(new_n267_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n254_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n263_), .A2(new_n267_), .ZN(new_n272_));
  INV_X1    g071(.A(G50gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n274_), .A2(KEYINPUT15), .A3(new_n268_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n243_), .A2(new_n253_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G232gat), .A2(G233gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n278_), .B(KEYINPUT74), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT34), .ZN(new_n280_));
  XOR2_X1   g079(.A(KEYINPUT75), .B(KEYINPUT35), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n280_), .A2(new_n282_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n228_), .A2(new_n242_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n269_), .A2(new_n270_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n284_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n277_), .A2(new_n283_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n283_), .B1(new_n277_), .B2(new_n287_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G190gat), .B(G218gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(G134gat), .B(G162gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT36), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n295_), .B(KEYINPUT77), .Z(new_n296_));
  AOI21_X1  g095(.A(new_n205_), .B1(new_n290_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n296_), .ZN(new_n298_));
  NOR4_X1   g097(.A1(new_n288_), .A2(new_n289_), .A3(KEYINPUT78), .A4(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n204_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT79), .B1(new_n288_), .B2(new_n289_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n277_), .A2(new_n287_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n283_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT79), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n277_), .A2(new_n287_), .A3(new_n283_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n293_), .B(KEYINPUT36), .ZN(new_n308_));
  AND4_X1   g107(.A1(KEYINPUT80), .A2(new_n301_), .A3(new_n307_), .A4(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n301_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n300_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n304_), .A2(new_n306_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n308_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n317_), .A2(KEYINPUT37), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT82), .B1(new_n314_), .B2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT78), .B1(new_n315_), .B2(new_n298_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n290_), .A2(new_n205_), .A3(new_n296_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n203_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n308_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n323_), .B1(new_n315_), .B2(KEYINPUT79), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT80), .B1(new_n324_), .B2(new_n307_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n322_), .B1(new_n325_), .B2(new_n309_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT82), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n317_), .A2(KEYINPUT37), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n319_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G127gat), .B(G155gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT16), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G183gat), .ZN(new_n333_));
  INV_X1    g132(.A(G211gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT17), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G57gat), .B(G64gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n339_), .A2(KEYINPUT11), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G71gat), .B(G78gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(KEYINPUT11), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n339_), .A2(new_n341_), .A3(KEYINPUT11), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT83), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G15gat), .B(G22gat), .ZN(new_n348_));
  INV_X1    g147(.A(G1gat), .ZN(new_n349_));
  INV_X1    g148(.A(G8gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT14), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G1gat), .B(G8gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G231gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n347_), .B(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n335_), .A2(new_n336_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n338_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n346_), .B(KEYINPUT70), .ZN(new_n360_));
  INV_X1    g159(.A(new_n356_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n361_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n337_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n359_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT84), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n330_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n241_), .B1(new_n252_), .B2(new_n215_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n346_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT12), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n369_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G230gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT64), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT12), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n360_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(new_n243_), .A3(new_n253_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n372_), .A2(new_n375_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n371_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n368_), .A2(new_n369_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n374_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n384_));
  XNOR2_X1  g183(.A(G120gat), .B(G148gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G176gat), .B(G204gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n388_), .B(KEYINPUT72), .Z(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n383_), .B2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n392_));
  OR2_X1    g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n202_), .B1(new_n367_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n393_), .A2(new_n395_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n330_), .A2(KEYINPUT85), .A3(new_n398_), .A4(new_n366_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT23), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n400_), .B1(G183gat), .B2(G190gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G183gat), .A2(G190gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT88), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT88), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(G183gat), .A3(G190gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n401_), .B1(new_n406_), .B2(new_n400_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT25), .B(G183gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT26), .B(G190gat), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n407_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G169gat), .A2(G176gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT24), .A4(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(KEYINPUT24), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT87), .B1(new_n418_), .B2(new_n413_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n402_), .A2(new_n400_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(new_n406_), .B2(KEYINPUT23), .ZN(new_n423_));
  NOR2_X1   g222(.A1(G183gat), .A2(G190gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT22), .B(G169gat), .ZN(new_n427_));
  INV_X1    g226(.A(G176gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n416_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n412_), .A2(new_n420_), .B1(new_n426_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT30), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G227gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n433_), .B(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT31), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n433_), .B(new_n434_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT31), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G71gat), .B(G99gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(G15gat), .B(G43gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT89), .B(KEYINPUT90), .Z(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(G127gat), .B(G134gat), .Z(new_n446_));
  XOR2_X1   g245(.A(G113gat), .B(G120gat), .Z(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n445_), .B(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n437_), .A2(new_n440_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n426_), .A2(new_n431_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n407_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n411_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n420_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G211gat), .B(G218gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G204gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G197gat), .ZN(new_n463_));
  INV_X1    g262(.A(G197gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(G204gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(KEYINPUT21), .A3(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT96), .B1(new_n464_), .B2(G204gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT96), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(new_n462_), .A3(G197gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n470_), .A3(new_n465_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n471_), .A2(KEYINPUT21), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n460_), .B1(new_n466_), .B2(KEYINPUT21), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n467_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n454_), .B1(new_n459_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n406_), .A2(KEYINPUT23), .ZN(new_n476_));
  INV_X1    g275(.A(new_n411_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n421_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT101), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n423_), .A2(KEYINPUT101), .A3(new_n477_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT26), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(G190gat), .ZN(new_n483_));
  INV_X1    g282(.A(G190gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n484_), .A2(KEYINPUT26), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT99), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(KEYINPUT26), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n482_), .A2(G190gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT99), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(new_n408_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT100), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n418_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n416_), .A2(KEYINPUT100), .A3(KEYINPUT24), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n414_), .A3(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n480_), .A2(new_n481_), .A3(new_n491_), .A4(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n474_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n430_), .B1(new_n456_), .B2(new_n425_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n475_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G226gat), .A2(G233gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT19), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT101), .B1(new_n423_), .B2(new_n477_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n491_), .A2(new_n495_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n498_), .B1(new_n507_), .B2(new_n481_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT102), .B1(new_n508_), .B2(new_n497_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT102), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n400_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n511_));
  NOR4_X1   g310(.A1(new_n511_), .A2(new_n422_), .A3(new_n479_), .A4(new_n411_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n505_), .A2(new_n506_), .A3(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n510_), .B(new_n474_), .C1(new_n513_), .C2(new_n498_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n454_), .B1(new_n432_), .B2(new_n497_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n509_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n504_), .B1(new_n516_), .B2(new_n503_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G8gat), .B(G36gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT18), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(G64gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(G92gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n522_), .A2(KEYINPUT32), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n517_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n497_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n515_), .B1(new_n525_), .B2(new_n510_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n514_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n503_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n503_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n475_), .A2(new_n500_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n446_), .B(new_n447_), .Z(new_n533_));
  NAND2_X1  g332(.A1(G141gat), .A2(G148gat), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT92), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT2), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT2), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n534_), .A2(new_n535_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n540_));
  OAI22_X1  g339(.A1(new_n540_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n541_));
  NOR2_X1   g340(.A1(G141gat), .A2(G148gat), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT3), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(KEYINPUT91), .A3(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n537_), .A2(new_n539_), .A3(new_n541_), .A4(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(G155gat), .A2(G162gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G155gat), .A2(G162gat), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n542_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n550_), .A2(new_n534_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT1), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n546_), .A2(new_n553_), .A3(new_n547_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n549_), .A2(new_n555_), .ZN(new_n556_));
  OR3_X1    g355(.A1(new_n533_), .A2(new_n556_), .A3(KEYINPUT103), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n533_), .A2(new_n556_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n545_), .A2(new_n548_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n448_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(KEYINPUT103), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G225gat), .A2(G233gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n557_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n557_), .A2(new_n561_), .A3(KEYINPUT4), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT4), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n558_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n563_), .B1(new_n567_), .B2(new_n562_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G57gat), .B(G85gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(G1gat), .B(G29gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(KEYINPUT104), .B(KEYINPUT0), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n568_), .A2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n568_), .A2(new_n574_), .ZN(new_n576_));
  OAI221_X1 g375(.A(new_n524_), .B1(new_n523_), .B2(new_n532_), .C1(new_n575_), .C2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n568_), .A2(new_n574_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT105), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT106), .B1(new_n557_), .B2(new_n561_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(new_n562_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n557_), .A2(new_n561_), .A3(KEYINPUT106), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n567_), .A2(new_n562_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n573_), .A3(new_n586_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n568_), .B(new_n574_), .C1(KEYINPUT105), .C2(KEYINPUT33), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n581_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT20), .B1(new_n459_), .B2(new_n474_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n474_), .B1(new_n513_), .B2(new_n498_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n591_), .B2(KEYINPUT102), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n529_), .B1(new_n592_), .B2(new_n514_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n521_), .B1(new_n593_), .B2(new_n530_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n528_), .A2(new_n522_), .A3(new_n531_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n577_), .B1(new_n589_), .B2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G22gat), .B(G50gat), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT29), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n549_), .A2(new_n600_), .A3(new_n555_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT28), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT93), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT28), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n559_), .A2(new_n604_), .A3(new_n600_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n602_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n603_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n599_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  AND4_X1   g407(.A1(new_n604_), .A2(new_n549_), .A3(new_n600_), .A4(new_n555_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n604_), .B1(new_n559_), .B2(new_n600_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT93), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n602_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n598_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT94), .B(G228gat), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT95), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n474_), .B(new_n616_), .C1(new_n600_), .C2(new_n559_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT97), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n615_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n559_), .A2(new_n600_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n620_), .B1(new_n621_), .B2(new_n497_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n556_), .A2(KEYINPUT29), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n623_), .A2(KEYINPUT97), .A3(new_n474_), .A4(new_n616_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n619_), .A2(new_n622_), .A3(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n608_), .A2(new_n613_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G78gat), .B(G106gat), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n608_), .A2(new_n613_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n625_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n630_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  AOI211_X1 g432(.A(new_n629_), .B(new_n625_), .C1(new_n608_), .C2(new_n613_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n628_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n611_), .A2(new_n598_), .A3(new_n612_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n598_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n632_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n629_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n631_), .A2(new_n632_), .A3(new_n630_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n639_), .A2(new_n627_), .A3(new_n640_), .A4(new_n626_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n635_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n597_), .A2(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n635_), .A2(new_n641_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n575_), .A2(new_n576_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT27), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n530_), .B1(new_n516_), .B2(new_n503_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n647_), .B2(new_n522_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n517_), .A2(new_n521_), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n596_), .A2(new_n646_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n644_), .A2(new_n645_), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n453_), .B1(new_n643_), .B2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n645_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n650_), .A2(KEYINPUT107), .A3(new_n642_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT107), .B1(new_n650_), .B2(new_n642_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n654_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT108), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n659_));
  AOI211_X1 g458(.A(new_n521_), .B(new_n530_), .C1(new_n516_), .C2(new_n503_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n522_), .B1(new_n528_), .B2(new_n531_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n646_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n649_), .A2(KEYINPUT27), .A3(new_n595_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n659_), .B1(new_n644_), .B2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n650_), .A2(KEYINPUT107), .A3(new_n642_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n654_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n652_), .B1(new_n658_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n276_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(new_n354_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(G229gat), .A2(G233gat), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n286_), .B2(new_n354_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n286_), .B(new_n354_), .ZN(new_n677_));
  AOI22_X1  g476(.A1(new_n673_), .A2(new_n676_), .B1(new_n677_), .B2(new_n675_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(G169gat), .B(G197gat), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT86), .ZN(new_n680_));
  XNOR2_X1  g479(.A(G113gat), .B(G141gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n678_), .B(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n670_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n397_), .A2(new_n399_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n397_), .A2(KEYINPUT109), .A3(new_n399_), .A4(new_n685_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n645_), .A2(G1gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT110), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n688_), .A2(new_n693_), .A3(new_n689_), .A4(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT38), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n643_), .A2(new_n651_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n452_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n668_), .B1(new_n667_), .B2(new_n654_), .ZN(new_n700_));
  AOI211_X1 g499(.A(KEYINPUT108), .B(new_n653_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n699_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n320_), .A2(new_n321_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n325_), .B2(new_n309_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(KEYINPUT112), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(KEYINPUT112), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n645_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n398_), .A2(new_n683_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n711_), .A2(new_n365_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT111), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n710_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G1gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n692_), .A2(KEYINPUT38), .A3(new_n694_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n697_), .A2(new_n715_), .A3(new_n716_), .ZN(G1324gat));
  NAND4_X1  g516(.A1(new_n688_), .A2(new_n350_), .A3(new_n664_), .A4(new_n689_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n713_), .B(new_n664_), .C1(new_n707_), .C2(new_n706_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT39), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(new_n720_), .A3(G8gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n719_), .B2(G8gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT40), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OAI211_X1 g524(.A(KEYINPUT40), .B(new_n718_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1325gat));
  NOR2_X1   g526(.A1(new_n452_), .A2(G15gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n688_), .A2(new_n689_), .A3(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n709_), .A2(new_n453_), .A3(new_n713_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n730_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT41), .B1(new_n730_), .B2(G15gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n729_), .B1(new_n731_), .B2(new_n732_), .ZN(G1326gat));
  NOR2_X1   g532(.A1(new_n642_), .A2(G22gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n688_), .A2(new_n689_), .A3(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n709_), .A2(new_n644_), .A3(new_n713_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G22gat), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n737_), .A2(KEYINPUT42), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(KEYINPUT42), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(G1327gat));
  INV_X1    g539(.A(new_n366_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n398_), .A2(new_n741_), .A3(new_n683_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n670_), .A2(new_n330_), .A3(KEYINPUT43), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n327_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n745_), .B1(new_n702_), .B2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n743_), .B1(new_n744_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(KEYINPUT43), .B1(new_n670_), .B2(new_n330_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n702_), .A2(new_n748_), .A3(new_n745_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(KEYINPUT44), .A3(new_n743_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n752_), .A2(new_n710_), .A3(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n258_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n759_), .B1(new_n758_), .B2(new_n757_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n670_), .A2(new_n704_), .A3(new_n742_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n258_), .A3(new_n710_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1328gat));
  NOR2_X1   g562(.A1(new_n650_), .A2(G36gat), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n761_), .A2(KEYINPUT45), .A3(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT44), .B1(new_n755_), .B2(new_n743_), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n751_), .B(new_n742_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n650_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n770_), .B1(new_n773_), .B2(new_n260_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT46), .B1(new_n774_), .B2(KEYINPUT114), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n752_), .A2(new_n664_), .A3(new_n756_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n769_), .B1(new_n776_), .B2(G36gat), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n775_), .A2(new_n780_), .ZN(G1329gat));
  NAND4_X1  g580(.A1(new_n752_), .A2(G43gat), .A3(new_n453_), .A4(new_n756_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n761_), .A2(new_n453_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(G43gat), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g584(.A1(new_n642_), .A2(G50gat), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT115), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n761_), .A2(new_n787_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n771_), .A2(new_n772_), .A3(new_n642_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(new_n273_), .ZN(G1331gat));
  NOR2_X1   g589(.A1(new_n398_), .A2(new_n683_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n708_), .A2(new_n741_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(G57gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT117), .B1(new_n645_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n367_), .A2(new_n792_), .A3(new_n670_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n645_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n796_), .B(new_n799_), .C1(new_n798_), .C2(new_n797_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n796_), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n800_), .A2(new_n794_), .B1(KEYINPUT117), .B2(new_n801_), .ZN(G1332gat));
  INV_X1    g601(.A(G64gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n797_), .A2(new_n803_), .A3(new_n664_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT48), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n793_), .A2(new_n664_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(G64gat), .ZN(new_n807_));
  AOI211_X1 g606(.A(KEYINPUT48), .B(new_n803_), .C1(new_n793_), .C2(new_n664_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(G1333gat));
  INV_X1    g608(.A(G71gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n797_), .A2(new_n810_), .A3(new_n453_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n793_), .B2(new_n453_), .ZN(new_n812_));
  XOR2_X1   g611(.A(KEYINPUT118), .B(KEYINPUT49), .Z(new_n813_));
  AND2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n812_), .A2(new_n813_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n811_), .B1(new_n814_), .B2(new_n815_), .ZN(G1334gat));
  INV_X1    g615(.A(G78gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n797_), .A2(new_n817_), .A3(new_n644_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n793_), .A2(new_n644_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(G78gat), .ZN(new_n821_));
  AOI211_X1 g620(.A(KEYINPUT50), .B(new_n817_), .C1(new_n793_), .C2(new_n644_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n818_), .B1(new_n821_), .B2(new_n822_), .ZN(G1335gat));
  NAND2_X1  g622(.A1(new_n791_), .A2(new_n741_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n824_), .A2(new_n670_), .A3(new_n704_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT119), .ZN(new_n826_));
  AOI21_X1  g625(.A(G85gat), .B1(new_n826_), .B2(new_n710_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n824_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n710_), .A2(new_n235_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n827_), .B1(new_n828_), .B2(new_n829_), .ZN(G1336gat));
  AOI21_X1  g629(.A(G92gat), .B1(new_n826_), .B2(new_n664_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n664_), .A2(G92gat), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n832_), .B(KEYINPUT120), .Z(new_n833_));
  AOI21_X1  g632(.A(new_n831_), .B1(new_n828_), .B2(new_n833_), .ZN(G1337gat));
  NAND3_X1  g633(.A1(new_n826_), .A2(new_n230_), .A3(new_n453_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n828_), .A2(new_n453_), .ZN(new_n836_));
  INV_X1    g635(.A(G99gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n835_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g638(.A1(new_n826_), .A2(new_n231_), .A3(new_n644_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n828_), .A2(new_n644_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(G106gat), .ZN(new_n843_));
  AOI211_X1 g642(.A(KEYINPUT52), .B(new_n231_), .C1(new_n828_), .C2(new_n644_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n840_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g645(.A1(new_n667_), .A2(new_n453_), .A3(new_n710_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(KEYINPUT59), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n678_), .A2(new_n682_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n682_), .B1(new_n677_), .B2(new_n674_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n286_), .A2(new_n354_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n675_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n672_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n391_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n372_), .A2(KEYINPUT55), .A3(new_n378_), .A4(new_n375_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n856_), .A2(KEYINPUT122), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(KEYINPUT122), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n372_), .A2(new_n378_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n374_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n379_), .A2(new_n861_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n857_), .A2(new_n858_), .A3(new_n860_), .A4(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n390_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n858_), .A2(new_n860_), .A3(new_n862_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n856_), .A2(KEYINPUT122), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT56), .B(new_n390_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT123), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n863_), .A2(new_n871_), .A3(KEYINPUT56), .A4(new_n390_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n866_), .A2(new_n870_), .A3(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n684_), .A2(new_n389_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n855_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n704_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(new_n879_));
  AOI211_X1 g678(.A(new_n389_), .B(new_n854_), .C1(new_n866_), .C2(new_n869_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n880_), .A2(KEYINPUT58), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(KEYINPUT58), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n748_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n366_), .B1(new_n879_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n396_), .A2(new_n683_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(new_n330_), .A3(new_n366_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n885_), .B1(new_n887_), .B2(KEYINPUT54), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n748_), .A2(new_n741_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n889_), .A2(KEYINPUT121), .A3(new_n890_), .A4(new_n886_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n887_), .A2(KEYINPUT54), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n888_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n848_), .B1(new_n884_), .B2(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n877_), .A2(new_n878_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n875_), .A2(new_n876_), .A3(KEYINPUT57), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n883_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n365_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n888_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n847_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n894_), .B(new_n683_), .C1(new_n900_), .C2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G113gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n898_), .A2(new_n899_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n847_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  OR3_X1    g705(.A1(new_n906_), .A2(G113gat), .A3(new_n684_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n907_), .ZN(G1340gat));
  OAI211_X1 g707(.A(new_n894_), .B(new_n396_), .C1(new_n900_), .C2(new_n901_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(G120gat), .ZN(new_n910_));
  INV_X1    g709(.A(G120gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n911_), .B1(new_n398_), .B2(KEYINPUT60), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n900_), .B(new_n912_), .C1(KEYINPUT60), .C2(new_n911_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n913_), .ZN(G1341gat));
  INV_X1    g713(.A(new_n365_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n894_), .B(new_n915_), .C1(new_n900_), .C2(new_n901_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G127gat), .ZN(new_n917_));
  OR3_X1    g716(.A1(new_n906_), .A2(G127gat), .A3(new_n741_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1342gat));
  OAI211_X1 g718(.A(new_n894_), .B(new_n748_), .C1(new_n900_), .C2(new_n901_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(G134gat), .ZN(new_n921_));
  OR3_X1    g720(.A1(new_n906_), .A2(G134gat), .A3(new_n704_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1343gat));
  NOR2_X1   g722(.A1(new_n453_), .A2(new_n642_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n664_), .A2(new_n645_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n904_), .A2(new_n683_), .A3(new_n924_), .A4(new_n925_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(KEYINPUT124), .B(G141gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1344gat));
  NAND4_X1  g727(.A1(new_n904_), .A2(new_n396_), .A3(new_n924_), .A4(new_n925_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g729(.A1(new_n904_), .A2(new_n366_), .A3(new_n924_), .A4(new_n925_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT61), .B(G155gat), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n931_), .B(new_n932_), .ZN(G1346gat));
  NAND3_X1  g732(.A1(new_n904_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n934_));
  OAI21_X1  g733(.A(G162gat), .B1(new_n934_), .B2(new_n330_), .ZN(new_n935_));
  OR2_X1    g734(.A1(new_n704_), .A2(G162gat), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n934_), .B2(new_n936_), .ZN(G1347gat));
  NOR2_X1   g736(.A1(new_n650_), .A2(new_n710_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n939_), .A2(new_n452_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n644_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n897_), .A2(new_n741_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n943_), .B1(new_n944_), .B2(new_n899_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  OAI211_X1 g745(.A(KEYINPUT62), .B(G169gat), .C1(new_n946_), .C2(new_n684_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n948_));
  AOI211_X1 g747(.A(new_n684_), .B(new_n943_), .C1(new_n944_), .C2(new_n899_), .ZN(new_n949_));
  INV_X1    g748(.A(G169gat), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n948_), .B1(new_n949_), .B2(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n949_), .A2(new_n427_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n947_), .A2(new_n951_), .A3(new_n952_), .ZN(G1348gat));
  AOI21_X1  g752(.A(G176gat), .B1(new_n945_), .B2(new_n396_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n644_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n941_), .A2(new_n398_), .A3(new_n428_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n954_), .B1(new_n955_), .B2(new_n956_), .ZN(G1349gat));
  NAND3_X1  g756(.A1(new_n955_), .A2(new_n366_), .A3(new_n940_), .ZN(new_n958_));
  INV_X1    g757(.A(G183gat), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n365_), .A2(new_n408_), .ZN(new_n960_));
  AOI22_X1  g759(.A1(new_n958_), .A2(new_n959_), .B1(new_n945_), .B2(new_n960_), .ZN(G1350gat));
  OAI21_X1  g760(.A(G190gat), .B1(new_n946_), .B2(new_n330_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n876_), .A2(new_n486_), .A3(new_n490_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n962_), .B1(new_n946_), .B2(new_n963_), .ZN(G1351gat));
  NAND4_X1  g763(.A1(new_n904_), .A2(new_n683_), .A3(new_n924_), .A4(new_n938_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g765(.A1(new_n904_), .A2(new_n396_), .A3(new_n924_), .A4(new_n938_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n462_), .A2(KEYINPUT125), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n967_), .B(new_n968_), .ZN(G1353gat));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n915_), .B1(new_n970_), .B2(new_n334_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(KEYINPUT126), .ZN(new_n972_));
  NAND4_X1  g771(.A1(new_n904_), .A2(new_n924_), .A3(new_n938_), .A4(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n970_), .A2(new_n334_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n973_), .B(new_n974_), .ZN(G1354gat));
  NAND3_X1  g774(.A1(new_n904_), .A2(new_n924_), .A3(new_n938_), .ZN(new_n976_));
  OAI21_X1  g775(.A(G218gat), .B1(new_n976_), .B2(new_n330_), .ZN(new_n977_));
  OR2_X1    g776(.A1(new_n704_), .A2(G218gat), .ZN(new_n978_));
  OAI21_X1  g777(.A(new_n977_), .B1(new_n976_), .B2(new_n978_), .ZN(G1355gat));
endmodule


