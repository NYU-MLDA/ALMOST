//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n208_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT26), .B(G190gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT25), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(G183gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n217_), .B(new_n220_), .C1(new_n221_), .C2(new_n218_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n216_), .A2(new_n222_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n213_), .B(new_n214_), .C1(G183gat), .C2(G190gat), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n204_), .A2(KEYINPUT78), .A3(KEYINPUT22), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT78), .B1(new_n204_), .B2(KEYINPUT22), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT79), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n204_), .B2(KEYINPUT22), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n205_), .A3(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n207_), .B(new_n224_), .C1(new_n227_), .C2(new_n232_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n223_), .A2(KEYINPUT30), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT30), .B1(new_n223_), .B2(new_n233_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n203_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n223_), .A2(new_n233_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT30), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n223_), .A2(KEYINPUT30), .A3(new_n233_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n202_), .A3(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G71gat), .B(G99gat), .ZN(new_n242_));
  INV_X1    g041(.A(G43gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n236_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n245_), .B1(new_n236_), .B2(new_n241_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT80), .B(G15gat), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT82), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n249_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n236_), .A2(new_n241_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n244_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n236_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n249_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT82), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n254_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(new_n251_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G127gat), .B(G134gat), .Z(new_n263_));
  XOR2_X1   g062(.A(G113gat), .B(G120gat), .Z(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n255_), .A2(new_n262_), .A3(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n266_), .B1(new_n255_), .B2(new_n262_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT85), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT84), .B(KEYINPUT2), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n270_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT2), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n275_), .A2(KEYINPUT84), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(KEYINPUT84), .ZN(new_n277_));
  OAI211_X1 g076(.A(KEYINPUT85), .B(new_n272_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G141gat), .A2(G148gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT3), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT3), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(G141gat), .B2(G148gat), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n280_), .A2(new_n282_), .B1(new_n273_), .B2(KEYINPUT2), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n274_), .A2(new_n278_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT83), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n290_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n287_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n285_), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n273_), .A2(new_n279_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n289_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n266_), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n284_), .A2(new_n288_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n265_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(KEYINPUT4), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G225gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT93), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n265_), .B1(new_n289_), .B2(new_n297_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT94), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT94), .ZN(new_n308_));
  NOR4_X1   g107(.A1(new_n300_), .A2(new_n308_), .A3(KEYINPUT4), .A4(new_n265_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n302_), .B(new_n304_), .C1(new_n307_), .C2(new_n309_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n299_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G1gat), .B(G29gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G57gat), .B(G85gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n310_), .A2(new_n312_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT98), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n310_), .A2(KEYINPUT98), .A3(new_n312_), .A4(new_n317_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n310_), .A2(new_n312_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n317_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G228gat), .A2(G233gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n327_), .B(KEYINPUT86), .Z(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(new_n289_), .B2(new_n297_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G197gat), .A2(G204gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G197gat), .A2(G204gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(KEYINPUT21), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT21), .ZN(new_n336_));
  INV_X1    g135(.A(new_n334_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(new_n332_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G211gat), .B(G218gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n340_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n335_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n329_), .B1(new_n331_), .B2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n342_), .B1(new_n335_), .B2(new_n338_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n342_), .A2(new_n335_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n348_), .B(new_n328_), .C1(new_n300_), .C2(new_n330_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G78gat), .B(G106gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n351_), .B(KEYINPUT87), .Z(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT88), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT88), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(new_n355_), .A3(new_n352_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n350_), .A2(new_n352_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n300_), .A2(new_n361_), .A3(new_n330_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n361_), .B1(new_n300_), .B2(new_n330_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n360_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n364_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(new_n362_), .A3(new_n359_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n345_), .A2(new_n349_), .A3(new_n351_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT89), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n350_), .A2(new_n371_), .A3(new_n352_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n358_), .A2(new_n368_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT27), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT19), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n224_), .A2(new_n207_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n230_), .A2(G169gat), .ZN(new_n382_));
  AOI21_X1  g181(.A(G176gat), .B1(new_n382_), .B2(new_n228_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n383_), .B(new_n231_), .C1(new_n226_), .C2(new_n225_), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n381_), .A2(new_n384_), .B1(new_n216_), .B2(new_n222_), .ZN(new_n385_));
  OAI211_X1 g184(.A(KEYINPUT20), .B(new_n380_), .C1(new_n385_), .C2(new_n344_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n204_), .A2(KEYINPUT22), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(new_n382_), .A3(new_n205_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n224_), .A2(new_n388_), .A3(new_n207_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n217_), .A2(new_n221_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n213_), .A2(new_n214_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .A4(new_n210_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT90), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT90), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n216_), .A2(new_n396_), .A3(new_n391_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n390_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT91), .B1(new_n386_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n397_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n224_), .A2(new_n207_), .A3(new_n388_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n401_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT20), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n237_), .B2(new_n348_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT91), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n403_), .A2(new_n405_), .A3(new_n406_), .A4(new_n380_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n399_), .A2(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G8gat), .B(G36gat), .Z(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G64gat), .B(G92gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n385_), .A2(new_n344_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n401_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n414_), .B(KEYINPUT20), .C1(new_n415_), .C2(new_n344_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n379_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n408_), .A2(new_n413_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n413_), .B1(new_n408_), .B2(new_n417_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n377_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n394_), .B(new_n389_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n421_), .B(KEYINPUT20), .C1(new_n385_), .C2(new_n344_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n379_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(new_n416_), .B2(new_n379_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT99), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n413_), .B(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n377_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n408_), .A2(new_n413_), .A3(new_n417_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT100), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n429_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n420_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n376_), .A2(new_n432_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n269_), .A2(new_n326_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT101), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n413_), .A2(KEYINPUT32), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n424_), .A2(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n408_), .A2(new_n417_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(new_n439_), .B2(new_n436_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n304_), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n289_), .A2(new_n297_), .A3(new_n265_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(new_n305_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n441_), .B1(new_n443_), .B2(KEYINPUT4), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n298_), .A2(new_n306_), .A3(new_n266_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n308_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n305_), .A2(KEYINPUT94), .A3(new_n306_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n311_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n321_), .B1(new_n449_), .B2(new_n317_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT98), .B1(new_n449_), .B2(new_n317_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n440_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n318_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT96), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT96), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n318_), .A2(new_n456_), .A3(new_n453_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n299_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n323_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n302_), .B(new_n303_), .C1(new_n307_), .C2(new_n309_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n460_), .B1(new_n461_), .B2(KEYINPUT97), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT97), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n448_), .A2(new_n463_), .A3(new_n302_), .A4(new_n303_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n419_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n310_), .A2(KEYINPUT33), .A3(new_n312_), .A4(new_n317_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n465_), .A2(new_n428_), .A3(new_n466_), .A4(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n452_), .B1(new_n458_), .B2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n375_), .A2(new_n325_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n427_), .A2(new_n428_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT100), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n466_), .A2(new_n428_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n472_), .A2(new_n473_), .B1(new_n474_), .B2(new_n377_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n469_), .A2(new_n375_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n435_), .B1(new_n476_), .B2(new_n269_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n252_), .B1(new_n250_), .B2(new_n254_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n261_), .A2(new_n251_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n265_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n255_), .A2(new_n262_), .A3(new_n266_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n310_), .A2(new_n312_), .A3(new_n317_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n483_), .A2(KEYINPUT33), .B1(new_n462_), .B2(new_n464_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n418_), .A2(new_n419_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n484_), .A2(new_n455_), .A3(new_n485_), .A4(new_n457_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n376_), .B1(new_n486_), .B2(new_n452_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n432_), .A2(new_n375_), .A3(new_n325_), .ZN(new_n488_));
  OAI211_X1 g287(.A(KEYINPUT101), .B(new_n482_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n434_), .B1(new_n477_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT10), .B(G99gat), .Z(new_n495_));
  INV_X1    g294(.A(G106gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G85gat), .B(G92gat), .Z(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT9), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT64), .B(G85gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT9), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(G92gat), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n494_), .A2(new_n497_), .A3(new_n499_), .A4(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  NOR2_X1   g304(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n498_), .B1(new_n507_), .B2(new_n493_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n508_), .A2(KEYINPUT8), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(KEYINPUT8), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n504_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n514_));
  XOR2_X1   g313(.A(G71gat), .B(G78gat), .Z(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n514_), .A2(new_n515_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(KEYINPUT66), .B(KEYINPUT12), .C1(new_n511_), .C2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n508_), .B(KEYINPUT8), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n503_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n518_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n519_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G230gat), .A2(G233gat), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n520_), .A2(new_n518_), .A3(new_n503_), .ZN(new_n527_));
  OR2_X1    g326(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n525_), .A2(new_n526_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n527_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n511_), .A2(new_n518_), .ZN(new_n533_));
  OAI211_X1 g332(.A(G230gat), .B(G233gat), .C1(new_n532_), .C2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G120gat), .B(G148gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G176gat), .B(G204gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT67), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n535_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT13), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT74), .B(G1gat), .ZN(new_n545_));
  INV_X1    g344(.A(G8gat), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT14), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G15gat), .B(G22gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G1gat), .B(G8gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n547_), .A2(new_n548_), .A3(new_n550_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G29gat), .B(G36gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G43gat), .B(G50gat), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n556_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT15), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n557_), .A2(KEYINPUT15), .A3(new_n558_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n562_), .A2(new_n553_), .A3(new_n552_), .A4(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT75), .Z(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(new_n564_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT76), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT76), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n560_), .A2(new_n564_), .A3(new_n569_), .A4(new_n566_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n554_), .A2(new_n559_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n559_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n553_), .B2(new_n552_), .ZN(new_n573_));
  OAI211_X1 g372(.A(G229gat), .B(G233gat), .C1(new_n571_), .C2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n568_), .A2(new_n570_), .A3(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G169gat), .B(G197gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n568_), .A2(new_n570_), .A3(new_n574_), .A4(new_n578_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n544_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n490_), .A2(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n562_), .A2(new_n563_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n521_), .A2(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n586_), .A2(KEYINPUT70), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT35), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n521_), .B2(new_n572_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT71), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI211_X1 g394(.A(KEYINPUT71), .B(new_n592_), .C1(new_n521_), .C2(new_n572_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n586_), .A2(KEYINPUT70), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n587_), .A2(new_n595_), .A3(new_n596_), .A4(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n590_), .A2(new_n591_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n586_), .B1(new_n591_), .B2(new_n590_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n601_), .A2(new_n593_), .ZN(new_n602_));
  XOR2_X1   g401(.A(G134gat), .B(G162gat), .Z(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT36), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT72), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n600_), .A2(new_n602_), .A3(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n600_), .A2(new_n602_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n605_), .B(new_n606_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n609_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(new_n609_), .B2(KEYINPUT73), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  OAI221_X1 g414(.A(new_n609_), .B1(KEYINPUT73), .B2(new_n613_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n518_), .B(new_n619_), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(new_n554_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT17), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT16), .ZN(new_n624_));
  XOR2_X1   g423(.A(G183gat), .B(G211gat), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n621_), .A2(new_n622_), .A3(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(KEYINPUT17), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n621_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n618_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n584_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n545_), .A3(new_n325_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT38), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n612_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n583_), .A2(new_n630_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n638_), .A2(KEYINPUT102), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(KEYINPUT102), .ZN(new_n640_));
  AOI211_X1 g439(.A(new_n637_), .B(new_n490_), .C1(new_n639_), .C2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n326_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n634_), .A2(new_n635_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n636_), .A2(new_n643_), .A3(new_n644_), .ZN(G1324gat));
  NAND3_X1  g444(.A1(new_n633_), .A2(new_n546_), .A3(new_n432_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n641_), .A2(new_n432_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n648_), .B2(G8gat), .ZN(new_n649_));
  AOI211_X1 g448(.A(KEYINPUT39), .B(new_n546_), .C1(new_n641_), .C2(new_n432_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT40), .B(new_n646_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1325gat));
  OR3_X1    g454(.A1(new_n632_), .A2(G15gat), .A3(new_n482_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n641_), .A2(new_n269_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT41), .B1(new_n657_), .B2(G15gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n656_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(KEYINPUT103), .B(new_n656_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1326gat));
  OAI21_X1  g463(.A(G22gat), .B1(new_n642_), .B2(new_n375_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT42), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n375_), .A2(G22gat), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT104), .Z(new_n668_));
  OAI21_X1  g467(.A(new_n666_), .B1(new_n632_), .B2(new_n668_), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n612_), .A2(new_n629_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n584_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G29gat), .B1(new_n671_), .B2(new_n325_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n583_), .A2(new_n629_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  INV_X1    g473(.A(new_n434_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n469_), .A2(new_n375_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n470_), .A2(new_n475_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT101), .B1(new_n678_), .B2(new_n482_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n489_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n675_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n674_), .B1(new_n681_), .B2(new_n618_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n490_), .A2(KEYINPUT43), .A3(new_n617_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n673_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT44), .B(new_n673_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n325_), .A2(G29gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n672_), .B1(new_n688_), .B2(new_n689_), .ZN(G1328gat));
  NAND3_X1  g489(.A1(new_n686_), .A2(new_n432_), .A3(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G36gat), .ZN(new_n692_));
  NOR2_X1   g491(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n693_));
  INV_X1    g492(.A(new_n583_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n475_), .A2(G36gat), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n681_), .A2(new_n694_), .A3(new_n670_), .A4(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT105), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n696_), .A2(KEYINPUT105), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT45), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n696_), .A2(KEYINPUT105), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT45), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n697_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n693_), .B1(new_n700_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT107), .Z(new_n706_));
  AND3_X1   g505(.A1(new_n692_), .A2(new_n704_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n692_), .B2(new_n704_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1329gat));
  NOR2_X1   g508(.A1(new_n482_), .A2(new_n243_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n686_), .A2(new_n687_), .A3(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT108), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n686_), .A2(new_n713_), .A3(new_n687_), .A4(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n671_), .A2(new_n269_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n243_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n712_), .A2(new_n714_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT47), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n712_), .A2(new_n719_), .A3(new_n714_), .A4(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1330gat));
  AOI21_X1  g520(.A(G50gat), .B1(new_n671_), .B2(new_n376_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n376_), .A2(G50gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n688_), .B2(new_n723_), .ZN(G1331gat));
  NOR3_X1   g523(.A1(new_n490_), .A2(new_n582_), .A3(new_n544_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n629_), .A3(new_n612_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G57gat), .B1(new_n726_), .B2(new_n326_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n725_), .A2(new_n629_), .A3(new_n617_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n326_), .A2(G57gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n728_), .B2(new_n729_), .ZN(G1332gat));
  OR3_X1    g529(.A1(new_n728_), .A2(G64gat), .A3(new_n475_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G64gat), .B1(new_n726_), .B2(new_n475_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n732_), .A2(KEYINPUT110), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(KEYINPUT110), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n731_), .B1(new_n736_), .B2(new_n737_), .ZN(G1333gat));
  OAI21_X1  g537(.A(G71gat), .B1(new_n726_), .B2(new_n482_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT49), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n482_), .A2(G71gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n740_), .B1(new_n728_), .B2(new_n741_), .ZN(G1334gat));
  OAI21_X1  g541(.A(G78gat), .B1(new_n726_), .B2(new_n375_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT50), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n375_), .A2(G78gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n728_), .B2(new_n745_), .ZN(G1335gat));
  AND2_X1   g545(.A1(new_n725_), .A2(new_n670_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n325_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n682_), .A2(new_n683_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n544_), .A2(new_n629_), .A3(new_n582_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n325_), .A2(new_n500_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n748_), .B1(new_n752_), .B2(new_n753_), .ZN(G1336gat));
  OAI21_X1  g553(.A(G92gat), .B1(new_n751_), .B2(new_n475_), .ZN(new_n755_));
  INV_X1    g554(.A(G92gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n747_), .A2(new_n756_), .A3(new_n432_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1337gat));
  NAND4_X1  g557(.A1(new_n725_), .A2(new_n495_), .A3(new_n269_), .A4(new_n670_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(KEYINPUT111), .B2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n749_), .A2(new_n269_), .A3(new_n750_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(G99gat), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n760_), .A2(KEYINPUT111), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n763_), .B(new_n764_), .ZN(G1338gat));
  NAND3_X1  g564(.A1(new_n747_), .A2(new_n496_), .A3(new_n376_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n376_), .B(new_n750_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n767_), .A2(new_n768_), .A3(G106gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n767_), .B2(G106gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g571(.A(new_n529_), .B1(new_n519_), .B2(new_n524_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT55), .B1(new_n773_), .B2(new_n526_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n531_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(KEYINPUT55), .A3(new_n526_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n540_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  INV_X1    g578(.A(new_n540_), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n779_), .B(new_n780_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n778_), .A2(new_n781_), .A3(KEYINPUT114), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n777_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n540_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n531_), .A2(new_n534_), .A3(new_n780_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(new_n582_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(new_n582_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n783_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n566_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n560_), .A2(new_n564_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n790_), .B(new_n579_), .C1(new_n791_), .C2(new_n566_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n581_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(new_n795_));
  OAI22_X1  g594(.A1(new_n782_), .A2(new_n789_), .B1(new_n542_), .B2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(KEYINPUT57), .A3(new_n612_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n542_), .A2(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n777_), .A2(new_n540_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n779_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n777_), .A2(KEYINPUT56), .A3(new_n540_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n801_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n783_), .A2(new_n788_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n799_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n798_), .B1(new_n806_), .B2(new_n637_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n784_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n795_), .A2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT58), .B(new_n809_), .C1(new_n778_), .C2(new_n781_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n618_), .A2(new_n810_), .A3(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n797_), .A2(new_n807_), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n630_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n542_), .A2(KEYINPUT13), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n542_), .A2(KEYINPUT13), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n582_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(new_n617_), .A3(new_n629_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n821_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n819_), .A2(new_n617_), .A3(new_n629_), .A4(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n816_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n269_), .A2(new_n325_), .A3(new_n433_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G113gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n582_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n582_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT59), .B1(new_n827_), .B2(new_n829_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n825_), .B1(new_n815_), .B2(new_n630_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n828_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n834_), .B1(new_n836_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n833_), .B1(new_n841_), .B2(new_n832_), .ZN(G1340gat));
  INV_X1    g641(.A(G120gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n544_), .B2(KEYINPUT60), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n831_), .B(new_n844_), .C1(KEYINPUT60), .C2(new_n843_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n544_), .B1(new_n836_), .B2(new_n840_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n843_), .ZN(G1341gat));
  XOR2_X1   g646(.A(KEYINPUT117), .B(G127gat), .Z(new_n848_));
  NOR2_X1   g647(.A1(new_n630_), .A2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n835_), .B2(new_n839_), .ZN(new_n850_));
  INV_X1    g649(.A(G127gat), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT116), .B(new_n851_), .C1(new_n830_), .C2(new_n630_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n837_), .A2(new_n630_), .A3(new_n828_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(G127gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n850_), .A2(new_n852_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n850_), .A2(new_n852_), .A3(new_n855_), .A4(KEYINPUT118), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1342gat));
  AOI21_X1  g659(.A(G134gat), .B1(new_n831_), .B2(new_n637_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n836_), .A2(new_n840_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n863_), .A2(G134gat), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(G134gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n617_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n861_), .B1(new_n862_), .B2(new_n866_), .ZN(G1343gat));
  NOR3_X1   g666(.A1(new_n432_), .A2(new_n326_), .A3(new_n375_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n827_), .A2(new_n482_), .A3(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n834_), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n544_), .ZN(new_n872_));
  XOR2_X1   g671(.A(new_n872_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g672(.A1(new_n869_), .A2(new_n630_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT61), .B(G155gat), .Z(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  OAI21_X1  g675(.A(G162gat), .B1(new_n869_), .B2(new_n617_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n612_), .A2(G162gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n869_), .B2(new_n878_), .ZN(G1347gat));
  XNOR2_X1  g678(.A(KEYINPUT120), .B(KEYINPUT62), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n837_), .A2(new_n475_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n482_), .A2(new_n376_), .A3(new_n325_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n834_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n880_), .B1(new_n884_), .B2(new_n204_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n880_), .ZN(new_n886_));
  OAI211_X1 g685(.A(G169gat), .B(new_n886_), .C1(new_n883_), .C2(new_n834_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n884_), .A2(new_n387_), .A3(new_n382_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n885_), .A2(new_n887_), .A3(new_n888_), .ZN(G1348gat));
  NOR2_X1   g688(.A1(new_n883_), .A2(new_n544_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n205_), .ZN(G1349gat));
  NOR2_X1   g690(.A1(new_n883_), .A2(new_n630_), .ZN(new_n892_));
  MUX2_X1   g691(.A(G183gat), .B(new_n221_), .S(new_n892_), .Z(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n883_), .B2(new_n617_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n637_), .A2(new_n217_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n883_), .B2(new_n895_), .ZN(G1351gat));
  NAND2_X1  g695(.A1(new_n482_), .A2(new_n470_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT121), .ZN(new_n898_));
  NOR4_X1   g697(.A1(new_n837_), .A2(new_n834_), .A3(new_n475_), .A4(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT123), .B1(new_n899_), .B2(KEYINPUT122), .ZN(new_n900_));
  AOI21_X1  g699(.A(G197gat), .B1(new_n899_), .B2(KEYINPUT122), .ZN(new_n901_));
  INV_X1    g700(.A(new_n898_), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n827_), .A2(new_n582_), .A3(new_n432_), .A4(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n900_), .A2(new_n901_), .A3(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n899_), .A2(KEYINPUT122), .ZN(new_n908_));
  INV_X1    g707(.A(G197gat), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n900_), .A2(new_n906_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n907_), .A2(new_n910_), .ZN(G1352gat));
  NAND2_X1  g710(.A1(new_n881_), .A2(new_n902_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n544_), .ZN(new_n913_));
  INV_X1    g712(.A(G204gat), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(KEYINPUT124), .ZN(new_n915_));
  XOR2_X1   g714(.A(new_n913_), .B(new_n915_), .Z(G1353gat));
  NOR2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n912_), .B2(new_n630_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  OAI211_X1 g719(.A(KEYINPUT126), .B(new_n917_), .C1(new_n912_), .C2(new_n630_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n837_), .A2(new_n475_), .A3(new_n898_), .ZN(new_n922_));
  XOR2_X1   g721(.A(KEYINPUT63), .B(G211gat), .Z(new_n923_));
  NAND3_X1  g722(.A1(new_n922_), .A2(new_n629_), .A3(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT125), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n922_), .A2(new_n926_), .A3(new_n629_), .A4(new_n923_), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n920_), .A2(new_n921_), .B1(new_n925_), .B2(new_n927_), .ZN(G1354gat));
  NAND2_X1  g727(.A1(new_n922_), .A2(new_n637_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT127), .B(G218gat), .Z(new_n930_));
  NOR2_X1   g729(.A1(new_n617_), .A2(new_n930_), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n929_), .A2(new_n930_), .B1(new_n922_), .B2(new_n931_), .ZN(G1355gat));
endmodule


