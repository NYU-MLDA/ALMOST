//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n911_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT78), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT78), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(G169gat), .B2(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n203_), .B1(new_n210_), .B2(KEYINPUT24), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT80), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(KEYINPUT24), .A3(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT25), .B(G183gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT26), .B(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT79), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n214_), .A2(KEYINPUT79), .A3(new_n217_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n212_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n213_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT81), .B(G176gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G169gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n222_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G71gat), .B(G99gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(G43gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n229_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n232_), .B(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(G15gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT31), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n236_), .B(new_n241_), .Z(new_n242_));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n243_));
  INV_X1    g042(.A(new_n235_), .ZN(new_n244_));
  AND2_X1   g043(.A1(G141gat), .A2(G148gat), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n245_), .A2(KEYINPUT2), .ZN(new_n246_));
  NOR2_X1   g045(.A1(G141gat), .A2(G148gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(KEYINPUT2), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n246_), .A2(new_n249_), .A3(new_n250_), .A4(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G155gat), .A2(G162gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT82), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(G155gat), .A3(G162gat), .ZN(new_n256_));
  INV_X1    g055(.A(G155gat), .ZN(new_n257_));
  INV_X1    g056(.A(G162gat), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n254_), .A2(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n254_), .A2(new_n256_), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n261_), .A2(KEYINPUT1), .B1(new_n257_), .B2(new_n258_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(KEYINPUT1), .B2(new_n261_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n245_), .A2(new_n247_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(KEYINPUT83), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT83), .B1(new_n263_), .B2(new_n264_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n260_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n244_), .B1(new_n268_), .B2(KEYINPUT98), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n263_), .A2(new_n264_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT83), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n265_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT98), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n273_), .A2(new_n274_), .A3(new_n260_), .A4(new_n235_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n243_), .B1(new_n269_), .B2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n268_), .A2(new_n243_), .A3(new_n235_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G225gat), .A2(G233gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT99), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT99), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(new_n276_), .B2(new_n280_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n269_), .A2(new_n275_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n278_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G1gat), .B(G29gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(G85gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT0), .B(G57gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(new_n292_), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n281_), .A2(KEYINPUT99), .B1(new_n285_), .B2(new_n278_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n294_), .A2(KEYINPUT100), .A3(new_n291_), .A4(new_n284_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT27), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT95), .ZN(new_n298_));
  INV_X1    g097(.A(G197gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G204gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT86), .ZN(new_n301_));
  INV_X1    g100(.A(G204gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G197gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT85), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n302_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(KEYINPUT87), .B(KEYINPUT21), .Z(new_n308_));
  OR3_X1    g107(.A1(new_n301_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G211gat), .B(G218gat), .Z(new_n310_));
  NAND2_X1  g109(.A1(new_n300_), .A2(new_n303_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(KEYINPUT21), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n301_), .A2(new_n307_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n310_), .A2(KEYINPUT21), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT88), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n309_), .A2(new_n312_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT88), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n220_), .A2(new_n221_), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n323_), .A2(new_n212_), .B1(new_n223_), .B2(new_n227_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n298_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G226gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n229_), .A2(KEYINPUT95), .A3(new_n318_), .A4(new_n321_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT94), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n223_), .B(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n226_), .B(KEYINPUT93), .Z(new_n333_));
  AOI21_X1  g132(.A(new_n224_), .B1(new_n333_), .B2(new_n225_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n210_), .A2(KEYINPUT92), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(new_n209_), .B2(new_n213_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n338_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n339_), .A2(new_n203_), .A3(new_n217_), .A4(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n335_), .A2(new_n319_), .A3(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n342_), .A2(KEYINPUT20), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n325_), .A2(new_n329_), .A3(new_n330_), .A4(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n335_), .A2(new_n341_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n317_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n319_), .B(KEYINPUT88), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n346_), .B(KEYINPUT20), .C1(new_n347_), .C2(new_n229_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n328_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(new_n349_), .A3(KEYINPUT96), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n330_), .A2(new_n343_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT96), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n329_), .A4(new_n325_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G8gat), .B(G36gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n350_), .A2(new_n353_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n297_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n350_), .A2(new_n353_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n358_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n325_), .A2(new_n330_), .A3(new_n343_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n328_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n328_), .B2(new_n348_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n359_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(KEYINPUT27), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n294_), .A2(new_n291_), .A3(new_n284_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT100), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n296_), .A2(new_n363_), .A3(new_n370_), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n268_), .A2(KEYINPUT29), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n317_), .ZN(new_n376_));
  AND2_X1   g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n322_), .A2(new_n377_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT89), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n375_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n380_), .B1(new_n379_), .B2(new_n375_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n378_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G78gat), .B(G106gat), .Z(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n384_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n378_), .B(new_n386_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n268_), .A2(KEYINPUT29), .ZN(new_n389_));
  XOR2_X1   g188(.A(G22gat), .B(G50gat), .Z(new_n390_));
  OR2_X1    g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n390_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n391_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n393_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n388_), .B(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n242_), .B1(new_n374_), .B2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n373_), .A2(new_n295_), .A3(new_n293_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n348_), .A2(new_n328_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n401_), .B1(new_n328_), .B2(new_n366_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n358_), .A2(KEYINPUT32), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n364_), .B2(new_n403_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n397_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n388_), .B(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n361_), .A2(new_n362_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n294_), .A2(KEYINPUT33), .A3(new_n291_), .A4(new_n284_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n371_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n291_), .B1(new_n285_), .B2(new_n279_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n277_), .A2(new_n278_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n413_), .B1(new_n276_), .B2(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n409_), .A2(new_n410_), .A3(new_n412_), .A4(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n406_), .A2(new_n408_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT101), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT27), .B1(new_n365_), .B2(new_n360_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT27), .B1(new_n402_), .B2(new_n358_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n420_), .A2(new_n362_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n418_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n363_), .A2(new_n370_), .A3(KEYINPUT101), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n398_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n242_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(new_n400_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n399_), .A2(new_n417_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT76), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G29gat), .B(G36gat), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n429_), .A2(KEYINPUT68), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(KEYINPUT68), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G43gat), .B(G50gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n430_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G15gat), .B(G22gat), .ZN(new_n438_));
  INV_X1    g237(.A(G1gat), .ZN(new_n439_));
  INV_X1    g238(.A(G8gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT14), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G1gat), .B(G8gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n437_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n437_), .A2(new_n444_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n428_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n430_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n433_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n444_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(new_n445_), .A3(KEYINPUT76), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G229gat), .A2(G233gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT15), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n458_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n435_), .A2(KEYINPUT15), .A3(new_n436_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n444_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n447_), .A2(new_n457_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n455_), .A2(new_n457_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G113gat), .B(G141gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT77), .ZN(new_n466_));
  XOR2_X1   g265(.A(G169gat), .B(G197gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n464_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n427_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT75), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G190gat), .B(G218gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT71), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G134gat), .B(G162gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT36), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT73), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT70), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G232gat), .A2(G233gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n481_), .B(KEYINPUT34), .Z(new_n482_));
  INV_X1    g281(.A(KEYINPUT35), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G85gat), .ZN(new_n485_));
  INV_X1    g284(.A(G92gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G85gat), .A2(G92gat), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT6), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(G99gat), .A3(G106gat), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT7), .ZN(new_n495_));
  INV_X1    g294(.A(G99gat), .ZN(new_n496_));
  INV_X1    g295(.A(G106gat), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .A4(KEYINPUT64), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT64), .ZN(new_n499_));
  OAI22_X1  g298(.A1(new_n499_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n489_), .B1(new_n494_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT8), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OAI211_X1 g303(.A(KEYINPUT8), .B(new_n489_), .C1(new_n494_), .C2(new_n501_), .ZN(new_n505_));
  OR2_X1    g304(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n497_), .A3(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n487_), .A2(KEYINPUT9), .A3(new_n488_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n488_), .A2(KEYINPUT9), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n504_), .A2(new_n505_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT65), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n502_), .A2(new_n503_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(KEYINPUT65), .A3(new_n505_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n451_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n482_), .A2(new_n483_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(KEYINPUT69), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n461_), .A2(new_n514_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT69), .B1(new_n519_), .B2(new_n520_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n480_), .B(new_n484_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n484_), .B1(new_n461_), .B2(new_n514_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(new_n520_), .A3(new_n519_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT72), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n526_), .A2(KEYINPUT72), .A3(new_n520_), .A4(new_n519_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n525_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n519_), .A2(new_n520_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT69), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n480_), .B1(new_n536_), .B2(new_n484_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n479_), .B1(new_n532_), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n484_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT70), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n476_), .A2(new_n477_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n540_), .A2(new_n541_), .A3(new_n525_), .A4(new_n531_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n472_), .B1(new_n538_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n538_), .B2(new_n542_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT37), .ZN(new_n546_));
  OAI22_X1  g345(.A1(KEYINPUT74), .A2(new_n543_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n538_), .A2(new_n542_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT75), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(new_n544_), .A3(KEYINPUT37), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(G78gat), .ZN(new_n555_));
  INV_X1    g354(.A(G78gat), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n556_), .A3(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(G64gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(G57gat), .ZN(new_n560_));
  INV_X1    g359(.A(G57gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(G64gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n562_), .A3(KEYINPUT11), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(new_n563_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n560_), .A2(new_n562_), .A3(KEYINPUT11), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT11), .B1(new_n560_), .B2(new_n562_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n555_), .B(new_n557_), .C1(new_n565_), .C2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n516_), .A2(new_n569_), .A3(new_n518_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT67), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT12), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n571_), .B1(new_n514_), .B2(new_n573_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n514_), .A2(new_n573_), .A3(new_n571_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n570_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n516_), .A2(new_n518_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT12), .B1(new_n577_), .B2(new_n568_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G230gat), .A2(G233gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n514_), .A2(new_n515_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT65), .B1(new_n517_), .B2(new_n505_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n568_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n570_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n580_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n581_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G120gat), .B(G148gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT5), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G176gat), .B(G204gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n581_), .A2(new_n587_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT13), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n593_), .A2(KEYINPUT13), .A3(new_n595_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n444_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n569_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT16), .ZN(new_n608_));
  XOR2_X1   g407(.A(G183gat), .B(G211gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n605_), .B1(new_n606_), .B2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n606_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n604_), .A2(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n551_), .A2(new_n601_), .A3(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n471_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n439_), .A3(new_n400_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n427_), .A2(new_n548_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n614_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n600_), .A2(new_n469_), .A3(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT102), .Z(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n400_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G1gat), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n617_), .A2(new_n618_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n619_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT103), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n619_), .A2(new_n630_), .A3(new_n626_), .A4(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(G1324gat));
  XNOR2_X1  g431(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n422_), .A2(new_n423_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(G8gat), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n471_), .A2(new_n615_), .A3(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT104), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n363_), .A2(new_n370_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n398_), .B1(new_n638_), .B2(new_n400_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n417_), .A2(new_n639_), .A3(new_n425_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n424_), .A2(new_n426_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n634_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n548_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n642_), .A2(new_n623_), .A3(new_n643_), .A4(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n646_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n647_), .A2(new_n648_), .A3(KEYINPUT39), .A4(G8gat), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n637_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(G8gat), .A3(new_n648_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT39), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n633_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n654_));
  AND4_X1   g453(.A1(new_n653_), .A2(new_n637_), .A3(new_n649_), .A4(new_n633_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1325gat));
  OAI21_X1  g455(.A(G15gat), .B1(new_n624_), .B2(new_n425_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n616_), .A2(new_n238_), .A3(new_n242_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(KEYINPUT107), .A3(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1326gat));
  OAI21_X1  g464(.A(G22gat), .B1(new_n624_), .B2(new_n408_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT42), .ZN(new_n667_));
  INV_X1    g466(.A(G22gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n616_), .A2(new_n668_), .A3(new_n398_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1327gat));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n601_), .A2(new_n470_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n614_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n547_), .A2(new_n550_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n427_), .A2(KEYINPUT43), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n642_), .B2(new_n551_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n676_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT43), .B1(new_n427_), .B2(new_n675_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n642_), .A2(new_n677_), .A3(new_n551_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(KEYINPUT44), .A3(new_n674_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n681_), .A2(new_n400_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G29gat), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n548_), .A2(new_n614_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n601_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n471_), .A2(new_n689_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n690_), .A2(G29gat), .A3(new_n625_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n671_), .B1(new_n687_), .B2(new_n692_), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT108), .B(new_n691_), .C1(new_n686_), .C2(G29gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1328gat));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  INV_X1    g495(.A(G36gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT44), .B1(new_n684_), .B2(new_n674_), .ZN(new_n698_));
  AOI211_X1 g497(.A(new_n680_), .B(new_n673_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n697_), .B1(new_n700_), .B2(new_n643_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n471_), .A2(new_n697_), .A3(new_n643_), .A4(new_n689_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT45), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n696_), .B1(new_n701_), .B2(new_n704_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n698_), .A2(new_n699_), .A3(new_n634_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT46), .B(new_n703_), .C1(new_n706_), .C2(new_n697_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1329gat));
  NAND4_X1  g507(.A1(new_n681_), .A2(G43gat), .A3(new_n242_), .A4(new_n685_), .ZN(new_n709_));
  INV_X1    g508(.A(G43gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n710_), .B1(new_n690_), .B2(new_n425_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g512(.A1(new_n690_), .A2(G50gat), .A3(new_n408_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n700_), .A2(KEYINPUT109), .A3(new_n398_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G50gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT109), .B1(new_n700_), .B2(new_n398_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n714_), .B1(new_n716_), .B2(new_n717_), .ZN(G1331gat));
  NOR2_X1   g517(.A1(new_n469_), .A2(new_n614_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n620_), .A2(new_n601_), .A3(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G57gat), .B1(new_n720_), .B2(new_n625_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n427_), .A2(new_n469_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n675_), .A2(new_n601_), .A3(new_n621_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n723_), .A2(new_n724_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n722_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n400_), .A2(new_n561_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n721_), .B1(new_n727_), .B2(new_n728_), .ZN(G1332gat));
  OAI21_X1  g528(.A(G64gat), .B1(new_n720_), .B2(new_n634_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT48), .ZN(new_n731_));
  INV_X1    g530(.A(new_n727_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n559_), .A3(new_n643_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1333gat));
  OAI21_X1  g533(.A(G71gat), .B1(new_n720_), .B2(new_n425_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT49), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n425_), .A2(G71gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT111), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n736_), .B1(new_n727_), .B2(new_n738_), .ZN(G1334gat));
  OAI21_X1  g538(.A(G78gat), .B1(new_n720_), .B2(new_n408_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT50), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n732_), .A2(new_n556_), .A3(new_n398_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1335gat));
  NOR3_X1   g542(.A1(new_n600_), .A2(new_n469_), .A3(new_n621_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n684_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745_), .B2(new_n625_), .ZN(new_n746_));
  NOR4_X1   g545(.A1(new_n427_), .A2(new_n469_), .A3(new_n600_), .A4(new_n688_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n485_), .A3(new_n400_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1336gat));
  OAI21_X1  g548(.A(G92gat), .B1(new_n745_), .B2(new_n634_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n747_), .A2(new_n486_), .A3(new_n643_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1337gat));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n242_), .B(new_n744_), .C1(new_n676_), .C2(new_n678_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n242_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n754_), .A2(G99gat), .B1(new_n747_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n757_));
  AOI211_X1 g556(.A(new_n753_), .B(KEYINPUT51), .C1(new_n756_), .C2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n757_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT112), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n756_), .B2(new_n753_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n758_), .B1(new_n760_), .B2(new_n762_), .ZN(G1338gat));
  NAND3_X1  g562(.A1(new_n747_), .A2(new_n497_), .A3(new_n398_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n684_), .A2(new_n398_), .A3(new_n744_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(G106gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(G106gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT53), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n764_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1339gat));
  NAND2_X1  g572(.A1(new_n455_), .A2(new_n456_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n447_), .A2(new_n456_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n468_), .B1(new_n775_), .B2(new_n462_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n464_), .A2(new_n468_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n596_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n469_), .A2(new_n595_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n582_), .A2(new_n583_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n514_), .A2(new_n573_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT67), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n514_), .A2(new_n573_), .A3(new_n571_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n780_), .A2(new_n569_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n584_), .A2(new_n572_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n784_), .A2(KEYINPUT55), .A3(new_n580_), .A4(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n579_), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n580_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n782_), .A2(new_n783_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n569_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n790_), .B(new_n570_), .C1(KEYINPUT12), .C2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n586_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(new_n792_), .B2(new_n586_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n788_), .A2(new_n789_), .A3(new_n793_), .A4(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n592_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n592_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n779_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n778_), .B1(new_n801_), .B2(KEYINPUT117), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n469_), .A2(new_n595_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n592_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT56), .B1(new_n796_), .B2(new_n592_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n803_), .B(KEYINPUT117), .C1(new_n804_), .C2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n644_), .B1(new_n802_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n548_), .A2(new_n809_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n802_), .B2(new_n807_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n777_), .A2(new_n595_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n777_), .A2(KEYINPUT118), .A3(new_n595_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820_));
  AOI22_X1  g619(.A1(new_n817_), .A2(new_n818_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n799_), .A2(new_n800_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n819_), .B1(KEYINPUT119), .B2(new_n820_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n821_), .A2(new_n822_), .A3(new_n824_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n551_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n803_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n829_), .A2(new_n830_), .B1(new_n596_), .B2(new_n777_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n806_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(KEYINPUT121), .A3(new_n811_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n810_), .A2(new_n814_), .A3(new_n828_), .A4(new_n833_), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n598_), .A2(new_n719_), .A3(new_n599_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n675_), .B2(new_n839_), .ZN(new_n840_));
  AOI211_X1 g639(.A(KEYINPUT115), .B(new_n838_), .C1(new_n547_), .C2(new_n550_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n836_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT115), .B1(new_n551_), .B2(new_n838_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n675_), .A2(new_n839_), .A3(new_n837_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n835_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n834_), .A2(new_n614_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n424_), .A2(new_n400_), .A3(new_n242_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(G113gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n469_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n847_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT121), .B1(new_n832_), .B2(new_n811_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n811_), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n813_), .B(new_n855_), .C1(new_n831_), .C2(new_n806_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n826_), .A2(new_n827_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n551_), .A2(new_n858_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n621_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n845_), .A2(new_n842_), .ZN(new_n861_));
  OAI211_X1 g660(.A(KEYINPUT59), .B(new_n853_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n470_), .B1(new_n852_), .B2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n850_), .B1(new_n863_), .B2(new_n849_), .ZN(G1340gat));
  INV_X1    g663(.A(G120gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n600_), .B2(KEYINPUT60), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n865_), .B2(KEYINPUT60), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n848_), .B(new_n869_), .C1(KEYINPUT122), .C2(new_n866_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n600_), .B1(new_n852_), .B2(new_n862_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n865_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  OAI211_X1 g673(.A(KEYINPUT123), .B(new_n870_), .C1(new_n871_), .C2(new_n865_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1341gat));
  INV_X1    g675(.A(G127gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n848_), .A2(new_n877_), .A3(new_n621_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n614_), .B1(new_n852_), .B2(new_n862_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n877_), .ZN(G1342gat));
  INV_X1    g679(.A(G134gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n848_), .A2(new_n881_), .A3(new_n548_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n675_), .B1(new_n852_), .B2(new_n862_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n881_), .ZN(G1343gat));
  NOR2_X1   g683(.A1(new_n408_), .A2(new_n242_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NOR4_X1   g685(.A1(new_n846_), .A2(new_n643_), .A3(new_n625_), .A4(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n469_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT124), .B(G141gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1344gat));
  NAND2_X1  g689(.A1(new_n887_), .A2(new_n601_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g691(.A1(new_n887_), .A2(new_n621_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT61), .B(G155gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1346gat));
  NAND3_X1  g694(.A1(new_n887_), .A2(new_n258_), .A3(new_n548_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n887_), .A2(new_n551_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n258_), .ZN(G1347gat));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n426_), .A2(new_n408_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n846_), .A2(new_n634_), .A3(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n470_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n899_), .B1(new_n903_), .B2(new_n204_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n333_), .ZN(new_n905_));
  OAI211_X1 g704(.A(KEYINPUT62), .B(G169gat), .C1(new_n902_), .C2(new_n470_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n904_), .A2(new_n905_), .A3(new_n906_), .ZN(G1348gat));
  NOR3_X1   g706(.A1(new_n902_), .A2(new_n205_), .A3(new_n600_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n901_), .A2(new_n601_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n225_), .B2(new_n909_), .ZN(G1349gat));
  NAND2_X1  g709(.A1(new_n901_), .A2(new_n621_), .ZN(new_n911_));
  MUX2_X1   g710(.A(new_n215_), .B(G183gat), .S(new_n911_), .Z(G1350gat));
  NAND3_X1  g711(.A1(new_n901_), .A2(new_n216_), .A3(new_n548_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(G190gat), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n915_), .B1(new_n901_), .B2(new_n551_), .ZN(new_n916_));
  OAI21_X1  g715(.A(KEYINPUT125), .B1(new_n914_), .B2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n916_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n918_), .A2(new_n919_), .A3(new_n913_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n917_), .A2(new_n920_), .ZN(G1351gat));
  NOR2_X1   g720(.A1(new_n886_), .A2(new_n400_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n643_), .B(new_n922_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n470_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(new_n299_), .ZN(G1352gat));
  NOR2_X1   g724(.A1(new_n923_), .A2(new_n600_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(new_n302_), .ZN(G1353gat));
  NOR2_X1   g726(.A1(new_n923_), .A2(new_n614_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n928_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT63), .B(G211gat), .Z(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n928_), .B2(new_n930_), .ZN(G1354gat));
  OR2_X1    g730(.A1(new_n644_), .A2(G218gat), .ZN(new_n932_));
  OR2_X1    g731(.A1(new_n923_), .A2(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(G218gat), .B1(new_n923_), .B2(new_n675_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n933_), .A2(KEYINPUT126), .A3(new_n934_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1355gat));
endmodule


