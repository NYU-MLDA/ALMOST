//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_;
  XNOR2_X1  g000(.A(KEYINPUT68), .B(G71gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G78gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n204_));
  INV_X1    g003(.A(G78gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G64gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G57gat), .ZN(new_n209_));
  INV_X1    g008(.A(G57gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G64gat), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT11), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT11), .B1(new_n209_), .B2(new_n211_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n203_), .B(new_n207_), .C1(new_n212_), .C2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT11), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n205_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n220_));
  INV_X1    g019(.A(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G85gat), .ZN(new_n224_));
  INV_X1    g023(.A(G92gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(KEYINPUT9), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT6), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n230_), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(KEYINPUT6), .ZN(new_n233_));
  OAI22_X1  g032(.A1(new_n231_), .A2(new_n233_), .B1(KEYINPUT9), .B2(new_n227_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT64), .B1(new_n229_), .B2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n227_), .A2(KEYINPUT9), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(KEYINPUT6), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n230_), .A2(G99gat), .A3(G106gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n223_), .A4(new_n228_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n226_), .A2(new_n227_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G99gat), .A2(G106gat), .ZN(new_n244_));
  AND2_X1   g043(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n245_));
  NOR2_X1   g044(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  OAI22_X1  g046(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n231_), .A2(new_n233_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n243_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT8), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n242_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n243_), .A2(KEYINPUT8), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT66), .B1(new_n231_), .B2(new_n233_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n237_), .A2(new_n238_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT67), .B1(new_n247_), .B2(new_n248_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n247_), .A2(KEYINPUT67), .A3(new_n248_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n255_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n219_), .B1(new_n254_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n235_), .A2(new_n241_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n237_), .A2(new_n238_), .A3(new_n257_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n257_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n249_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n271_), .A3(new_n262_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n255_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n219_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n266_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n264_), .A2(new_n265_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G230gat), .A2(G233gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n277_), .B(new_n279_), .C1(new_n265_), .C2(new_n264_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT12), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n264_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n266_), .A2(new_n274_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n219_), .A2(KEYINPUT70), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n214_), .A2(new_n285_), .A3(new_n218_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n283_), .A2(KEYINPUT12), .A3(new_n287_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n282_), .A2(new_n278_), .A3(new_n288_), .A4(new_n276_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n280_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G120gat), .B(G148gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT5), .ZN(new_n292_));
  XOR2_X1   g091(.A(G176gat), .B(G204gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n290_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT13), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(KEYINPUT71), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n296_), .A2(KEYINPUT71), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n295_), .B1(new_n299_), .B2(new_n297_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT72), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n298_), .A2(new_n303_), .A3(new_n300_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G1gat), .B(G8gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT77), .ZN(new_n307_));
  OR2_X1    g106(.A1(G15gat), .A2(G22gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G15gat), .A2(G22gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G1gat), .A2(G8gat), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n308_), .A2(new_n309_), .B1(KEYINPUT14), .B2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n307_), .B(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G29gat), .B(G36gat), .Z(new_n313_));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G29gat), .B(G36gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT74), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G43gat), .B(G50gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n315_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n312_), .B(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G229gat), .A2(G233gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n321_), .A2(KEYINPUT15), .A3(new_n322_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT15), .B1(new_n321_), .B2(new_n322_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n312_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n326_), .B1(new_n312_), .B2(new_n323_), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n324_), .A2(new_n326_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G113gat), .B(G141gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT78), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G169gat), .B(G197gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n333_), .B(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n305_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT80), .ZN(new_n346_));
  INV_X1    g145(.A(G176gat), .ZN(new_n347_));
  INV_X1    g146(.A(G169gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT22), .B1(new_n348_), .B2(KEYINPUT79), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n348_), .A2(KEYINPUT22), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n347_), .B(new_n349_), .C1(new_n350_), .C2(KEYINPUT79), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n346_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n345_), .A2(KEYINPUT80), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n342_), .A2(new_n344_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT24), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT25), .B(G183gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT26), .B(G190gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n356_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(KEYINPUT24), .A3(new_n352_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  OAI22_X1  g164(.A1(new_n353_), .A2(new_n354_), .B1(new_n359_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G227gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G15gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n366_), .B(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G71gat), .B(G99gat), .Z(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT82), .B(G43gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT81), .B(KEYINPUT30), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n369_), .B(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G127gat), .B(G134gat), .Z(new_n376_));
  XOR2_X1   g175(.A(G113gat), .B(G120gat), .Z(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT31), .ZN(new_n379_));
  OR3_X1    g178(.A1(new_n375_), .A2(KEYINPUT83), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n375_), .A2(KEYINPUT83), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n379_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n375_), .A2(KEYINPUT83), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n380_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G197gat), .B(G204gat), .Z(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT21), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G197gat), .B(G204gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT21), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G211gat), .B(G218gat), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n386_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  OR3_X1    g190(.A1(new_n387_), .A2(new_n390_), .A3(new_n388_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G155gat), .A2(G162gat), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G155gat), .A2(G162gat), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n400_));
  INV_X1    g199(.A(G141gat), .ZN(new_n401_));
  INV_X1    g200(.A(G148gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G141gat), .A2(G148gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT2), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n403_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT85), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n399_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n401_), .A2(new_n402_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n404_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n396_), .A2(new_n397_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT1), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n398_), .B(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n413_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n411_), .A2(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(KEYINPUT88), .B(KEYINPUT29), .Z(new_n419_));
  OAI21_X1  g218(.A(new_n393_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(G228gat), .A3(G233gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G228gat), .A2(G233gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT86), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n393_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT87), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT29), .B1(new_n411_), .B2(new_n417_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n426_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n421_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n411_), .A2(new_n417_), .A3(KEYINPUT29), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT28), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n432_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n434_), .B(new_n421_), .C1(new_n429_), .C2(new_n428_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G78gat), .B(G106gat), .Z(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT89), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G22gat), .B(G50gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n436_), .A2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n378_), .B1(new_n417_), .B2(new_n411_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n417_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n376_), .B(new_n377_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT85), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n409_), .B(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n403_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n414_), .B(new_n398_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n446_), .A2(new_n447_), .A3(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n445_), .A2(KEYINPUT4), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n378_), .B(new_n454_), .C1(new_n417_), .C2(new_n411_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n444_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G1gat), .B(G29gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(G85gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT0), .B(G57gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n444_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n462_), .B1(new_n445_), .B2(new_n452_), .ZN(new_n463_));
  OR3_X1    g262(.A1(new_n456_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n461_), .B1(new_n456_), .B2(new_n463_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n442_), .A2(new_n443_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT90), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n365_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n359_), .A2(KEYINPUT91), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n362_), .A2(KEYINPUT90), .A3(new_n364_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT91), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n355_), .A2(new_n473_), .A3(new_n358_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .A4(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n391_), .A2(new_n392_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT22), .B(G169gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n347_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n478_), .A2(KEYINPUT92), .A3(new_n352_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT92), .B1(new_n478_), .B2(new_n352_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n345_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n475_), .A2(new_n476_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT93), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n475_), .A2(new_n476_), .A3(new_n481_), .A4(KEYINPUT93), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT20), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(new_n366_), .B2(new_n393_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G226gat), .A2(G233gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT19), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n476_), .B1(new_n475_), .B2(new_n481_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT20), .B1(new_n366_), .B2(new_n393_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n491_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G8gat), .B(G36gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT18), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G64gat), .B(G92gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n495_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n501_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT27), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n493_), .A2(new_n494_), .A3(new_n490_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n491_), .B1(new_n487_), .B2(new_n482_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n504_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n502_), .A2(KEYINPUT27), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n508_), .A2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT98), .B1(new_n468_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT98), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n467_), .A2(new_n508_), .A3(new_n515_), .A4(new_n512_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n442_), .A2(new_n443_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n453_), .A2(new_n455_), .A3(new_n444_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n445_), .A2(new_n462_), .A3(new_n452_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n460_), .A3(new_n519_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n502_), .A2(new_n520_), .A3(new_n505_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n465_), .A2(KEYINPUT95), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT33), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT95), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n524_), .B(new_n461_), .C1(new_n456_), .C2(new_n463_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n522_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT96), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n522_), .A2(new_n528_), .A3(new_n523_), .A4(new_n525_), .ZN(new_n529_));
  OAI211_X1 g328(.A(KEYINPUT33), .B(new_n461_), .C1(new_n456_), .C2(new_n463_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT94), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n521_), .A2(new_n527_), .A3(new_n529_), .A4(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(KEYINPUT32), .B(new_n501_), .C1(new_n509_), .C2(new_n510_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n501_), .A2(KEYINPUT32), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n533_), .B(new_n466_), .C1(new_n503_), .C2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n517_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT97), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n514_), .B(new_n516_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n532_), .A2(new_n535_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n517_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(KEYINPUT97), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n384_), .B1(new_n538_), .B2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n513_), .B(KEYINPUT99), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n384_), .A2(new_n466_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n544_), .A2(KEYINPUT100), .A3(new_n540_), .A4(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n513_), .A2(KEYINPUT99), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT99), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n540_), .B(new_n545_), .C1(new_n547_), .C2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT100), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n546_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n339_), .B1(new_n543_), .B2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT36), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT34), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT35), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT73), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n329_), .A2(new_n283_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT75), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n254_), .A2(new_n263_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n323_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n560_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT35), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n563_), .A2(new_n567_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n565_), .A2(new_n571_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n329_), .A2(new_n283_), .B1(new_n569_), .B2(new_n568_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT75), .B1(new_n329_), .B2(new_n283_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n573_), .B(new_n567_), .C1(new_n574_), .C2(new_n562_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n557_), .A2(KEYINPUT36), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n572_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n558_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT37), .B1(new_n577_), .B2(KEYINPUT76), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT37), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n572_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT76), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n582_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n585_), .B(new_n558_), .C1(new_n577_), .C2(new_n578_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G127gat), .B(G155gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT16), .ZN(new_n590_));
  XOR2_X1   g389(.A(G183gat), .B(G211gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n312_), .B(new_n593_), .ZN(new_n594_));
  AOI211_X1 g393(.A(new_n588_), .B(new_n592_), .C1(new_n594_), .C2(new_n287_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n594_), .B2(new_n287_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n594_), .A2(new_n275_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n275_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n592_), .B(KEYINPUT17), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n587_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n554_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n466_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n603_), .A2(G1gat), .A3(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT102), .Z(new_n609_));
  NOR2_X1   g408(.A1(new_n605_), .A2(new_n607_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT103), .ZN(new_n611_));
  INV_X1    g410(.A(new_n579_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n601_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n554_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n616_), .B2(new_n604_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n609_), .A2(new_n611_), .A3(new_n617_), .ZN(G1324gat));
  NAND2_X1  g417(.A1(new_n543_), .A2(new_n553_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n339_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n544_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .A4(new_n615_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT104), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n622_), .A2(new_n623_), .A3(G8gat), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n622_), .B2(G8gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT39), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT105), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n622_), .A2(G8gat), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT104), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n622_), .A2(new_n623_), .A3(G8gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT106), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(KEYINPUT105), .B(KEYINPUT39), .C1(new_n624_), .C2(new_n625_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n630_), .A2(KEYINPUT106), .A3(new_n631_), .A4(new_n632_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n628_), .A2(new_n635_), .A3(new_n636_), .A4(new_n637_), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n603_), .A2(G8gat), .A3(new_n544_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n638_), .A2(KEYINPUT40), .A3(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1325gat));
  NOR3_X1   g443(.A1(new_n603_), .A2(G15gat), .A3(new_n384_), .ZN(new_n645_));
  INV_X1    g444(.A(G15gat), .ZN(new_n646_));
  INV_X1    g445(.A(new_n616_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n384_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n650_));
  AOI21_X1  g449(.A(new_n645_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n649_), .B2(new_n650_), .ZN(G1326gat));
  OAI21_X1  g451(.A(G22gat), .B1(new_n616_), .B2(new_n540_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n540_), .A2(G22gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n603_), .B2(new_n656_), .ZN(G1327gat));
  NOR2_X1   g456(.A1(new_n612_), .A2(new_n613_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n554_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(G29gat), .B1(new_n659_), .B2(new_n466_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n620_), .A2(new_n601_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n619_), .A2(new_n587_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT43), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n619_), .A2(new_n664_), .A3(new_n587_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n661_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n466_), .A2(G29gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n660_), .B1(new_n668_), .B2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  INV_X1    g470(.A(G36gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n668_), .B2(new_n621_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n659_), .A2(new_n672_), .A3(new_n621_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT45), .Z(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n666_), .B(KEYINPUT44), .ZN(new_n677_));
  OAI21_X1  g476(.A(G36gat), .B1(new_n677_), .B2(new_n544_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n675_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(KEYINPUT46), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n676_), .A2(new_n680_), .ZN(G1329gat));
  NAND2_X1  g480(.A1(new_n648_), .A2(G43gat), .ZN(new_n682_));
  INV_X1    g481(.A(new_n659_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n384_), .ZN(new_n684_));
  OAI22_X1  g483(.A1(new_n677_), .A2(new_n682_), .B1(G43gat), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g485(.A1(new_n683_), .A2(G50gat), .A3(new_n540_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT109), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n668_), .A2(new_n688_), .A3(new_n517_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G50gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n668_), .B2(new_n517_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1331gat));
  AOI211_X1 g491(.A(new_n338_), .B(new_n305_), .C1(new_n543_), .C2(new_n553_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(new_n615_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n210_), .B1(new_n694_), .B2(new_n466_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n602_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n696_), .A2(G57gat), .A3(new_n604_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT110), .Z(G1332gat));
  AOI21_X1  g498(.A(new_n208_), .B1(new_n694_), .B2(new_n621_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT48), .Z(new_n701_));
  NAND2_X1  g500(.A1(new_n621_), .A2(new_n208_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n696_), .B2(new_n702_), .ZN(G1333gat));
  INV_X1    g502(.A(G71gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n694_), .B2(new_n648_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT49), .Z(new_n706_));
  NAND2_X1  g505(.A1(new_n648_), .A2(new_n704_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT111), .Z(new_n708_));
  OAI21_X1  g507(.A(new_n706_), .B1(new_n696_), .B2(new_n708_), .ZN(G1334gat));
  AOI21_X1  g508(.A(new_n205_), .B1(new_n694_), .B2(new_n517_), .ZN(new_n710_));
  XOR2_X1   g509(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n517_), .A2(new_n205_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n696_), .B2(new_n713_), .ZN(G1335gat));
  NAND2_X1  g513(.A1(new_n663_), .A2(new_n665_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n305_), .A2(new_n613_), .A3(new_n338_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G85gat), .B1(new_n717_), .B2(new_n604_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n693_), .A2(new_n658_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n224_), .A3(new_n466_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(G1336gat));
  OAI21_X1  g521(.A(G92gat), .B1(new_n717_), .B2(new_n544_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n720_), .A2(new_n225_), .A3(new_n621_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1337gat));
  OAI21_X1  g524(.A(G99gat), .B1(new_n717_), .B2(new_n384_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n648_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n726_), .B(KEYINPUT113), .C1(new_n719_), .C2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g528(.A1(new_n720_), .A2(new_n221_), .A3(new_n517_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n715_), .A2(new_n517_), .A3(new_n716_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n731_), .A2(new_n732_), .A3(G106gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n731_), .B2(G106gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n735_), .B(new_n737_), .ZN(G1339gat));
  INV_X1    g537(.A(new_n338_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n602_), .A2(new_n739_), .A3(new_n301_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT54), .Z(new_n741_));
  OR2_X1    g540(.A1(new_n290_), .A2(new_n294_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n333_), .A2(new_n337_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n337_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n325_), .B1(new_n312_), .B2(new_n323_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n331_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n743_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n742_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT115), .B1(new_n289_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n286_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n285_), .B1(new_n214_), .B2(new_n218_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT12), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n276_), .B1(new_n566_), .B2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n275_), .B1(new_n266_), .B2(new_n274_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(KEYINPUT12), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(KEYINPUT55), .A4(new_n278_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n289_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n288_), .B(new_n276_), .C1(KEYINPUT12), .C2(new_n757_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n751_), .B1(new_n763_), .B2(new_n279_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n752_), .B(new_n761_), .C1(new_n762_), .C2(new_n764_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n294_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n294_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n750_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT58), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  OAI211_X1 g569(.A(KEYINPUT58), .B(new_n750_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n587_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n742_), .A2(new_n338_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n765_), .A2(new_n294_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n294_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n295_), .A2(new_n749_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT57), .B(new_n612_), .C1(new_n778_), .C2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n772_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n612_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n613_), .B1(new_n783_), .B2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n741_), .A2(new_n787_), .ZN(new_n788_));
  NOR4_X1   g587(.A1(new_n621_), .A2(new_n384_), .A3(new_n604_), .A4(new_n517_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT59), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n788_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n338_), .A2(G113gat), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT119), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n740_), .B(KEYINPUT54), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n338_), .B(new_n742_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n579_), .B1(new_n798_), .B2(new_n779_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n797_), .B1(new_n799_), .B2(KEYINPUT57), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n784_), .A2(KEYINPUT116), .A3(new_n785_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n782_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n601_), .B1(new_n802_), .B2(KEYINPUT117), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n804_), .B(new_n782_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n796_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT118), .B(new_n796_), .C1(new_n803_), .C2(new_n805_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(new_n789_), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n792_), .B(new_n795_), .C1(new_n810_), .C2(KEYINPUT59), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n808_), .A2(new_n809_), .A3(new_n789_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G113gat), .B1(new_n812_), .B2(new_n338_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT120), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n810_), .A2(KEYINPUT59), .ZN(new_n815_));
  INV_X1    g614(.A(new_n792_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n794_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT120), .ZN(new_n818_));
  INV_X1    g617(.A(G113gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n810_), .B2(new_n739_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n814_), .A2(new_n821_), .ZN(G1340gat));
  INV_X1    g621(.A(new_n305_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n816_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n810_), .B2(KEYINPUT59), .ZN(new_n825_));
  OAI21_X1  g624(.A(G120gat), .B1(new_n825_), .B2(KEYINPUT122), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827_));
  AOI211_X1 g626(.A(new_n827_), .B(new_n824_), .C1(KEYINPUT59), .C2(new_n810_), .ZN(new_n828_));
  INV_X1    g627(.A(G120gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT121), .B1(new_n829_), .B2(KEYINPUT60), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n305_), .B2(KEYINPUT60), .ZN(new_n831_));
  MUX2_X1   g630(.A(KEYINPUT121), .B(new_n830_), .S(new_n831_), .Z(new_n832_));
  OAI22_X1  g631(.A1(new_n826_), .A2(new_n828_), .B1(new_n810_), .B2(new_n832_), .ZN(G1341gat));
  INV_X1    g632(.A(G127gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n812_), .A2(new_n834_), .A3(new_n613_), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n601_), .B(new_n792_), .C1(new_n810_), .C2(KEYINPUT59), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n834_), .ZN(G1342gat));
  NAND2_X1  g636(.A1(new_n581_), .A2(new_n586_), .ZN(new_n838_));
  INV_X1    g637(.A(G134gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  AOI211_X1 g640(.A(new_n792_), .B(new_n841_), .C1(new_n810_), .C2(KEYINPUT59), .ZN(new_n842_));
  AOI21_X1  g641(.A(G134gat), .B1(new_n812_), .B2(new_n579_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT123), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n815_), .A2(new_n816_), .A3(new_n840_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n839_), .B1(new_n810_), .B2(new_n612_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n844_), .A2(new_n848_), .ZN(G1343gat));
  XNOR2_X1  g648(.A(KEYINPUT124), .B(G141gat), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n808_), .A2(new_n384_), .A3(new_n809_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n621_), .A2(new_n604_), .A3(new_n540_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n850_), .B1(new_n853_), .B2(new_n338_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n852_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n850_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n855_), .A2(new_n739_), .A3(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n854_), .A2(new_n857_), .ZN(G1344gat));
  XNOR2_X1  g657(.A(KEYINPUT125), .B(G148gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n853_), .A2(new_n823_), .A3(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n859_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n855_), .B2(new_n305_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1345gat));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  OR3_X1    g663(.A1(new_n855_), .A2(new_n601_), .A3(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n855_), .B2(new_n601_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1346gat));
  OAI21_X1  g666(.A(G162gat), .B1(new_n855_), .B2(new_n838_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n612_), .A2(G162gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n855_), .B2(new_n869_), .ZN(G1347gat));
  NAND2_X1  g669(.A1(new_n621_), .A2(new_n545_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n517_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n741_), .B2(new_n787_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n348_), .B1(new_n874_), .B2(new_n338_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n875_), .A2(KEYINPUT62), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(new_n338_), .A3(new_n477_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(KEYINPUT62), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n877_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT126), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT126), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n876_), .A2(new_n877_), .A3(new_n881_), .A4(new_n878_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1348gat));
  AOI21_X1  g682(.A(G176gat), .B1(new_n874_), .B2(new_n823_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n808_), .A2(new_n540_), .A3(new_n809_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n871_), .A2(new_n305_), .A3(new_n347_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(G1349gat));
  NOR3_X1   g686(.A1(new_n873_), .A2(new_n601_), .A3(new_n360_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT127), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n885_), .A2(new_n613_), .A3(new_n621_), .A4(new_n545_), .ZN(new_n890_));
  INV_X1    g689(.A(G183gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n873_), .B2(new_n838_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n579_), .A2(new_n361_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n873_), .B2(new_n894_), .ZN(G1351gat));
  NOR2_X1   g694(.A1(new_n544_), .A2(new_n468_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n851_), .A2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G197gat), .B1(new_n897_), .B2(new_n338_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n851_), .A2(new_n896_), .ZN(new_n899_));
  INV_X1    g698(.A(G197gat), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n899_), .A2(new_n900_), .A3(new_n739_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n898_), .A2(new_n901_), .ZN(G1352gat));
  OR3_X1    g701(.A1(new_n899_), .A2(G204gat), .A3(new_n305_), .ZN(new_n903_));
  OAI21_X1  g702(.A(G204gat), .B1(new_n899_), .B2(new_n305_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1353gat));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(new_n899_), .B2(new_n601_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT63), .B(G211gat), .Z(new_n908_));
  NAND4_X1  g707(.A1(new_n851_), .A2(new_n613_), .A3(new_n896_), .A4(new_n908_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1354gat));
  OAI21_X1  g709(.A(G218gat), .B1(new_n899_), .B2(new_n838_), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n612_), .A2(G218gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n899_), .B2(new_n912_), .ZN(G1355gat));
endmodule


