//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202_));
  AND2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  AOI22_X1  g008(.A1(new_n203_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n207_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n208_), .B(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT85), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n216_), .A2(G141gat), .A3(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT85), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT2), .ZN(new_n219_));
  AOI22_X1  g018(.A1(new_n216_), .A2(new_n219_), .B1(G141gat), .B2(G148gat), .ZN(new_n220_));
  OR3_X1    g019(.A1(new_n214_), .A2(new_n217_), .A3(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n212_), .B1(new_n221_), .B2(new_n205_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G22gat), .B(G50gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n222_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  NOR3_X1   g025(.A1(new_n214_), .A2(new_n217_), .A3(new_n220_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n205_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n211_), .B(new_n223_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(new_n224_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n226_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n231_), .B1(new_n226_), .B2(new_n230_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n202_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n226_), .A2(new_n230_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n231_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(KEYINPUT87), .A3(new_n232_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n235_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G211gat), .B(G218gat), .Z(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G204gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT88), .B1(new_n243_), .B2(G197gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT88), .ZN(new_n245_));
  INV_X1    g044(.A(G197gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(G204gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(G197gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n242_), .B1(new_n250_), .B2(KEYINPUT89), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT21), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n244_), .A2(new_n247_), .B1(G197gat), .B2(new_n243_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT89), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n252_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n246_), .A2(G204gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n252_), .B1(new_n258_), .B2(new_n249_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n259_), .A2(new_n241_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT90), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n262_), .B(KEYINPUT90), .C1(new_n222_), .C2(new_n223_), .ZN(new_n266_));
  INV_X1    g065(.A(G228gat), .ZN(new_n267_));
  INV_X1    g066(.A(G233gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n265_), .A2(new_n266_), .A3(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G78gat), .B(G106gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT91), .Z(new_n272_));
  OAI211_X1 g071(.A(new_n263_), .B(new_n264_), .C1(new_n267_), .C2(new_n268_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n270_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n272_), .B1(new_n270_), .B2(new_n273_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n240_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n270_), .A2(new_n273_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n272_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n233_), .A2(new_n234_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n270_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n276_), .A2(new_n282_), .A3(KEYINPUT92), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT92), .B1(new_n276_), .B2(new_n282_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT23), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(G183gat), .A3(G190gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT82), .B(G176gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT22), .B(G169gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G169gat), .ZN(new_n296_));
  INV_X1    g095(.A(G176gat), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n292_), .B(new_n295_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G190gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT24), .B1(new_n296_), .B2(new_n297_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT81), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT24), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n287_), .A2(new_n289_), .B1(new_n306_), .B2(new_n304_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(G169gat), .B2(G176gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT81), .ZN(new_n309_));
  INV_X1    g108(.A(new_n304_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n302_), .A2(new_n305_), .A3(new_n307_), .A4(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n285_), .B1(new_n298_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n298_), .A2(new_n312_), .A3(new_n285_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G71gat), .B(G99gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G227gat), .A2(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n314_), .A2(new_n315_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n315_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n318_), .B1(new_n321_), .B2(new_n313_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G15gat), .B(G43gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n320_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(KEYINPUT83), .A3(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G127gat), .B(G134gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G113gat), .ZN(new_n330_));
  INV_X1    g129(.A(G120gat), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n331_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT31), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n328_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT84), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT83), .ZN(new_n338_));
  INV_X1    g137(.A(new_n327_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n324_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(new_n328_), .A3(new_n335_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n336_), .A2(new_n337_), .A3(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n337_), .B1(new_n336_), .B2(new_n342_), .ZN(new_n344_));
  OAI22_X1  g143(.A1(new_n283_), .A2(new_n284_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT92), .ZN(new_n346_));
  INV_X1    g145(.A(new_n281_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n280_), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n347_), .A2(new_n275_), .A3(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n270_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n279_), .A2(new_n350_), .B1(new_n239_), .B2(new_n235_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n346_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n276_), .A2(new_n282_), .A3(KEYINPUT92), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n336_), .A2(new_n342_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n345_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n298_), .A2(new_n312_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT20), .B1(new_n262_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT93), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n294_), .B(KEYINPUT96), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n360_), .A2(new_n293_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n292_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n303_), .A2(KEYINPUT94), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n310_), .B1(new_n303_), .B2(KEYINPUT94), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n302_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n307_), .B(KEYINPUT95), .ZN(new_n366_));
  OAI22_X1  g165(.A1(new_n361_), .A2(new_n362_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n262_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT93), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n369_), .B(KEYINPUT20), .C1(new_n262_), .C2(new_n357_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n359_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT19), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n251_), .A2(new_n255_), .B1(new_n260_), .B2(new_n257_), .ZN(new_n375_));
  OAI221_X1 g174(.A(new_n375_), .B1(new_n365_), .B2(new_n366_), .C1(new_n362_), .C2(new_n361_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n373_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT20), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n262_), .B2(new_n357_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n376_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n374_), .A2(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G8gat), .B(G36gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  NOR2_X1   g186(.A1(new_n382_), .A2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n380_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n387_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT98), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n382_), .A2(KEYINPUT98), .A3(new_n387_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n392_), .A2(KEYINPUT27), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n376_), .A2(new_n379_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n373_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n396_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n397_), .A2(new_n387_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT27), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n388_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n394_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n222_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n334_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n222_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n403_), .A2(KEYINPUT4), .A3(new_n404_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n402_), .A2(new_n334_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n406_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT0), .B(G57gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(G85gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(G1gat), .B(G29gat), .Z(new_n415_));
  XOR2_X1   g214(.A(new_n414_), .B(new_n415_), .Z(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  OR3_X1    g216(.A1(new_n408_), .A2(new_n412_), .A3(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n417_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n356_), .A2(new_n401_), .A3(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n419_), .B(KEYINPUT33), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n409_), .A2(new_n406_), .A3(new_n411_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT99), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n405_), .A2(new_n407_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n416_), .A3(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n423_), .B(new_n427_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n390_), .A2(KEYINPUT32), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n397_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT100), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n382_), .A2(new_n429_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n420_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n283_), .A2(new_n284_), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n343_), .A2(new_n344_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n422_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT67), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT66), .ZN(new_n440_));
  INV_X1    g239(.A(G99gat), .ZN(new_n441_));
  INV_X1    g240(.A(G106gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT7), .ZN(new_n444_));
  AND3_X1   g243(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT7), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n440_), .A2(new_n448_), .A3(new_n441_), .A4(new_n442_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n444_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(G92gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G85gat), .ZN(new_n452_));
  INV_X1    g251(.A(G85gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G92gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT8), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT8), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n450_), .A2(new_n458_), .A3(new_n455_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT65), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT9), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(G85gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n453_), .A2(KEYINPUT65), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n451_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n462_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G99gat), .A2(G106gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n465_), .A2(new_n466_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n441_), .A2(KEYINPUT10), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT10), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G99gat), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n473_), .A2(new_n475_), .A3(KEYINPUT64), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT64), .B1(new_n473_), .B2(new_n475_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n442_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n472_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n439_), .B1(new_n460_), .B2(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n450_), .A2(new_n458_), .A3(new_n455_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n458_), .B1(new_n450_), .B2(new_n455_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n439_), .B(new_n479_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G57gat), .B(G64gat), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n485_), .A2(KEYINPUT11), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(KEYINPUT11), .ZN(new_n487_));
  XOR2_X1   g286(.A(G71gat), .B(G78gat), .Z(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n487_), .A2(new_n488_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OR4_X1    g290(.A1(KEYINPUT68), .A2(new_n480_), .A3(new_n484_), .A4(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n491_), .B1(new_n480_), .B2(new_n484_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n479_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT67), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n489_), .A2(new_n490_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n483_), .A3(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(KEYINPUT68), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G230gat), .A2(G233gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n492_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n481_), .A2(new_n482_), .A3(KEYINPUT69), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT69), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n479_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n496_), .A2(KEYINPUT12), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n503_), .A2(new_n499_), .A3(new_n510_), .A4(new_n493_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n501_), .A2(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G120gat), .B(G148gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G176gat), .B(G204gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n512_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n501_), .A2(new_n511_), .A3(new_n517_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT13), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n519_), .B(new_n520_), .C1(KEYINPUT72), .C2(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n519_), .A2(new_n520_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n522_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(G1gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT75), .B(G8gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT14), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n526_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT14), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n531_), .A3(new_n526_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  OR3_X1    g332(.A1(new_n530_), .A2(G8gat), .A3(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(G8gat), .B1(new_n530_), .B2(new_n533_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G29gat), .B(G36gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(G43gat), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G50gat), .ZN(new_n540_));
  INV_X1    g339(.A(G50gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT78), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n536_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n534_), .A2(new_n535_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT78), .B1(new_n547_), .B2(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT15), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n543_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n540_), .A2(new_n542_), .A3(KEYINPUT15), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n547_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n549_), .A2(new_n550_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n547_), .A2(new_n543_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n550_), .B1(new_n549_), .B2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT79), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G113gat), .B(G141gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(new_n296_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(new_n246_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT80), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n559_), .A2(new_n564_), .ZN(new_n565_));
  OAI211_X1 g364(.A(KEYINPUT79), .B(new_n563_), .C1(new_n556_), .C2(new_n558_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n525_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT17), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n491_), .B(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(new_n536_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n536_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G183gat), .B(G211gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  AND4_X1   g379(.A1(new_n570_), .A2(new_n574_), .A3(new_n575_), .A4(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n570_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n575_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(new_n573_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT77), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n583_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  OAI211_X1 g386(.A(KEYINPUT77), .B(new_n582_), .C1(new_n584_), .C2(new_n573_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n581_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n569_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT34), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n543_), .B1(new_n495_), .B2(new_n483_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT73), .ZN(new_n594_));
  OAI211_X1 g393(.A(KEYINPUT35), .B(new_n592_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n554_), .A2(new_n507_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n592_), .A2(KEYINPUT35), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n595_), .A2(new_n598_), .A3(new_n597_), .A4(new_n599_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(G134gat), .ZN(new_n605_));
  INV_X1    g404(.A(G162gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(KEYINPUT36), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n603_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n601_), .A2(new_n609_), .A3(new_n602_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n608_), .A2(KEYINPUT36), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(KEYINPUT74), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT37), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n615_), .A2(new_n617_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n438_), .A2(new_n590_), .A3(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT101), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n526_), .A3(new_n420_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT38), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n438_), .A2(new_n590_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n615_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G1gat), .B1(new_n628_), .B2(new_n421_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n623_), .A2(new_n624_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n625_), .A2(new_n629_), .A3(new_n630_), .ZN(G1324gat));
  OAI21_X1  g430(.A(G8gat), .B1(new_n628_), .B2(new_n401_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT39), .ZN(new_n633_));
  INV_X1    g432(.A(new_n401_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n622_), .A2(new_n527_), .A3(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(KEYINPUT102), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(KEYINPUT102), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n633_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g438(.A(new_n436_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n627_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G15gat), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n642_), .A2(KEYINPUT103), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(KEYINPUT103), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT41), .ZN(new_n645_));
  OR3_X1    g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n645_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n647_));
  INV_X1    g446(.A(G15gat), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n622_), .A2(new_n648_), .A3(new_n640_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n646_), .A2(new_n647_), .A3(new_n649_), .ZN(G1326gat));
  INV_X1    g449(.A(G22gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n435_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n627_), .B2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT42), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n622_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1327gat));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n618_), .A2(new_n619_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n438_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n438_), .A2(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT43), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n438_), .A2(KEYINPUT104), .A3(new_n658_), .A4(new_n657_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n661_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n589_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n569_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n665_), .A2(KEYINPUT44), .A3(new_n667_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(new_n420_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G29gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n615_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n422_), .B2(new_n437_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(new_n667_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n421_), .A2(G29gat), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT105), .Z(new_n679_));
  OAI21_X1  g478(.A(new_n673_), .B1(new_n677_), .B2(new_n679_), .ZN(G1328gat));
  INV_X1    g479(.A(G36gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n676_), .A2(new_n681_), .A3(new_n634_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT45), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n670_), .A2(new_n634_), .A3(new_n671_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n684_), .B2(new_n681_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT46), .Z(G1329gat));
  NAND2_X1  g485(.A1(new_n670_), .A2(new_n354_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n671_), .A2(G43gat), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n677_), .A2(new_n436_), .ZN(new_n689_));
  OAI22_X1  g488(.A1(new_n687_), .A2(new_n688_), .B1(G43gat), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g490(.A1(new_n676_), .A2(new_n541_), .A3(new_n652_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n670_), .A2(new_n652_), .A3(new_n671_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(G50gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n693_), .B2(G50gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n692_), .B1(new_n696_), .B2(new_n697_), .ZN(G1331gat));
  INV_X1    g497(.A(new_n525_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n438_), .A2(new_n699_), .A3(new_n567_), .A4(new_n666_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(new_n658_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT107), .ZN(new_n702_));
  AOI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n420_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n700_), .A2(new_n421_), .A3(new_n615_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(G57gat), .B2(new_n704_), .ZN(G1332gat));
  INV_X1    g504(.A(G64gat), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n700_), .A2(new_n615_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(new_n634_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT108), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT48), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n702_), .A2(new_n706_), .A3(new_n634_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1333gat));
  INV_X1    g511(.A(G71gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n707_), .B2(new_n640_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT49), .Z(new_n715_));
  NAND3_X1  g514(.A1(new_n702_), .A2(new_n713_), .A3(new_n640_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1334gat));
  INV_X1    g516(.A(G78gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n707_), .B2(new_n652_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT50), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n702_), .A2(new_n718_), .A3(new_n652_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1335gat));
  NOR3_X1   g521(.A1(new_n525_), .A2(new_n568_), .A3(new_n666_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n675_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G85gat), .B1(new_n724_), .B2(new_n420_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n665_), .A2(new_n723_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n461_), .A2(G85gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n421_), .B1(new_n464_), .B2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n725_), .B1(new_n727_), .B2(new_n729_), .ZN(G1336gat));
  NOR3_X1   g529(.A1(new_n726_), .A2(new_n451_), .A3(new_n401_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G92gat), .B1(new_n724_), .B2(new_n634_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT109), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1337gat));
  OAI21_X1  g533(.A(G99gat), .B1(new_n726_), .B2(new_n436_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n724_), .B(new_n354_), .C1(new_n477_), .C2(new_n476_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(KEYINPUT110), .A3(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g537(.A1(new_n665_), .A2(new_n652_), .A3(new_n723_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n665_), .A2(KEYINPUT111), .A3(new_n652_), .A4(new_n723_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(G106gat), .A3(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT52), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n741_), .A2(new_n745_), .A3(G106gat), .A4(new_n742_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n724_), .A2(new_n442_), .A3(new_n652_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT53), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n747_), .A2(new_n751_), .A3(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1339gat));
  NOR3_X1   g552(.A1(new_n634_), .A2(new_n421_), .A3(new_n355_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT118), .Z(new_n755_));
  NAND2_X1  g554(.A1(new_n549_), .A2(new_n555_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n562_), .B1(new_n756_), .B2(new_n550_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n758_));
  AOI22_X1  g557(.A1(new_n549_), .A2(new_n557_), .B1(G229gat), .B2(G233gat), .ZN(new_n759_));
  OR3_X1    g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  OR3_X1    g559(.A1(new_n556_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n758_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n760_), .A2(new_n520_), .A3(new_n761_), .A4(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT69), .B1(new_n481_), .B2(new_n482_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n457_), .A2(new_n505_), .A3(new_n459_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n508_), .B1(new_n767_), .B2(new_n479_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n496_), .B1(new_n495_), .B2(new_n483_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AOI211_X1 g569(.A(new_n764_), .B(new_n499_), .C1(new_n770_), .C2(new_n503_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n503_), .A2(new_n510_), .A3(new_n493_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT114), .B1(new_n772_), .B2(new_n500_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n511_), .A2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n770_), .A2(KEYINPUT55), .A3(new_n499_), .A4(new_n503_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT115), .B1(new_n774_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n772_), .A2(new_n500_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n764_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n772_), .A2(KEYINPUT114), .A3(new_n500_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n776_), .A2(new_n777_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n779_), .A2(new_n786_), .A3(KEYINPUT56), .A4(new_n518_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n763_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n779_), .A2(new_n518_), .A3(new_n786_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(KEYINPUT117), .A3(new_n787_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n790_), .A2(KEYINPUT58), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT58), .B1(new_n790_), .B2(new_n794_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n620_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n568_), .A2(new_n520_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n793_), .B2(new_n787_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n760_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(new_n523_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n674_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT57), .B(new_n674_), .C1(new_n799_), .C2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n589_), .B1(new_n797_), .B2(new_n806_), .ZN(new_n807_));
  AOI211_X1 g606(.A(KEYINPUT112), .B(new_n589_), .C1(new_n565_), .C2(new_n566_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n567_), .B2(new_n666_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(new_n525_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n813_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT54), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n812_), .A2(new_n813_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n814_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n755_), .B1(new_n807_), .B2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(G113gat), .B1(new_n821_), .B2(new_n568_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT59), .B1(new_n821_), .B2(KEYINPUT119), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n793_), .A2(KEYINPUT117), .A3(new_n787_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n763_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n787_), .B2(KEYINPUT117), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n825_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n790_), .A2(new_n794_), .A3(KEYINPUT58), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n658_), .A3(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n819_), .B1(new_n832_), .B2(new_n589_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT59), .ZN(new_n835_));
  NOR4_X1   g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .A4(new_n755_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n567_), .B1(new_n824_), .B2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n822_), .B1(new_n838_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g638(.A(new_n331_), .B1(new_n525_), .B2(KEYINPUT60), .ZN(new_n840_));
  XOR2_X1   g639(.A(new_n840_), .B(KEYINPUT120), .Z(new_n841_));
  OAI211_X1 g640(.A(new_n821_), .B(new_n841_), .C1(KEYINPUT60), .C2(new_n331_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n525_), .B1(new_n824_), .B2(new_n837_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n331_), .ZN(G1341gat));
  AOI21_X1  g643(.A(G127gat), .B1(new_n821_), .B2(new_n666_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT121), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n589_), .B1(new_n824_), .B2(new_n837_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(G127gat), .ZN(G1342gat));
  OAI211_X1 g647(.A(G134gat), .B(new_n658_), .C1(new_n823_), .C2(new_n836_), .ZN(new_n849_));
  INV_X1    g648(.A(G134gat), .ZN(new_n850_));
  INV_X1    g649(.A(new_n821_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n674_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n849_), .A2(KEYINPUT122), .A3(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1343gat));
  NOR2_X1   g656(.A1(new_n833_), .A2(new_n345_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n634_), .A2(new_n421_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n568_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n699_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g664(.A1(new_n860_), .A2(new_n589_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT61), .B(G155gat), .Z(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1346gat));
  NOR3_X1   g667(.A1(new_n860_), .A2(new_n606_), .A3(new_n620_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n861_), .A2(new_n615_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n606_), .B2(new_n870_), .ZN(G1347gat));
  INV_X1    g670(.A(KEYINPUT62), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n401_), .A2(new_n420_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n640_), .ZN(new_n874_));
  NOR4_X1   g673(.A1(new_n833_), .A2(new_n567_), .A3(new_n652_), .A4(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n872_), .B1(new_n875_), .B2(new_n296_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n833_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n874_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n877_), .A2(new_n568_), .A3(new_n435_), .A4(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n875_), .A2(new_n360_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n876_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT123), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n876_), .A2(new_n880_), .A3(new_n884_), .A4(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1348gat));
  NOR3_X1   g685(.A1(new_n833_), .A2(new_n652_), .A3(new_n874_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n699_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n297_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(new_n293_), .B2(new_n888_), .ZN(G1349gat));
  INV_X1    g689(.A(new_n887_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n589_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n892_), .A2(KEYINPUT124), .A3(G183gat), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n301_), .B1(new_n894_), .B2(new_n300_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n892_), .B2(new_n895_), .ZN(G1350gat));
  OAI21_X1  g695(.A(G190gat), .B1(new_n891_), .B2(new_n620_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n887_), .A2(new_n615_), .A3(new_n299_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1351gat));
  AND2_X1   g698(.A1(new_n858_), .A2(new_n873_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n568_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n699_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g703(.A(KEYINPUT63), .ZN(new_n905_));
  INV_X1    g704(.A(G211gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n666_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT125), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n907_), .A2(KEYINPUT125), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n900_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n905_), .A2(new_n906_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1354gat));
  NAND3_X1  g711(.A1(new_n858_), .A2(new_n615_), .A3(new_n873_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n913_), .A2(KEYINPUT126), .ZN(new_n914_));
  INV_X1    g713(.A(G218gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(KEYINPUT126), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n658_), .A2(G218gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT127), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n900_), .A2(new_n919_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n917_), .A2(new_n920_), .ZN(G1355gat));
endmodule


