//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n956_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT74), .B(G8gat), .ZN(new_n205_));
  INV_X1    g004(.A(G1gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT75), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n208_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G1gat), .B(G8gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n211_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n207_), .A2(new_n209_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT75), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n213_), .B1(new_n217_), .B2(new_n210_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n204_), .B1(new_n215_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G229gat), .A2(G233gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n215_), .A2(new_n218_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n219_), .B(new_n220_), .C1(new_n222_), .C2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n218_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n204_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n217_), .A2(new_n210_), .A3(new_n213_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(new_n219_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n220_), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT79), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT79), .ZN(new_n233_));
  AOI211_X1 g032(.A(new_n233_), .B(new_n220_), .C1(new_n229_), .C2(new_n219_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n225_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT82), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT80), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G169gat), .B(G197gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT81), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n235_), .A2(new_n236_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n240_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n225_), .B(new_n243_), .C1(new_n232_), .C2(new_n234_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n236_), .B1(new_n235_), .B2(new_n241_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT83), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n235_), .A2(new_n241_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT82), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT83), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(new_n244_), .A4(new_n242_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT24), .ZN(new_n253_));
  INV_X1    g052(.A(G169gat), .ZN(new_n254_));
  INV_X1    g053(.A(G176gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT23), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n256_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT85), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT85), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n256_), .A2(new_n259_), .A3(new_n263_), .A4(new_n260_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n254_), .A2(new_n255_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(KEYINPUT24), .A3(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G190gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT84), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT25), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(G183gat), .ZN(new_n271_));
  INV_X1    g070(.A(G183gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT25), .B1(new_n272_), .B2(KEYINPUT84), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n268_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n262_), .A2(new_n264_), .A3(new_n267_), .A4(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n259_), .A2(new_n277_), .A3(new_n260_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT22), .ZN(new_n279_));
  OAI21_X1  g078(.A(G169gat), .B1(new_n279_), .B2(KEYINPUT86), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n254_), .A2(KEYINPUT22), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n280_), .B1(KEYINPUT86), .B2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(KEYINPUT87), .B(G176gat), .Z(new_n283_));
  OAI211_X1 g082(.A(new_n278_), .B(new_n266_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n275_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G227gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(G15gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n285_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT31), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G71gat), .B(G99gat), .ZN(new_n291_));
  INV_X1    g090(.A(G43gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT88), .B(KEYINPUT30), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n288_), .A2(new_n289_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n290_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n295_), .B1(new_n290_), .B2(new_n296_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT90), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n290_), .A2(new_n296_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n295_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT90), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n290_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G127gat), .B(G134gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT89), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT89), .ZN(new_n308_));
  INV_X1    g107(.A(G127gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n309_), .A2(G134gat), .ZN(new_n310_));
  INV_X1    g109(.A(G134gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(G127gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n308_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G113gat), .B(G120gat), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n307_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n314_), .B1(new_n307_), .B2(new_n313_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n299_), .A2(new_n305_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n299_), .B2(new_n305_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(G197gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G204gat), .ZN(new_n323_));
  INV_X1    g122(.A(G204gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G197gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT21), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n323_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G218gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(G211gat), .ZN(new_n329_));
  INV_X1    g128(.A(G211gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(G218gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n323_), .A2(new_n325_), .A3(KEYINPUT96), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT21), .B1(new_n323_), .B2(KEYINPUT96), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n327_), .B(new_n333_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G197gat), .B(G204gat), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n337_), .A2(new_n326_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n332_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n341_));
  INV_X1    g140(.A(G141gat), .ZN(new_n342_));
  INV_X1    g141(.A(G148gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G141gat), .A2(G148gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n344_), .A2(new_n347_), .A3(new_n348_), .A4(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  OR3_X1    g150(.A1(KEYINPUT91), .A2(G155gat), .A3(G162gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT91), .B1(G155gat), .B2(G162gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT92), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(G155gat), .B2(G162gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n356_), .A2(KEYINPUT92), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n352_), .B(new_n353_), .C1(new_n355_), .C2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT93), .B1(new_n351_), .B2(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n352_), .A2(new_n353_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(KEYINPUT92), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n354_), .A2(G155gat), .A3(G162gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT93), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n360_), .A2(new_n350_), .A3(new_n363_), .A4(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(KEYINPUT1), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n361_), .A2(new_n362_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n360_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G141gat), .B(G148gat), .Z(new_n370_));
  AOI22_X1  g169(.A1(new_n359_), .A2(new_n365_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  OAI211_X1 g171(.A(KEYINPUT97), .B(new_n340_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT94), .ZN(new_n374_));
  OAI21_X1  g173(.A(G228gat), .B1(new_n374_), .B2(G233gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n374_), .B2(G233gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G22gat), .B(G50gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT28), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n371_), .A2(new_n379_), .A3(new_n372_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n378_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n382_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n378_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n380_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n377_), .B1(new_n383_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G106gat), .ZN(new_n389_));
  OAI211_X1 g188(.A(KEYINPUT95), .B(new_n340_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT97), .ZN(new_n391_));
  INV_X1    g190(.A(G78gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n392_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n389_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n395_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n397_), .A2(G106gat), .A3(new_n393_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n383_), .A2(new_n386_), .A3(new_n377_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n388_), .A2(new_n396_), .A3(new_n398_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT104), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n359_), .A2(new_n365_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n369_), .A2(new_n370_), .ZN(new_n404_));
  AND4_X1   g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .A4(new_n317_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n317_), .B1(new_n371_), .B2(new_n402_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n401_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n403_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n317_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n371_), .A2(new_n402_), .A3(new_n317_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n408_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n401_), .B(KEYINPUT105), .Z(new_n414_));
  NAND2_X1  g213(.A1(new_n317_), .A2(new_n408_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n414_), .B1(new_n415_), .B2(new_n371_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n407_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G1gat), .B(G29gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(G85gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT0), .B(G57gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n407_), .B(new_n421_), .C1(new_n413_), .C2(new_n416_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n394_), .A2(new_n389_), .A3(new_n395_), .ZN(new_n427_));
  AOI21_X1  g226(.A(G106gat), .B1(new_n397_), .B2(new_n393_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n383_), .A2(new_n386_), .A3(new_n377_), .ZN(new_n429_));
  OAI22_X1  g228(.A1(new_n427_), .A2(new_n428_), .B1(new_n429_), .B2(new_n387_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT102), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n285_), .A2(KEYINPUT100), .A3(new_n340_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT100), .B1(new_n285_), .B2(new_n340_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n276_), .A2(KEYINPUT26), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT26), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G190gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n270_), .A2(G183gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n272_), .A2(KEYINPUT25), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n435_), .A2(new_n437_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT98), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n253_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(KEYINPUT98), .A2(KEYINPUT24), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n265_), .A2(new_n442_), .A3(new_n266_), .A4(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n260_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G169gat), .A2(G176gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n443_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(KEYINPUT98), .A2(KEYINPUT24), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n440_), .A2(new_n444_), .A3(new_n447_), .A4(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT99), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n266_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(KEYINPUT99), .A2(G169gat), .A3(G176gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n279_), .A2(G169gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n281_), .A2(new_n457_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n278_), .B(new_n456_), .C1(new_n283_), .C2(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n336_), .A2(new_n452_), .A3(new_n339_), .A4(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT101), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n332_), .B1(new_n326_), .B2(new_n337_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n323_), .A2(new_n325_), .A3(KEYINPUT96), .ZN(new_n463_));
  OR3_X1    g262(.A1(new_n324_), .A2(KEYINPUT96), .A3(G197gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(KEYINPUT21), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n462_), .A2(new_n465_), .B1(new_n332_), .B2(new_n338_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT101), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n466_), .A2(new_n467_), .A3(new_n459_), .A4(new_n452_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G226gat), .A2(G233gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT19), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n461_), .A2(new_n468_), .A3(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n431_), .B1(new_n434_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n285_), .A2(new_n340_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT100), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n285_), .A2(KEYINPUT100), .A3(new_n340_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n461_), .A2(new_n468_), .A3(new_n472_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(KEYINPUT102), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n452_), .A2(new_n459_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n471_), .B1(new_n340_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n466_), .A2(new_n284_), .A3(new_n275_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n470_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G8gat), .B(G36gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT18), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G64gat), .B(G92gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n474_), .A2(new_n481_), .A3(new_n486_), .A4(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n485_), .A2(new_n470_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n479_), .A2(KEYINPUT20), .A3(new_n460_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(new_n470_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n491_), .B(KEYINPUT27), .C1(new_n494_), .C2(new_n490_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n400_), .A2(new_n426_), .A3(new_n430_), .A4(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(KEYINPUT103), .ZN(new_n497_));
  INV_X1    g296(.A(new_n486_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n473_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n498_), .B1(new_n499_), .B2(KEYINPUT102), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT103), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n474_), .A4(new_n490_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n474_), .A2(new_n486_), .A3(new_n481_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n490_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n497_), .A2(new_n502_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT27), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT109), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n506_), .A2(KEYINPUT109), .A3(new_n507_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n496_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n400_), .A2(new_n430_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n497_), .A2(new_n505_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT106), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT33), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n424_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n424_), .A2(new_n515_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n411_), .A2(new_n412_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT107), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT107), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n411_), .A2(new_n521_), .A3(new_n412_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n414_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n519_), .A2(KEYINPUT4), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n415_), .A2(new_n371_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(G225gat), .B2(G233gat), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n421_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n518_), .A2(KEYINPUT33), .B1(new_n523_), .B2(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n514_), .A2(new_n502_), .A3(new_n517_), .A4(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n490_), .A2(KEYINPUT32), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n494_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n530_), .B(KEYINPUT108), .Z(new_n532_));
  OAI211_X1 g331(.A(new_n531_), .B(new_n425_), .C1(new_n503_), .C2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n513_), .B1(new_n529_), .B2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n321_), .B1(new_n512_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n510_), .A2(new_n511_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n318_), .A2(new_n319_), .A3(new_n425_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n400_), .A2(new_n430_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .A4(new_n495_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n252_), .B1(new_n535_), .B2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G127gat), .B(G155gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(G183gat), .B(G211gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT78), .B1(new_n545_), .B2(KEYINPUT17), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  XNOR2_X1  g347(.A(G71gat), .B(G78gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(G57gat), .B(G64gat), .Z(new_n550_));
  INV_X1    g349(.A(KEYINPUT11), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n549_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT67), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G71gat), .B(G78gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(G57gat), .B(G64gat), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n555_), .B1(KEYINPUT11), .B2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n557_), .A2(KEYINPUT67), .ZN(new_n558_));
  OAI22_X1  g357(.A1(new_n554_), .A2(new_n558_), .B1(new_n551_), .B2(new_n550_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n552_), .A2(new_n553_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(KEYINPUT67), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n550_), .A2(new_n551_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT76), .Z(new_n565_));
  NAND2_X1  g364(.A1(new_n548_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n548_), .A2(new_n565_), .ZN(new_n568_));
  OR3_X1    g367(.A1(new_n567_), .A2(new_n221_), .A3(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n221_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n545_), .A2(KEYINPUT17), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT8), .ZN(new_n573_));
  XOR2_X1   g372(.A(G85gat), .B(G92gat), .Z(new_n574_));
  NOR2_X1   g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT7), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT6), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n574_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(KEYINPUT9), .B2(new_n574_), .ZN(new_n582_));
  XOR2_X1   g381(.A(KEYINPUT10), .B(G99gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT65), .B(G85gat), .ZN(new_n584_));
  INV_X1    g383(.A(G92gat), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(KEYINPUT9), .ZN(new_n586_));
  AOI22_X1  g385(.A1(new_n583_), .A2(new_n389_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n573_), .A2(new_n581_), .B1(new_n582_), .B2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n575_), .B(KEYINPUT7), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT66), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n577_), .A2(KEYINPUT66), .ZN(new_n592_));
  INV_X1    g391(.A(new_n580_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n574_), .A2(KEYINPUT8), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n588_), .A2(new_n597_), .A3(new_n204_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT70), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT70), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n588_), .A2(new_n597_), .A3(new_n600_), .A4(new_n204_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n588_), .A2(new_n597_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT35), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n223_), .A2(new_n603_), .B1(new_n604_), .B2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n604_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n602_), .A2(new_n608_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n610_), .B1(new_n602_), .B2(new_n608_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT72), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n602_), .A2(new_n608_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n609_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT72), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(new_n617_), .A3(new_n611_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT36), .Z(new_n622_));
  NAND3_X1  g421(.A1(new_n614_), .A2(new_n618_), .A3(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(KEYINPUT36), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n616_), .A2(new_n624_), .A3(new_n611_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n623_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n625_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n622_), .B(KEYINPUT71), .Z(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n616_), .B2(new_n611_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT37), .B1(new_n628_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n563_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n562_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n581_), .A2(new_n573_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n574_), .A2(KEYINPUT9), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n587_), .A2(new_n593_), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n580_), .B1(new_n577_), .B2(KEYINPUT66), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n595_), .B1(new_n639_), .B2(new_n591_), .ZN(new_n640_));
  OAI22_X1  g439(.A1(new_n633_), .A2(new_n634_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n559_), .A2(new_n588_), .A3(new_n597_), .A4(new_n563_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT64), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT68), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n641_), .A2(new_n642_), .A3(KEYINPUT12), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT12), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n564_), .A2(new_n603_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n645_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n649_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT5), .ZN(new_n657_));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n657_), .B(new_n658_), .Z(new_n659_));
  NAND2_X1  g458(.A1(new_n655_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n659_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n649_), .A2(new_n654_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT13), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(KEYINPUT13), .A3(new_n662_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n572_), .A2(new_n632_), .A3(new_n665_), .A4(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n540_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n206_), .A3(new_n425_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(KEYINPUT38), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT110), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n623_), .A2(new_n625_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n535_), .B2(new_n539_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n665_), .A2(new_n666_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n252_), .A2(new_n678_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n677_), .A2(new_n572_), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n206_), .B1(new_n680_), .B2(new_n425_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n672_), .B2(KEYINPUT38), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n674_), .A2(new_n682_), .ZN(G1324gat));
  NAND2_X1  g482(.A1(new_n536_), .A2(new_n495_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n670_), .A2(new_n205_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n680_), .A2(new_n684_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G8gat), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(KEYINPUT39), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(KEYINPUT39), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(G1325gat));
  NAND2_X1  g491(.A1(new_n680_), .A2(new_n320_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G15gat), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT41), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n669_), .A2(G15gat), .A3(new_n321_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1326gat));
  NAND2_X1  g496(.A1(new_n680_), .A2(new_n513_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G22gat), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(KEYINPUT42), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(KEYINPUT42), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n538_), .A2(G22gat), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT111), .ZN(new_n703_));
  OAI22_X1  g502(.A1(new_n700_), .A2(new_n701_), .B1(new_n669_), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT112), .ZN(G1327gat));
  NOR3_X1   g504(.A1(new_n678_), .A2(new_n675_), .A3(new_n572_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n540_), .A2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G29gat), .B1(new_n707_), .B2(new_n425_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n627_), .A2(KEYINPUT113), .A3(new_n631_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT43), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n535_), .A2(new_n539_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n632_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  AOI211_X1 g514(.A(new_n632_), .B(new_n711_), .C1(new_n535_), .C2(new_n539_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n709_), .B(new_n679_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT44), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n425_), .A2(G29gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n708_), .B1(new_n718_), .B2(new_n719_), .ZN(G1328gat));
  NOR2_X1   g519(.A1(KEYINPUT114), .A2(KEYINPUT46), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(G36gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n707_), .A2(new_n723_), .A3(new_n684_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT45), .Z(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n718_), .A2(new_n684_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n722_), .B(new_n726_), .C1(new_n727_), .C2(new_n723_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n723_), .B1(new_n718_), .B2(new_n684_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n721_), .B1(new_n729_), .B2(new_n725_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1329gat));
  NAND3_X1  g530(.A1(new_n718_), .A2(G43gat), .A3(new_n320_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n707_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n292_), .B1(new_n733_), .B2(new_n321_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT47), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n732_), .A2(new_n737_), .A3(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1330gat));
  AOI21_X1  g538(.A(G50gat), .B1(new_n707_), .B2(new_n513_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n513_), .A2(G50gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n718_), .B2(new_n741_), .ZN(G1331gat));
  NAND2_X1  g541(.A1(new_n713_), .A2(new_n252_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(KEYINPUT115), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(KEYINPUT115), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n678_), .A2(new_n572_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n746_), .A2(new_n714_), .A3(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(G57gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n425_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n247_), .A2(new_n251_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n747_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n677_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G57gat), .B1(new_n753_), .B2(new_n426_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n750_), .A2(new_n754_), .ZN(G1332gat));
  INV_X1    g554(.A(G64gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n748_), .A2(new_n756_), .A3(new_n684_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n684_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G64gat), .B1(new_n753_), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT48), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n757_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(G1333gat));
  INV_X1    g562(.A(G71gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n748_), .A2(new_n764_), .A3(new_n320_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G71gat), .B1(new_n753_), .B2(new_n321_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT49), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1334gat));
  NAND3_X1  g567(.A1(new_n748_), .A2(new_n392_), .A3(new_n513_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G78gat), .B1(new_n753_), .B2(new_n538_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT50), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1335gat));
  NAND2_X1  g571(.A1(new_n678_), .A2(new_n709_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n746_), .A2(new_n675_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(G85gat), .B1(new_n774_), .B2(new_n425_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n773_), .A2(new_n751_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n496_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n506_), .A2(KEYINPUT109), .A3(new_n507_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT109), .B1(new_n506_), .B2(new_n507_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n528_), .A2(new_n517_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n533_), .B1(new_n782_), .B2(new_n506_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n538_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n320_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n538_), .B(new_n495_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n320_), .A2(new_n426_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n714_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n711_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n713_), .A2(new_n714_), .A3(new_n712_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n777_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n425_), .A2(new_n584_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n775_), .B1(new_n792_), .B2(new_n793_), .ZN(G1336gat));
  NAND3_X1  g593(.A1(new_n774_), .A2(new_n585_), .A3(new_n684_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n792_), .ZN(new_n796_));
  OAI21_X1  g595(.A(G92gat), .B1(new_n796_), .B2(new_n758_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1337gat));
  AND2_X1   g597(.A1(new_n320_), .A2(new_n583_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n792_), .A2(new_n320_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n774_), .A2(new_n799_), .B1(G99gat), .B2(new_n800_), .ZN(new_n801_));
  XOR2_X1   g600(.A(new_n801_), .B(KEYINPUT51), .Z(G1338gat));
  OAI211_X1 g601(.A(new_n513_), .B(new_n776_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n803_));
  OAI21_X1  g602(.A(G106gat), .B1(new_n803_), .B2(KEYINPUT117), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n792_), .B2(new_n513_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT52), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n792_), .A2(new_n805_), .A3(new_n513_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n803_), .A2(KEYINPUT117), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n808_), .A2(new_n809_), .A3(new_n810_), .A4(G106gat), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n807_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n774_), .A2(new_n389_), .A3(new_n513_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT53), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n816_), .A3(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1339gat));
  INV_X1    g617(.A(KEYINPUT121), .ZN(new_n819_));
  XNOR2_X1  g618(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT119), .Z(new_n821_));
  NAND3_X1  g620(.A1(new_n668_), .A2(new_n252_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n821_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n667_), .B2(new_n751_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n646_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n650_), .A2(new_n646_), .A3(new_n652_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(KEYINPUT55), .B2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n653_), .A2(KEYINPUT55), .A3(new_n645_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT56), .B(new_n659_), .C1(new_n829_), .C2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n662_), .B1(new_n832_), .B2(KEYINPUT120), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n828_), .A2(KEYINPUT55), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n654_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n830_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT56), .B1(new_n836_), .B2(new_n659_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n838_), .B(new_n661_), .C1(new_n835_), .C2(new_n830_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n833_), .B1(new_n840_), .B2(KEYINPUT120), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n243_), .B1(new_n230_), .B2(new_n220_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n222_), .A2(new_n224_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n219_), .A2(new_n231_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n244_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n841_), .A2(new_n751_), .B1(new_n663_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n826_), .B1(new_n848_), .B2(new_n676_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n663_), .A2(new_n847_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n659_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n838_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(KEYINPUT120), .A3(new_n832_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n832_), .A2(KEYINPUT120), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n662_), .A3(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n850_), .B1(new_n252_), .B2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(KEYINPUT57), .A3(new_n675_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n847_), .A2(new_n662_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n840_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n714_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n840_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n849_), .A2(new_n857_), .A3(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n825_), .B1(new_n864_), .B2(new_n709_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n320_), .A2(new_n425_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n786_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n865_), .A2(new_n252_), .A3(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n819_), .B1(new_n869_), .B2(G113gat), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n867_), .A2(KEYINPUT122), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n867_), .A2(KEYINPUT122), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n871_), .B1(new_n865_), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT59), .B1(new_n865_), .B2(new_n868_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n875_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n861_), .A2(new_n862_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n856_), .A2(new_n675_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n826_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n572_), .B1(new_n881_), .B2(new_n857_), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT123), .B(new_n878_), .C1(new_n882_), .C2(new_n825_), .ZN(new_n883_));
  INV_X1    g682(.A(G113gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n252_), .A2(new_n884_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n876_), .A2(new_n877_), .A3(new_n883_), .A4(new_n885_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n751_), .B(new_n867_), .C1(new_n882_), .C2(new_n825_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(KEYINPUT121), .A3(new_n884_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n870_), .A2(new_n886_), .A3(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n870_), .A2(new_n886_), .A3(KEYINPUT124), .A4(new_n888_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1340gat));
  AND4_X1   g692(.A1(new_n678_), .A2(new_n876_), .A3(new_n877_), .A4(new_n883_), .ZN(new_n894_));
  INV_X1    g693(.A(G120gat), .ZN(new_n895_));
  INV_X1    g694(.A(new_n865_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n867_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n678_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n895_), .B1(new_n898_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(KEYINPUT60), .B2(new_n895_), .ZN(new_n900_));
  OAI22_X1  g699(.A1(new_n894_), .A2(new_n895_), .B1(new_n897_), .B2(new_n900_), .ZN(G1341gat));
  AND4_X1   g700(.A1(new_n572_), .A2(new_n876_), .A3(new_n877_), .A4(new_n883_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n572_), .A2(new_n309_), .ZN(new_n903_));
  OAI22_X1  g702(.A1(new_n902_), .A2(new_n309_), .B1(new_n897_), .B2(new_n903_), .ZN(G1342gat));
  AND4_X1   g703(.A1(new_n714_), .A2(new_n876_), .A3(new_n877_), .A4(new_n883_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n676_), .A2(new_n311_), .ZN(new_n906_));
  OAI22_X1  g705(.A1(new_n905_), .A2(new_n311_), .B1(new_n897_), .B2(new_n906_), .ZN(G1343gat));
  NAND4_X1  g706(.A1(new_n758_), .A2(new_n513_), .A3(new_n425_), .A4(new_n321_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n865_), .A2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n751_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n678_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g712(.A1(new_n909_), .A2(new_n572_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT61), .B(G155gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1346gat));
  INV_X1    g715(.A(new_n909_), .ZN(new_n917_));
  OR3_X1    g716(.A1(new_n917_), .A2(G162gat), .A3(new_n675_), .ZN(new_n918_));
  OAI21_X1  g717(.A(G162gat), .B1(new_n917_), .B2(new_n632_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1347gat));
  XNOR2_X1  g719(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n758_), .A2(new_n513_), .A3(new_n787_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n896_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n252_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n921_), .B1(new_n924_), .B2(new_n254_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n921_), .ZN(new_n926_));
  OAI211_X1 g725(.A(G169gat), .B(new_n926_), .C1(new_n923_), .C2(new_n252_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n924_), .A2(new_n281_), .A3(new_n457_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n925_), .A2(new_n927_), .A3(new_n928_), .ZN(G1348gat));
  NOR2_X1   g728(.A1(new_n923_), .A2(new_n898_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(new_n283_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n931_), .B1(G176gat), .B2(new_n930_), .ZN(G1349gat));
  NOR2_X1   g731(.A1(new_n923_), .A2(new_n709_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(G183gat), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n438_), .A2(new_n439_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n934_), .B1(new_n935_), .B2(new_n933_), .ZN(G1350gat));
  OAI21_X1  g735(.A(G190gat), .B1(new_n923_), .B2(new_n632_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n676_), .A2(new_n268_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n923_), .B2(new_n938_), .ZN(G1351gat));
  NOR3_X1   g738(.A1(new_n320_), .A2(new_n538_), .A3(new_n425_), .ZN(new_n940_));
  XOR2_X1   g739(.A(new_n940_), .B(KEYINPUT126), .Z(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n684_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n865_), .A2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n751_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n678_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g746(.A1(new_n943_), .A2(new_n572_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n949_));
  AND2_X1   g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n948_), .A2(new_n949_), .A3(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n951_), .B1(new_n948_), .B2(new_n949_), .ZN(G1354gat));
  NAND3_X1  g751(.A1(new_n943_), .A2(new_n328_), .A3(new_n676_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n865_), .A2(new_n632_), .A3(new_n942_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n328_), .B2(new_n954_), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n955_), .B(new_n956_), .ZN(G1355gat));
endmodule


