//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  OAI21_X1  g001(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n208_), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n203_), .B(new_n207_), .C1(new_n209_), .C2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n212_), .A2(KEYINPUT65), .A3(new_n217_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(KEYINPUT8), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n226_), .A2(G85gat), .A3(G92gat), .A4(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n215_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n216_), .ZN(new_n229_));
  OR2_X1    g028(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n206_), .A3(new_n231_), .ZN(new_n232_));
  AND4_X1   g031(.A1(new_n225_), .A2(new_n228_), .A3(new_n229_), .A4(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT65), .B1(new_n212_), .B2(new_n217_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT8), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT12), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n222_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G57gat), .B(G64gat), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n241_));
  XOR2_X1   g040(.A(G71gat), .B(G78gat), .Z(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n241_), .A2(new_n242_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n238_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n237_), .A2(KEYINPUT66), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n249_), .B1(new_n222_), .B2(new_n236_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n222_), .A2(new_n236_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(KEYINPUT12), .A4(new_n245_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n202_), .B1(new_n251_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G120gat), .B(G148gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT5), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G176gat), .B(G204gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n252_), .A2(new_n245_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n202_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n212_), .A2(KEYINPUT65), .A3(new_n217_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n264_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n218_), .A2(new_n219_), .A3(new_n235_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n233_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n263_), .B1(new_n269_), .B2(new_n246_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n256_), .B(new_n261_), .C1(new_n262_), .C2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n248_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(new_n246_), .A3(new_n238_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n263_), .B1(new_n273_), .B2(new_n254_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n270_), .A2(new_n262_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n260_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n271_), .A2(KEYINPUT13), .A3(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT13), .B1(new_n271_), .B2(new_n276_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT67), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT68), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT37), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G190gat), .B(G218gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT71), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G134gat), .B(G162gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G29gat), .B(G36gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G43gat), .B(G50gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n269_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT69), .B(KEYINPUT15), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n289_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n252_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G232gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT34), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n297_), .A2(KEYINPUT35), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n291_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT70), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n291_), .A2(new_n295_), .A3(new_n301_), .A4(new_n298_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n291_), .A2(new_n295_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n297_), .A2(KEYINPUT35), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n298_), .A2(new_n304_), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n300_), .A2(new_n302_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT36), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n286_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n300_), .A2(new_n302_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n303_), .A2(new_n305_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n286_), .A2(new_n307_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n308_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n312_), .B1(new_n308_), .B2(new_n313_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n282_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n308_), .A2(new_n313_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n312_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n308_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(KEYINPUT37), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G231gat), .A2(G233gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n246_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n246_), .A2(new_n324_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT73), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G15gat), .B(G22gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G1gat), .A2(G8gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT14), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G1gat), .B(G8gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n245_), .A2(new_n323_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(new_n325_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n328_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n335_), .B1(new_n328_), .B2(new_n338_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n253_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n341_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(KEYINPUT66), .A3(new_n339_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G127gat), .B(G155gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT16), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G183gat), .B(G211gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT17), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n349_), .B(KEYINPUT74), .Z(new_n350_));
  NAND3_X1  g149(.A1(new_n342_), .A2(new_n344_), .A3(new_n350_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n348_), .A2(KEYINPUT17), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n352_), .B(new_n349_), .C1(new_n340_), .C2(new_n341_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n322_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n281_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT90), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT84), .ZN(new_n358_));
  INV_X1    g157(.A(G197gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(G204gat), .ZN(new_n360_));
  INV_X1    g159(.A(G204gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(KEYINPUT84), .A3(G197gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(G204gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT21), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G211gat), .B(G218gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT85), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n367_), .B1(new_n359_), .B2(G204gat), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n361_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n369_));
  OAI22_X1  g168(.A1(new_n368_), .A2(new_n369_), .B1(new_n359_), .B2(G204gat), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n365_), .B(new_n366_), .C1(new_n370_), .C2(KEYINPUT21), .ZN(new_n371_));
  INV_X1    g170(.A(new_n366_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(KEYINPUT21), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT88), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT83), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(G141gat), .A2(G148gat), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n381_), .A2(KEYINPUT2), .ZN(new_n382_));
  NOR2_X1   g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n381_), .A2(KEYINPUT2), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n382_), .A2(new_n385_), .A3(new_n386_), .A4(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n380_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT1), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n379_), .B(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n378_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n381_), .A2(new_n383_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT29), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT87), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n380_), .A2(new_n388_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399_));
  OR3_X1    g198(.A1(new_n398_), .A2(KEYINPUT87), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n375_), .A2(new_n397_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(G228gat), .ZN(new_n402_));
  INV_X1    g201(.A(G233gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT86), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n374_), .B(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n395_), .B2(KEYINPUT29), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(KEYINPUT89), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n405_), .A2(new_n413_), .A3(new_n409_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G22gat), .B(G50gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT28), .B1(new_n395_), .B2(KEYINPUT29), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n395_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n416_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n419_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(new_n417_), .A3(new_n415_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n414_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n357_), .B1(new_n412_), .B2(new_n425_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n401_), .A2(new_n404_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n423_), .B1(new_n427_), .B2(new_n413_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n410_), .A2(new_n411_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(KEYINPUT90), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n413_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n410_), .A2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n424_), .B1(new_n433_), .B2(new_n414_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT91), .B1(new_n431_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT91), .ZN(new_n437_));
  AOI211_X1 g236(.A(new_n437_), .B(new_n434_), .C1(new_n426_), .C2(new_n430_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G183gat), .A2(G190gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT23), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n441_), .B1(G183gat), .B2(G190gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(G169gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT25), .B(G183gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT26), .B(G190gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(G169gat), .ZN(new_n451_));
  INV_X1    g250(.A(G176gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  OR3_X1    g252(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n448_), .A2(new_n453_), .A3(new_n441_), .A4(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n445_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n439_), .B1(new_n374_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n441_), .A2(new_n454_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT78), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n450_), .B(KEYINPUT76), .C1(new_n451_), .C2(new_n452_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n461_), .A2(new_n448_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT76), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n453_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(KEYINPUT77), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT77), .B1(new_n462_), .B2(new_n464_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n445_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n457_), .B1(new_n468_), .B2(new_n407_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G226gat), .A2(G233gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT19), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n439_), .B1(new_n468_), .B2(new_n407_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n374_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n456_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n471_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n472_), .A2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G8gat), .B(G36gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(G64gat), .B(G92gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n481_), .B(new_n482_), .Z(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n472_), .A2(new_n477_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n483_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n471_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n375_), .A2(new_n456_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n491_), .B1(new_n492_), .B2(new_n473_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n469_), .A2(new_n471_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n486_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n484_), .A2(KEYINPUT27), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n490_), .A2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G127gat), .B(G134gat), .Z(new_n498_));
  XOR2_X1   g297(.A(G113gat), .B(G120gat), .Z(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  NAND2_X1  g299(.A1(new_n395_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n500_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n398_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n503_), .A3(KEYINPUT4), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G225gat), .A2(G233gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT93), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n504_), .B(new_n506_), .C1(KEYINPUT4), .C2(new_n501_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n501_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G1gat), .B(G29gat), .Z(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G85gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n507_), .A2(new_n508_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT96), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n507_), .A2(new_n508_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n513_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n507_), .A2(new_n508_), .A3(KEYINPUT96), .A4(new_n514_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  OAI22_X1  g320(.A1(new_n436_), .A2(new_n438_), .B1(new_n497_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n430_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT90), .B1(new_n428_), .B2(new_n429_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n435_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n437_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n431_), .A2(KEYINPUT91), .A3(new_n435_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n501_), .A2(new_n503_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT95), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT95), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n501_), .A2(new_n503_), .A3(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n506_), .A3(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n504_), .B(new_n505_), .C1(KEYINPUT4), .C2(new_n501_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n532_), .A2(new_n513_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT33), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n515_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n515_), .A2(new_n535_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n536_), .A2(new_n484_), .A3(new_n487_), .A4(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT32), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n478_), .B1(new_n539_), .B2(new_n486_), .ZN(new_n540_));
  OAI211_X1 g339(.A(KEYINPUT32), .B(new_n483_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(new_n521_), .A3(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n526_), .A2(new_n527_), .A3(new_n538_), .A4(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G15gat), .B(G43gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT79), .B(KEYINPUT81), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G227gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT80), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n546_), .B(new_n548_), .Z(new_n549_));
  XNOR2_X1  g348(.A(G71gat), .B(G99gat), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n468_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n468_), .A2(new_n551_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n550_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n554_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n550_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n552_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n549_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT82), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n555_), .A2(new_n558_), .A3(new_n549_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT82), .B1(new_n564_), .B2(new_n559_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n500_), .B(KEYINPUT31), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n563_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n566_), .ZN(new_n568_));
  OAI211_X1 g367(.A(KEYINPUT82), .B(new_n568_), .C1(new_n564_), .C2(new_n559_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n522_), .A2(new_n543_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n521_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n567_), .A2(new_n572_), .A3(new_n569_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n436_), .A2(new_n438_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n497_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n293_), .A2(new_n334_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n335_), .A2(new_n289_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT75), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G229gat), .A2(G233gat), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n334_), .A2(new_n290_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n583_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n582_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(new_n580_), .B2(new_n587_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G113gat), .B(G141gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G169gat), .B(G197gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n591_), .B(new_n592_), .Z(new_n593_));
  NOR2_X1   g392(.A1(new_n590_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n593_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n584_), .B2(new_n589_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT98), .B1(new_n577_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n601_));
  AOI211_X1 g400(.A(new_n601_), .B(new_n597_), .C1(new_n571_), .C2(new_n576_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n356_), .B1(new_n600_), .B2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n572_), .A2(G1gat), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT38), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n609_));
  INV_X1    g408(.A(new_n280_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n609_), .B1(new_n610_), .B2(new_n597_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n354_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n280_), .A2(KEYINPUT100), .A3(new_n598_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n314_), .A2(new_n315_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n571_), .B2(new_n576_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n614_), .A2(KEYINPUT101), .A3(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT101), .B1(new_n614_), .B2(new_n616_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n521_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(G1gat), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n608_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n604_), .A2(KEYINPUT99), .A3(KEYINPUT38), .A4(new_n605_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n624_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .A4(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n625_), .A2(new_n623_), .A3(new_n608_), .A4(new_n620_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT102), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1324gat));
  NAND2_X1  g428(.A1(new_n614_), .A2(new_n616_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G8gat), .B1(new_n630_), .B2(new_n575_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT39), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n575_), .A2(G8gat), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n633_), .B1(new_n604_), .B2(new_n634_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n604_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n632_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n632_), .B(KEYINPUT40), .C1(new_n635_), .C2(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1325gat));
  INV_X1    g440(.A(new_n604_), .ZN(new_n642_));
  OR3_X1    g441(.A1(new_n642_), .A2(G15gat), .A3(new_n570_), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n617_), .A2(new_n618_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n570_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n646_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT41), .B1(new_n646_), .B2(G15gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n643_), .B1(new_n647_), .B2(new_n648_), .ZN(G1326gat));
  OR3_X1    g448(.A1(new_n642_), .A2(G22gat), .A3(new_n574_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n574_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n644_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n652_), .A2(new_n653_), .A3(G22gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n652_), .B2(G22gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n650_), .B1(new_n654_), .B2(new_n655_), .ZN(G1327gat));
  NAND2_X1  g455(.A1(new_n600_), .A2(new_n603_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n615_), .A2(new_n354_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n610_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(G29gat), .B1(new_n661_), .B2(new_n521_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n611_), .A2(new_n354_), .A3(new_n613_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT43), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n577_), .A2(new_n322_), .A3(new_n665_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n664_), .A2(KEYINPUT43), .ZN(new_n667_));
  AOI22_X1  g466(.A1(new_n577_), .A2(new_n322_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n663_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n663_), .B(KEYINPUT44), .C1(new_n666_), .C2(new_n668_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n521_), .A2(G29gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n662_), .B1(new_n673_), .B2(new_n674_), .ZN(G1328gat));
  NAND3_X1  g474(.A1(new_n671_), .A2(new_n497_), .A3(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(G36gat), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT45), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n575_), .A2(G36gat), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n659_), .B(new_n679_), .C1(new_n599_), .C2(new_n602_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(KEYINPUT105), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(KEYINPUT105), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n680_), .A2(KEYINPUT105), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n680_), .A2(KEYINPUT105), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(KEYINPUT45), .A3(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n677_), .A2(new_n683_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(KEYINPUT46), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n689_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n677_), .A2(new_n683_), .A3(new_n686_), .A4(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1329gat));
  NAND4_X1  g492(.A1(new_n671_), .A2(G43gat), .A3(new_n645_), .A4(new_n672_), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT107), .B(G43gat), .Z(new_n695_));
  OAI21_X1  g494(.A(new_n695_), .B1(new_n660_), .B2(new_n570_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g497(.A(G50gat), .B1(new_n661_), .B2(new_n651_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n651_), .A2(G50gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n673_), .B2(new_n700_), .ZN(G1331gat));
  AOI21_X1  g500(.A(new_n598_), .B1(new_n571_), .B2(new_n576_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n702_), .A2(new_n610_), .A3(new_n355_), .ZN(new_n703_));
  INV_X1    g502(.A(G57gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n704_), .A3(new_n521_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n351_), .A2(new_n597_), .A3(new_n353_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n281_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n616_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT108), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(new_n521_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n710_), .B2(new_n704_), .ZN(G1332gat));
  INV_X1    g510(.A(G64gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n703_), .A2(new_n712_), .A3(new_n497_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n709_), .A2(new_n497_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(G64gat), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n714_), .B2(G64gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(G1333gat));
  INV_X1    g517(.A(G71gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n703_), .A2(new_n719_), .A3(new_n645_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT49), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n709_), .A2(new_n645_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(G71gat), .ZN(new_n723_));
  AOI211_X1 g522(.A(KEYINPUT49), .B(new_n719_), .C1(new_n709_), .C2(new_n645_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(G1334gat));
  NOR2_X1   g524(.A1(new_n574_), .A2(G78gat), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT110), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n703_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n709_), .A2(new_n651_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT50), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(G78gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n729_), .B2(G78gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(G1335gat));
  NAND2_X1  g532(.A1(new_n577_), .A2(new_n597_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n734_), .A2(new_n281_), .A3(new_n658_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n213_), .A3(new_n521_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n610_), .A2(new_n597_), .A3(new_n354_), .ZN(new_n737_));
  OR3_X1    g536(.A1(new_n666_), .A2(new_n668_), .A3(KEYINPUT111), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT111), .B1(new_n666_), .B2(new_n668_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(new_n521_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n736_), .B1(new_n741_), .B2(new_n213_), .ZN(G1336gat));
  NAND3_X1  g541(.A1(new_n735_), .A2(new_n214_), .A3(new_n497_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n740_), .A2(new_n497_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(new_n214_), .ZN(G1337gat));
  AOI21_X1  g544(.A(new_n205_), .B1(new_n740_), .B2(new_n645_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n735_), .A2(new_n645_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT51), .B1(new_n746_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750_));
  AOI211_X1 g549(.A(new_n570_), .B(new_n737_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n750_), .B(new_n747_), .C1(new_n751_), .C2(new_n205_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n752_), .ZN(G1338gat));
  NAND3_X1  g552(.A1(new_n735_), .A2(new_n206_), .A3(new_n651_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n666_), .A2(new_n668_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n737_), .A2(new_n574_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n755_), .B1(new_n758_), .B2(G106gat), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT52), .B(new_n206_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n754_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n754_), .B(new_n762_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1339gat));
  NOR3_X1   g565(.A1(new_n706_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n316_), .A2(new_n321_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT113), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n316_), .A2(new_n321_), .A3(new_n767_), .A4(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n769_), .A2(KEYINPUT54), .A3(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT57), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n615_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n271_), .A2(new_n276_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n596_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n587_), .B1(new_n581_), .B2(KEYINPUT118), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(KEYINPUT118), .B2(new_n581_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n586_), .A2(new_n583_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n595_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n780_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n271_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n597_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n256_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n274_), .A2(KEYINPUT55), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n273_), .A2(new_n263_), .A3(new_n254_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n273_), .A2(KEYINPUT114), .A3(new_n263_), .A4(new_n254_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n794_), .A2(new_n795_), .A3(new_n798_), .A4(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT115), .B1(new_n800_), .B2(new_n260_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(KEYINPUT56), .A3(new_n260_), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n792_), .A2(new_n801_), .B1(new_n802_), .B2(KEYINPUT116), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n792_), .A2(KEYINPUT116), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n798_), .A2(new_n799_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n273_), .A2(new_n254_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT55), .B1(new_n806_), .B2(new_n202_), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n793_), .B(new_n263_), .C1(new_n273_), .C2(new_n254_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n261_), .B1(new_n805_), .B2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n804_), .B1(new_n810_), .B2(KEYINPUT115), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n791_), .B1(new_n803_), .B2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n788_), .B1(new_n812_), .B2(KEYINPUT117), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n802_), .A2(KEYINPUT116), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n800_), .A2(new_n260_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n792_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n811_), .A2(new_n814_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n790_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n778_), .B1(new_n813_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT120), .B1(new_n810_), .B2(KEYINPUT56), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n815_), .A2(new_n824_), .A3(new_n792_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n802_), .A2(KEYINPUT119), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n810_), .A2(new_n827_), .A3(KEYINPUT56), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n823_), .A2(new_n825_), .A3(new_n826_), .A4(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n786_), .A2(new_n789_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n829_), .A2(KEYINPUT58), .A3(new_n830_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n322_), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n787_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n812_), .A2(KEYINPUT117), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n615_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n822_), .B(new_n835_), .C1(new_n838_), .C2(KEYINPUT57), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n776_), .B1(new_n839_), .B2(new_n354_), .ZN(new_n840_));
  NOR4_X1   g639(.A1(new_n651_), .A2(new_n497_), .A3(new_n572_), .A4(new_n570_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(G113gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n598_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n836_), .A2(new_n837_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n834_), .A2(new_n322_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n848_), .A2(new_n778_), .B1(new_n849_), .B2(new_n833_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n615_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n813_), .B2(new_n821_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n777_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n612_), .B1(new_n850_), .B2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT59), .B(new_n841_), .C1(new_n854_), .C2(new_n776_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n597_), .B1(new_n847_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n845_), .B1(new_n856_), .B2(new_n844_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT121), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n859_), .B(new_n845_), .C1(new_n856_), .C2(new_n844_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(G1340gat));
  NOR2_X1   g660(.A1(new_n280_), .A2(KEYINPUT60), .ZN(new_n862_));
  MUX2_X1   g661(.A(new_n862_), .B(KEYINPUT60), .S(G120gat), .Z(new_n863_));
  NAND2_X1  g662(.A1(new_n843_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n281_), .B1(new_n847_), .B2(new_n855_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n865_), .A2(KEYINPUT122), .ZN(new_n866_));
  OAI21_X1  g665(.A(G120gat), .B1(new_n865_), .B2(KEYINPUT122), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n864_), .B1(new_n866_), .B2(new_n867_), .ZN(G1341gat));
  INV_X1    g667(.A(G127gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n843_), .A2(new_n869_), .A3(new_n612_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n354_), .B1(new_n847_), .B2(new_n855_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n869_), .ZN(G1342gat));
  INV_X1    g671(.A(G134gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n843_), .A2(new_n873_), .A3(new_n615_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n322_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n847_), .B2(new_n855_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n874_), .B1(new_n876_), .B2(new_n873_), .ZN(G1343gat));
  NOR2_X1   g676(.A1(new_n574_), .A2(new_n645_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR4_X1   g678(.A1(new_n840_), .A2(new_n497_), .A3(new_n572_), .A4(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n598_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g681(.A1(new_n840_), .A2(new_n879_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n497_), .A2(new_n572_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n281_), .ZN(new_n886_));
  XOR2_X1   g685(.A(KEYINPUT123), .B(G148gat), .Z(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1345gat));
  NAND2_X1  g687(.A1(new_n880_), .A2(new_n612_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT61), .B(G155gat), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1346gat));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892_));
  INV_X1    g691(.A(G162gat), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n893_), .B1(new_n880_), .B2(new_n322_), .ZN(new_n894_));
  AND4_X1   g693(.A1(new_n893_), .A2(new_n883_), .A3(new_n615_), .A4(new_n884_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n892_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G162gat), .B1(new_n885_), .B2(new_n875_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n880_), .A2(new_n893_), .A3(new_n615_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n897_), .A2(new_n898_), .A3(KEYINPUT124), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n899_), .ZN(G1347gat));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n839_), .A2(new_n354_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n776_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n573_), .A2(new_n574_), .A3(new_n497_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n598_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n901_), .B1(new_n908_), .B2(G169gat), .ZN(new_n909_));
  AOI211_X1 g708(.A(KEYINPUT62), .B(new_n451_), .C1(new_n907_), .C2(new_n598_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT22), .B(G169gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n598_), .A2(new_n911_), .ZN(new_n912_));
  XOR2_X1   g711(.A(new_n912_), .B(KEYINPUT125), .Z(new_n913_));
  OAI22_X1  g712(.A1(new_n909_), .A2(new_n910_), .B1(new_n906_), .B2(new_n913_), .ZN(G1348gat));
  OAI21_X1  g713(.A(G176gat), .B1(new_n906_), .B2(new_n281_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n610_), .A2(new_n452_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n906_), .B2(new_n916_), .ZN(G1349gat));
  NOR2_X1   g716(.A1(new_n906_), .A2(new_n354_), .ZN(new_n918_));
  MUX2_X1   g717(.A(G183gat), .B(new_n446_), .S(new_n918_), .Z(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n906_), .B2(new_n875_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n615_), .A2(new_n447_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n906_), .B2(new_n921_), .ZN(G1351gat));
  NOR2_X1   g721(.A1(new_n575_), .A2(new_n521_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n883_), .A2(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n597_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n359_), .ZN(G1352gat));
  NOR2_X1   g725(.A1(new_n924_), .A2(new_n281_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(new_n361_), .ZN(G1353gat));
  NOR2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n929_), .B1(new_n924_), .B2(new_n354_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  OAI211_X1 g731(.A(KEYINPUT127), .B(new_n929_), .C1(new_n924_), .C2(new_n354_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n883_), .A2(new_n923_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935_));
  XOR2_X1   g734(.A(KEYINPUT63), .B(G211gat), .Z(new_n936_));
  NAND4_X1  g735(.A1(new_n934_), .A2(new_n935_), .A3(new_n612_), .A4(new_n936_), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n883_), .A2(new_n612_), .A3(new_n923_), .A4(new_n936_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(KEYINPUT126), .ZN(new_n939_));
  AOI22_X1  g738(.A1(new_n932_), .A2(new_n933_), .B1(new_n937_), .B2(new_n939_), .ZN(G1354gat));
  OAI21_X1  g739(.A(G218gat), .B1(new_n924_), .B2(new_n875_), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n851_), .A2(G218gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n924_), .B2(new_n942_), .ZN(G1355gat));
endmodule


