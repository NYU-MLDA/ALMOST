//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n839_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_;
  INV_X1    g000(.A(G230gat), .ZN(new_n202_));
  INV_X1    g001(.A(G233gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G57gat), .ZN(new_n205_));
  INV_X1    g004(.A(G64gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G57gat), .A2(G64gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT11), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(new_n211_), .A3(new_n208_), .ZN(new_n212_));
  AND2_X1   g011(.A1(KEYINPUT65), .A2(G71gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT65), .A2(G71gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(G78gat), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(KEYINPUT65), .A2(G71gat), .ZN(new_n216_));
  INV_X1    g015(.A(G78gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(KEYINPUT65), .A2(G71gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n210_), .A2(new_n212_), .A3(new_n215_), .A4(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n215_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n211_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(G99gat), .ZN(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT6), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n228_), .A2(new_n231_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT8), .ZN(new_n235_));
  AND2_X1   g034(.A1(G85gat), .A2(G92gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G85gat), .A2(G92gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n234_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n235_), .B1(new_n234_), .B2(new_n238_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT9), .ZN(new_n243_));
  INV_X1    g042(.A(G85gat), .ZN(new_n244_));
  INV_X1    g043(.A(G92gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G85gat), .A2(G92gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n243_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n243_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n242_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n226_), .A2(KEYINPUT10), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT10), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G99gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(G106gat), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n231_), .A2(new_n232_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(KEYINPUT64), .B(new_n249_), .C1(new_n238_), .C2(new_n243_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n251_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n224_), .B1(new_n241_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n220_), .A2(new_n223_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n251_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n261_), .B(new_n262_), .C1(new_n240_), .C2(new_n239_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(KEYINPUT12), .A3(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n262_), .B1(new_n240_), .B2(new_n239_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT12), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(new_n224_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n204_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n260_), .A2(new_n263_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n204_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G120gat), .B(G148gat), .ZN(new_n273_));
  INV_X1    g072(.A(G204gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT5), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(G176gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n272_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT13), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n274_), .A2(G197gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT21), .B1(new_n281_), .B2(KEYINPUT88), .ZN(new_n282_));
  XOR2_X1   g081(.A(G211gat), .B(G218gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(G197gat), .B(G204gat), .ZN(new_n284_));
  OR3_X1    g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT21), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n284_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT89), .Z(new_n290_));
  NAND2_X1  g089(.A1(G228gat), .A2(G233gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n291_), .B(KEYINPUT87), .Z(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G155gat), .B(G162gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n294_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n294_), .B(KEYINPUT3), .Z(new_n302_));
  XOR2_X1   g101(.A(new_n300_), .B(KEYINPUT2), .Z(new_n303_));
  OAI21_X1  g102(.A(new_n296_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT29), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n290_), .A2(new_n293_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n306_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n292_), .B1(new_n308_), .B2(new_n289_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n305_), .A2(KEYINPUT29), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n310_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G22gat), .B(G50gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(G78gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(G106gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n314_), .A2(new_n318_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G127gat), .B(G134gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G113gat), .B(G120gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n327_), .A2(KEYINPUT31), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(KEYINPUT31), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(KEYINPUT83), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G227gat), .A2(G233gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT80), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(KEYINPUT23), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(KEYINPUT23), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT80), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n335_), .B(new_n337_), .C1(KEYINPUT23), .C2(new_n333_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(G183gat), .B2(G190gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT81), .ZN(new_n340_));
  AND2_X1   g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT22), .B(G169gat), .ZN(new_n342_));
  INV_X1    g141(.A(G176gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n341_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n340_), .B(new_n346_), .C1(new_n345_), .C2(new_n344_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT77), .B1(new_n333_), .B2(KEYINPUT23), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(new_n336_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT24), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n353_), .B(KEYINPUT78), .Z(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT25), .B(G183gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G190gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n341_), .A2(new_n350_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n355_), .A2(new_n356_), .B1(new_n357_), .B2(KEYINPUT24), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n354_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n347_), .A2(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(KEYINPUT82), .B(KEYINPUT30), .Z(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n332_), .B(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G15gat), .B(G43gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(G71gat), .B(G99gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n363_), .A2(new_n366_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n305_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n327_), .B(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(KEYINPUT4), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n327_), .A2(new_n305_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(KEYINPUT4), .B2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n374_), .B1(new_n377_), .B2(new_n373_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G1gat), .B(G29gat), .Z(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G57gat), .B(G85gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n378_), .B(new_n383_), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n289_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n360_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT19), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n349_), .B1(G183gat), .B2(G190gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n358_), .A2(new_n338_), .A3(new_n352_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n289_), .A3(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT90), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n387_), .A2(KEYINPUT20), .A3(new_n390_), .A4(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT91), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n394_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n386_), .ZN(new_n400_));
  OAI211_X1 g199(.A(KEYINPUT20), .B(new_n400_), .C1(new_n360_), .C2(new_n386_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n389_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(G8gat), .B(G36gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n406_), .B(new_n407_), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT32), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n385_), .B1(new_n403_), .B2(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n401_), .A2(new_n389_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n387_), .B(KEYINPUT20), .C1(new_n290_), .C2(new_n399_), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n413_), .A2(KEYINPUT95), .B1(new_n389_), .B2(new_n414_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n414_), .A2(KEYINPUT95), .A3(new_n389_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n411_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT96), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n417_), .A2(new_n418_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n412_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n403_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n409_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n378_), .A2(new_n383_), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n424_), .B(KEYINPUT33), .Z(new_n425_));
  NAND2_X1  g224(.A1(new_n403_), .A2(new_n408_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n373_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n372_), .A2(new_n427_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n383_), .B(new_n428_), .C1(new_n377_), .C2(new_n427_), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n429_), .B(KEYINPUT94), .Z(new_n430_));
  AND4_X1   g229(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .A4(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n322_), .B(new_n370_), .C1(new_n421_), .C2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n370_), .A2(new_n322_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n423_), .A2(new_n426_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n385_), .B1(new_n369_), .B2(new_n321_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n408_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n423_), .A2(KEYINPUT27), .A3(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n433_), .A2(new_n436_), .A3(new_n437_), .A4(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n280_), .B1(new_n432_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT37), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G190gat), .B(G218gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(G134gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(G162gat), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(KEYINPUT36), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G29gat), .B(G36gat), .ZN(new_n447_));
  INV_X1    g246(.A(G43gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(G50gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT15), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n265_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G232gat), .A2(G233gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT34), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT35), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n450_), .A2(new_n265_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n453_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n456_), .A2(new_n457_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n461_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n453_), .A2(new_n463_), .A3(new_n458_), .A4(new_n459_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n446_), .B1(new_n465_), .B2(KEYINPUT66), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT66), .ZN(new_n467_));
  INV_X1    g266(.A(new_n446_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n462_), .A2(new_n467_), .A3(new_n468_), .A4(new_n464_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n465_), .A2(KEYINPUT36), .A3(new_n445_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n466_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n442_), .B1(new_n472_), .B2(KEYINPUT67), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT67), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n474_), .A3(KEYINPUT37), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G231gat), .A2(G233gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n224_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G8gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G15gat), .ZN(new_n482_));
  INV_X1    g281(.A(G22gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G15gat), .A2(G22gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G1gat), .A2(G8gat), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n484_), .A2(new_n485_), .B1(KEYINPUT14), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n481_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n478_), .B(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G127gat), .B(G155gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT70), .B(KEYINPUT16), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G183gat), .B(G211gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n489_), .A2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n497_), .B(KEYINPUT71), .Z(new_n498_));
  AND2_X1   g297(.A1(new_n494_), .A2(new_n495_), .ZN(new_n499_));
  OR3_X1    g298(.A1(new_n489_), .A2(new_n496_), .A3(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n476_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n452_), .A2(new_n488_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT73), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G229gat), .A2(G233gat), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n488_), .A2(new_n450_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT72), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n452_), .A2(KEYINPUT73), .A3(new_n488_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n506_), .A2(new_n507_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n488_), .A2(new_n450_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n507_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n512_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G169gat), .B(G197gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(G141gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT75), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(G113gat), .Z(new_n521_));
  OR2_X1    g320(.A1(new_n521_), .A2(KEYINPUT74), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n517_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT76), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n512_), .A2(new_n516_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(new_n522_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT76), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n441_), .A2(new_n503_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(G1gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n384_), .B(KEYINPUT97), .Z(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT38), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n535_), .B(KEYINPUT98), .Z(new_n536_));
  AOI21_X1  g335(.A(new_n471_), .B1(new_n432_), .B2(new_n440_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n523_), .A2(new_n279_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT99), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n537_), .A2(new_n501_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n531_), .B1(new_n540_), .B2(new_n385_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n534_), .B2(new_n533_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n536_), .A2(new_n542_), .ZN(G1324gat));
  INV_X1    g342(.A(G8gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n436_), .A2(new_n439_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n530_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT100), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n530_), .A2(KEYINPUT100), .A3(new_n544_), .A4(new_n545_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n544_), .B1(new_n540_), .B2(new_n545_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT39), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT39), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n537_), .A2(new_n501_), .A3(new_n539_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n545_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n553_), .B1(new_n556_), .B2(new_n544_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n550_), .A2(new_n552_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT101), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT101), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n550_), .A2(new_n557_), .A3(new_n560_), .A4(new_n552_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT40), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n559_), .A2(new_n561_), .A3(KEYINPUT40), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(G1325gat));
  NAND3_X1  g365(.A1(new_n530_), .A2(new_n482_), .A3(new_n369_), .ZN(new_n567_));
  OAI21_X1  g366(.A(G15gat), .B1(new_n554_), .B2(new_n370_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT102), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(KEYINPUT102), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n570_), .A2(KEYINPUT41), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT41), .B1(new_n570_), .B2(new_n571_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n567_), .B1(new_n572_), .B2(new_n573_), .ZN(G1326gat));
  OAI21_X1  g373(.A(G22gat), .B1(new_n554_), .B2(new_n322_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT42), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n321_), .A2(new_n483_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT103), .Z(new_n578_));
  NAND2_X1  g377(.A1(new_n530_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT104), .Z(G1327gat));
  NOR2_X1   g380(.A1(new_n472_), .A2(new_n501_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n441_), .A2(new_n529_), .A3(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(G29gat), .B1(new_n583_), .B2(new_n385_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n432_), .A2(new_n440_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n476_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT43), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT43), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n588_), .A3(new_n476_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n590_), .A2(KEYINPUT44), .A3(new_n502_), .A4(new_n539_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n588_), .B1(new_n585_), .B2(new_n476_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n476_), .ZN(new_n593_));
  AOI211_X1 g392(.A(KEYINPUT43), .B(new_n593_), .C1(new_n432_), .C2(new_n440_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n502_), .B(new_n539_), .C1(new_n592_), .C2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT44), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n591_), .A2(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n598_), .A2(G29gat), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n584_), .B1(new_n599_), .B2(new_n532_), .ZN(G1328gat));
  INV_X1    g399(.A(KEYINPUT105), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT46), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n591_), .A2(new_n597_), .A3(new_n545_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(G36gat), .ZN(new_n605_));
  INV_X1    g404(.A(G36gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n583_), .A2(new_n606_), .A3(new_n545_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT45), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n603_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(G1329gat));
  NOR2_X1   g410(.A1(new_n370_), .A2(new_n448_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n591_), .A2(new_n597_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT106), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n591_), .A2(new_n597_), .A3(KEYINPUT106), .A4(new_n612_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n583_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n448_), .B1(new_n618_), .B2(new_n370_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT47), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT47), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(new_n622_), .A3(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(G1330gat));
  AOI21_X1  g423(.A(G50gat), .B1(new_n583_), .B2(new_n321_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n321_), .A2(G50gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n598_), .B2(new_n626_), .ZN(G1331gat));
  INV_X1    g426(.A(new_n529_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n537_), .A2(new_n501_), .A3(new_n628_), .A4(new_n280_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT107), .Z(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(G57gat), .A3(new_n385_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n523_), .A2(new_n279_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n585_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n503_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n532_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n205_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n631_), .A2(new_n636_), .ZN(G1332gat));
  INV_X1    g436(.A(new_n634_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n206_), .A3(new_n545_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n630_), .A2(new_n545_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G64gat), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(KEYINPUT48), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(KEYINPUT48), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n639_), .B1(new_n642_), .B2(new_n643_), .ZN(G1333gat));
  OR3_X1    g443(.A1(new_n634_), .A2(G71gat), .A3(new_n370_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n630_), .A2(new_n369_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(G71gat), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(KEYINPUT49), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(KEYINPUT49), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(G1334gat));
  NAND3_X1  g449(.A1(new_n638_), .A2(new_n217_), .A3(new_n321_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n630_), .A2(new_n321_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(G78gat), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n653_), .A2(KEYINPUT50), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(KEYINPUT50), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n651_), .B1(new_n654_), .B2(new_n655_), .ZN(G1335gat));
  AND2_X1   g455(.A1(new_n633_), .A2(new_n582_), .ZN(new_n657_));
  AOI21_X1  g456(.A(G85gat), .B1(new_n657_), .B2(new_n532_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n632_), .A2(new_n502_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT109), .Z(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n592_), .A2(new_n594_), .A3(KEYINPUT108), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(new_n384_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n658_), .B1(new_n666_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g466(.A(G92gat), .B1(new_n657_), .B2(new_n545_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n665_), .A2(new_n555_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(G92gat), .ZN(G1337gat));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n369_), .B(new_n661_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G99gat), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n252_), .A2(new_n254_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n657_), .A2(new_n674_), .A3(new_n369_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n671_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n673_), .A2(new_n671_), .A3(new_n675_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(KEYINPUT51), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT51), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n673_), .A2(new_n671_), .A3(new_n675_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n681_), .B2(new_n676_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(G1338gat));
  NAND3_X1  g482(.A1(new_n590_), .A2(new_n321_), .A3(new_n661_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G106gat), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT52), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n657_), .A2(new_n227_), .A3(new_n321_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT53), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT53), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n686_), .A2(new_n690_), .A3(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1339gat));
  NOR2_X1   g491(.A1(new_n545_), .A2(new_n635_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(new_n322_), .A3(new_n369_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n264_), .A2(new_n204_), .A3(new_n267_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT113), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(new_n697_), .A3(KEYINPUT55), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n696_), .B2(KEYINPUT55), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n269_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n696_), .A2(KEYINPUT55), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT113), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n696_), .A2(new_n697_), .A3(KEYINPUT55), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n268_), .A3(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n700_), .A2(new_n704_), .A3(new_n277_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT56), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n506_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n515_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n510_), .A2(new_n507_), .A3(new_n513_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n521_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n521_), .B2(new_n517_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n707_), .A2(new_n712_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n272_), .A2(new_n277_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT117), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT58), .ZN(new_n716_));
  AOI22_X1  g515(.A1(new_n713_), .A2(new_n714_), .B1(KEYINPUT116), .B2(new_n716_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n707_), .A2(new_n712_), .A3(KEYINPUT116), .A4(new_n714_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT58), .B1(new_n718_), .B2(new_n715_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n476_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT114), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n705_), .A2(new_n721_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n700_), .A2(new_n704_), .A3(KEYINPUT114), .A4(new_n277_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n706_), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT115), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n705_), .A2(new_n706_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT115), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n722_), .A2(new_n727_), .A3(new_n706_), .A4(new_n723_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n725_), .A2(new_n726_), .A3(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n523_), .A2(new_n714_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n712_), .A2(new_n278_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n471_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n720_), .B1(new_n733_), .B2(KEYINPUT57), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT118), .B1(new_n733_), .B2(KEYINPUT57), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n729_), .A2(new_n730_), .B1(new_n278_), .B2(new_n712_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT118), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT57), .ZN(new_n738_));
  NOR4_X1   g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .A4(new_n471_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n734_), .A2(new_n735_), .A3(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(new_n501_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n525_), .A2(new_n501_), .A3(new_n528_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n525_), .A2(KEYINPUT111), .A3(new_n501_), .A4(new_n528_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n593_), .A2(new_n744_), .A3(new_n279_), .A4(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT112), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n745_), .A2(new_n475_), .A3(new_n473_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n279_), .A4(new_n744_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT54), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n747_), .A2(new_n750_), .A3(KEYINPUT54), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n695_), .B1(new_n741_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G113gat), .B1(new_n757_), .B2(new_n523_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT120), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n759_), .B1(new_n740_), .B2(new_n501_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n754_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT54), .B1(new_n747_), .B2(new_n750_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n733_), .A2(KEYINPUT57), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n737_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n733_), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(KEYINPUT120), .B(new_n502_), .C1(new_n767_), .C2(new_n734_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n760_), .A2(new_n763_), .A3(new_n768_), .ZN(new_n769_));
  XOR2_X1   g568(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n695_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n756_), .A2(KEYINPUT59), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n773_), .A2(new_n628_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n758_), .B1(new_n774_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g574(.A(KEYINPUT122), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(new_n773_), .B2(new_n279_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n771_), .A2(new_n772_), .A3(KEYINPUT122), .A4(new_n280_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(G120gat), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(G120gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n279_), .B2(KEYINPUT60), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT121), .B1(new_n780_), .B2(KEYINPUT60), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n756_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT121), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n779_), .A2(new_n785_), .ZN(G1341gat));
  AOI21_X1  g585(.A(G127gat), .B1(new_n757_), .B2(new_n501_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n771_), .A2(G127gat), .A3(new_n772_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n501_), .ZN(G1342gat));
  NAND2_X1  g588(.A1(new_n476_), .A2(G134gat), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT123), .Z(new_n791_));
  NOR2_X1   g590(.A1(new_n756_), .A2(new_n472_), .ZN(new_n792_));
  OAI22_X1  g591(.A1(new_n773_), .A2(new_n791_), .B1(G134gat), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT124), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(G1343gat));
  NOR2_X1   g594(.A1(new_n741_), .A2(new_n755_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(new_n322_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n797_), .A2(new_n370_), .A3(new_n693_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(new_n527_), .ZN(new_n799_));
  INV_X1    g598(.A(G141gat), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(G1344gat));
  NOR2_X1   g600(.A1(new_n798_), .A2(new_n279_), .ZN(new_n802_));
  INV_X1    g601(.A(G148gat), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n802_), .B(new_n803_), .ZN(G1345gat));
  NOR2_X1   g603(.A1(new_n798_), .A2(new_n502_), .ZN(new_n805_));
  XOR2_X1   g604(.A(KEYINPUT61), .B(G155gat), .Z(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1346gat));
  NOR2_X1   g606(.A1(new_n798_), .A2(new_n472_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n808_), .A2(G162gat), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n798_), .A2(new_n593_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(G162gat), .B2(new_n810_), .ZN(G1347gat));
  NOR3_X1   g610(.A1(new_n555_), .A2(new_n532_), .A3(new_n370_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n812_), .A2(new_n523_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n769_), .A2(new_n322_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(G169gat), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT62), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n769_), .A2(new_n322_), .A3(new_n342_), .A4(new_n813_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n814_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT125), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n817_), .A2(new_n818_), .A3(KEYINPUT125), .A4(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1348gat));
  OAI211_X1 g623(.A(new_n322_), .B(new_n812_), .C1(new_n741_), .C2(new_n755_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n825_), .A2(new_n343_), .A3(new_n279_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n769_), .A2(new_n322_), .A3(new_n812_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n280_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n826_), .B1(new_n828_), .B2(new_n343_), .ZN(G1349gat));
  INV_X1    g628(.A(new_n355_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(new_n501_), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT126), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n831_), .A2(new_n832_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n825_), .A2(new_n502_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(G183gat), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n833_), .A2(new_n834_), .A3(new_n836_), .ZN(G1350gat));
  INV_X1    g636(.A(new_n827_), .ZN(new_n838_));
  OAI21_X1  g637(.A(G190gat), .B1(new_n838_), .B2(new_n593_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n827_), .A2(new_n471_), .A3(new_n356_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1351gat));
  NAND2_X1  g640(.A1(new_n437_), .A2(new_n321_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n796_), .B1(KEYINPUT127), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT127), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n555_), .B1(new_n845_), .B2(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n527_), .ZN(new_n848_));
  INV_X1    g647(.A(G197gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1352gat));
  NOR2_X1   g649(.A1(new_n847_), .A2(new_n279_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(new_n274_), .ZN(G1353gat));
  INV_X1    g651(.A(new_n847_), .ZN(new_n853_));
  XOR2_X1   g652(.A(KEYINPUT63), .B(G211gat), .Z(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n501_), .A3(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n847_), .B2(new_n502_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1354gat));
  AOI21_X1  g657(.A(G218gat), .B1(new_n853_), .B2(new_n471_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n847_), .A2(new_n593_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(G218gat), .B2(new_n860_), .ZN(G1355gat));
endmodule


