//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n943_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_, new_n962_;
  INV_X1    g000(.A(G141gat), .ZN(new_n202_));
  INV_X1    g001(.A(G148gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT88), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209_));
  AND2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n211_), .A2(KEYINPUT89), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT89), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n208_), .B(new_n213_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n210_), .A2(new_n209_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n206_), .B1(new_n212_), .B2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n204_), .B(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n205_), .B(KEYINPUT2), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n210_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n208_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n217_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G127gat), .B(G134gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT87), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G120gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n224_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n223_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n211_), .A2(KEYINPUT89), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(new_n215_), .A3(new_n214_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n231_), .B1(new_n233_), .B2(new_n206_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n228_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(new_n235_), .A3(KEYINPUT4), .ZN(new_n236_));
  OR3_X1    g035(.A1(new_n234_), .A2(KEYINPUT4), .A3(new_n228_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G1gat), .B(G29gat), .Z(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT99), .B(G85gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT0), .B(G57gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n230_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n240_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n246_), .B1(new_n240_), .B2(new_n247_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT79), .B(G183gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT25), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT80), .B(G190gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT26), .ZN(new_n255_));
  OR2_X1    g054(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n251_), .A2(new_n253_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT24), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(G169gat), .B2(G176gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT81), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(G169gat), .B2(G176gat), .ZN(new_n261_));
  INV_X1    g060(.A(G169gat), .ZN(new_n262_));
  INV_X1    g061(.A(G176gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT81), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n259_), .A2(new_n261_), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT24), .B1(new_n264_), .B2(new_n261_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n257_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT23), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n268_), .B(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n271_), .B1(new_n273_), .B2(new_n270_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n269_), .A2(KEYINPUT23), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n276_), .B1(new_n273_), .B2(KEYINPUT23), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT22), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT83), .B1(new_n279_), .B2(G169gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT22), .B(G169gat), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n263_), .B(new_n280_), .C1(new_n281_), .C2(KEYINPUT83), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n267_), .A2(new_n275_), .B1(new_n278_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G227gat), .A2(G233gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n286_), .B(KEYINPUT86), .Z(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n285_), .A2(new_n288_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n292_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n294_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G15gat), .B(G43gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT85), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G71gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n299_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n293_), .A2(new_n295_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n228_), .B(KEYINPUT31), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(G99gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n305_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n250_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G22gat), .B(G50gat), .Z(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n217_), .A2(new_n312_), .A3(new_n223_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT28), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT28), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n234_), .A2(new_n315_), .A3(new_n312_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT91), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n314_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n311_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n314_), .A2(new_n316_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT91), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n314_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n310_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n224_), .A2(KEYINPUT29), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G211gat), .B(G218gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n327_), .B(KEYINPUT93), .Z(new_n328_));
  INV_X1    g127(.A(G197gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT92), .B1(new_n329_), .B2(G204gat), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT92), .ZN(new_n331_));
  INV_X1    g130(.A(G204gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(G197gat), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n330_), .B(new_n333_), .C1(G197gat), .C2(new_n332_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n328_), .A2(KEYINPUT21), .A3(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n334_), .A2(KEYINPUT21), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n327_), .B(KEYINPUT93), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n329_), .A2(G204gat), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n332_), .A2(G197gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT21), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(new_n337_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT94), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n336_), .A2(new_n337_), .A3(KEYINPUT94), .A4(new_n340_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n335_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G228gat), .A2(G233gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n326_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n312_), .B1(new_n217_), .B2(new_n223_), .ZN(new_n349_));
  OAI211_X1 g148(.A(G228gat), .B(G233gat), .C1(new_n349_), .C2(new_n345_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G78gat), .B(G106gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n351_), .B(KEYINPUT95), .Z(new_n352_));
  AND3_X1   g151(.A1(new_n348_), .A2(new_n350_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n352_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n325_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n351_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n353_), .A2(new_n359_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n325_), .A2(new_n360_), .A3(KEYINPUT96), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT96), .B1(new_n325_), .B2(new_n360_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n357_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT18), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n281_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370_));
  OAI221_X1 g169(.A(new_n283_), .B1(G176gat), .B2(new_n369_), .C1(new_n274_), .C2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n259_), .A2(KEYINPUT98), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n259_), .A2(KEYINPUT98), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n261_), .A4(new_n264_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT25), .B(G183gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT26), .B(G190gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n258_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n374_), .A2(new_n277_), .A3(new_n377_), .A4(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n371_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n345_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT20), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G226gat), .A2(G233gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n345_), .A2(new_n285_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n382_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n345_), .A2(new_n380_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT20), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n345_), .B2(new_n285_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n385_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n368_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n391_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n386_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n387_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n396_), .A2(KEYINPUT20), .A3(new_n385_), .A4(new_n381_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n395_), .A2(new_n367_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT27), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n393_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(KEYINPUT101), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT101), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n395_), .A2(new_n397_), .A3(new_n402_), .A4(new_n367_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n386_), .B1(new_n382_), .B2(new_n387_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n389_), .A2(new_n385_), .A3(new_n391_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n368_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n401_), .A2(new_n403_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n400_), .B1(new_n408_), .B2(KEYINPUT27), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n309_), .A2(new_n363_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n325_), .A2(new_n360_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT96), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n325_), .A2(new_n360_), .A3(KEYINPUT96), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n356_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n367_), .A2(KEYINPUT32), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT100), .B1(new_n406_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT100), .ZN(new_n419_));
  AOI211_X1 g218(.A(new_n419_), .B(new_n416_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n395_), .A2(new_n397_), .A3(new_n416_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n422_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n240_), .A2(KEYINPUT33), .A3(new_n246_), .A4(new_n247_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n230_), .A2(new_n235_), .A3(new_n239_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n245_), .A3(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n393_), .A2(new_n398_), .A3(new_n424_), .A4(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n248_), .A2(KEYINPUT33), .ZN(new_n429_));
  OAI22_X1  g228(.A1(new_n421_), .A2(new_n423_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n415_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n363_), .A2(new_n250_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n431_), .B1(new_n432_), .B2(new_n409_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n307_), .A2(new_n308_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n410_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G29gat), .B(G36gat), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n436_), .A2(KEYINPUT72), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(KEYINPUT72), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G43gat), .B(G50gat), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n439_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G15gat), .B(G22gat), .ZN(new_n443_));
  INV_X1    g242(.A(G1gat), .ZN(new_n444_));
  INV_X1    g243(.A(G8gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT14), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G1gat), .B(G8gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n442_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n449_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G229gat), .A2(G233gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT15), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n437_), .A2(new_n438_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n439_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(KEYINPUT15), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n450_), .B1(new_n458_), .B2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n454_), .B(KEYINPUT77), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n451_), .A2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n456_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G113gat), .B(G141gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G169gat), .B(G197gat), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n468_), .B(new_n469_), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n467_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT78), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n456_), .B(new_n470_), .C1(new_n464_), .C2(new_n466_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n467_), .A2(KEYINPUT78), .A3(new_n471_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n435_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G120gat), .B(G148gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT5), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G176gat), .B(G204gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT69), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT68), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G230gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  AND2_X1   g287(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(G78gat), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT66), .ZN(new_n492_));
  INV_X1    g291(.A(G71gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G78gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n491_), .A2(new_n497_), .B1(new_n498_), .B2(KEYINPUT11), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT11), .ZN(new_n500_));
  INV_X1    g299(.A(G57gat), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n501_), .A2(G64gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(G64gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n500_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n491_), .A2(new_n497_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n499_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT7), .ZN(new_n509_));
  INV_X1    g308(.A(G99gat), .ZN(new_n510_));
  INV_X1    g309(.A(G106gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT65), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT6), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(G99gat), .A3(G106gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT65), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n512_), .A2(new_n521_), .A3(new_n513_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n515_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(G85gat), .ZN(new_n524_));
  INV_X1    g323(.A(G92gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n528_), .A2(KEYINPUT8), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n517_), .A2(new_n519_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n528_), .B1(new_n530_), .B2(new_n514_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT8), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n523_), .A2(new_n529_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT64), .ZN(new_n534_));
  OR2_X1    g333(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n511_), .A3(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n526_), .A2(KEYINPUT9), .A3(new_n527_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT9), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(G85gat), .A3(G92gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n520_), .A2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n534_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n527_), .A2(KEYINPUT9), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n545_), .A2(KEYINPUT64), .A3(new_n537_), .A4(new_n538_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n508_), .B1(new_n533_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT67), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n523_), .A2(new_n529_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n531_), .A2(new_n532_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n547_), .A2(new_n508_), .A3(new_n550_), .A4(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n548_), .B1(new_n549_), .B2(new_n552_), .ZN(new_n553_));
  AOI211_X1 g352(.A(KEYINPUT67), .B(new_n508_), .C1(new_n533_), .C2(new_n547_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n486_), .B(new_n488_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(KEYINPUT12), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(new_n548_), .ZN(new_n557_));
  AOI211_X1 g356(.A(KEYINPUT12), .B(new_n508_), .C1(new_n533_), .C2(new_n547_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n487_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n552_), .A2(new_n549_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n533_), .A2(new_n547_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n508_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n562_), .A2(new_n563_), .A3(new_n549_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n486_), .B1(new_n567_), .B2(new_n488_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n485_), .B1(new_n560_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT70), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n488_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT68), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n572_), .A2(new_n559_), .A3(new_n555_), .A4(new_n483_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n569_), .A2(new_n570_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n570_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT13), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT13), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n578_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT71), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT71), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n458_), .A2(new_n463_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n562_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT34), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT35), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n590_), .A2(new_n591_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n442_), .A2(new_n533_), .A3(new_n547_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n587_), .A2(new_n593_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n594_), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n458_), .A2(new_n463_), .B1(new_n533_), .B2(new_n547_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n592_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(G190gat), .B(G218gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT73), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  OAI22_X1  g403(.A1(new_n600_), .A2(KEYINPUT74), .B1(KEYINPUT36), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT74), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n604_), .A2(KEYINPUT36), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n596_), .A2(new_n599_), .A3(new_n606_), .A4(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n600_), .A2(KEYINPUT36), .A3(new_n604_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT37), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n609_), .A2(new_n613_), .A3(new_n610_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n449_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(new_n508_), .ZN(new_n618_));
  XOR2_X1   g417(.A(G127gat), .B(G155gat), .Z(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT17), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n618_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n617_), .B(new_n563_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(KEYINPUT17), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT76), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n625_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n625_), .B2(new_n628_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AND4_X1   g432(.A1(new_n479_), .A2(new_n585_), .A3(new_n615_), .A4(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n250_), .A2(G1gat), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OR3_X1    g435(.A1(new_n636_), .A2(KEYINPUT103), .A3(KEYINPUT38), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT103), .B1(new_n636_), .B2(KEYINPUT38), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n435_), .A2(new_n611_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n581_), .A2(new_n478_), .A3(new_n632_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n250_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n444_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n636_), .A2(KEYINPUT102), .A3(KEYINPUT38), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n634_), .A2(KEYINPUT38), .A3(new_n635_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n644_), .B1(new_n645_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n639_), .A2(new_n649_), .ZN(G1324gat));
  NAND3_X1  g449(.A1(new_n640_), .A2(new_n409_), .A3(new_n641_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G8gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT39), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n634_), .A2(new_n445_), .A3(new_n409_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n655_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1325gat));
  INV_X1    g458(.A(G15gat), .ZN(new_n660_));
  INV_X1    g459(.A(new_n434_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n634_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n642_), .A2(new_n661_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n663_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT41), .B1(new_n663_), .B2(G15gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n662_), .B1(new_n664_), .B2(new_n665_), .ZN(G1326gat));
  INV_X1    g465(.A(G22gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n634_), .A2(new_n667_), .A3(new_n363_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n642_), .A2(new_n363_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G22gat), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n670_), .A2(KEYINPUT42), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(KEYINPUT42), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(G1327gat));
  NAND2_X1  g472(.A1(new_n611_), .A2(new_n632_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n581_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n479_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G29gat), .B1(new_n677_), .B2(new_n643_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT43), .B1(new_n435_), .B2(new_n615_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n612_), .A2(new_n614_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n409_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n250_), .A3(new_n363_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n661_), .B1(new_n683_), .B2(new_n431_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n680_), .B(new_n681_), .C1(new_n684_), .C2(new_n410_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n679_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n580_), .A2(new_n477_), .A3(new_n632_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT44), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  AOI211_X1 g489(.A(new_n690_), .B(new_n687_), .C1(new_n679_), .C2(new_n685_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n643_), .A2(G29gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n678_), .B1(new_n692_), .B2(new_n693_), .ZN(G1328gat));
  NOR2_X1   g493(.A1(new_n682_), .A2(G36gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OR3_X1    g495(.A1(new_n676_), .A2(KEYINPUT45), .A3(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT45), .B1(new_n676_), .B2(new_n696_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n689_), .A2(new_n691_), .A3(new_n682_), .ZN(new_n700_));
  INV_X1    g499(.A(G36gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n699_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(KEYINPUT46), .B(new_n699_), .C1(new_n700_), .C2(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  AOI21_X1  g505(.A(G43gat), .B1(new_n677_), .B2(new_n661_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n661_), .A2(G43gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n692_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT47), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(G1330gat));
  OR3_X1    g510(.A1(new_n676_), .A2(G50gat), .A3(new_n415_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n692_), .A2(new_n713_), .A3(new_n363_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G50gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n713_), .B1(new_n692_), .B2(new_n363_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(G1331gat));
  NOR2_X1   g516(.A1(new_n435_), .A2(new_n477_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n580_), .A2(new_n681_), .A3(new_n632_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n501_), .B1(new_n720_), .B2(new_n250_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT106), .Z(new_n722_));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n723_));
  INV_X1    g522(.A(new_n585_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n477_), .A2(new_n632_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n640_), .A2(new_n723_), .A3(new_n724_), .A4(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n611_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n727_), .B1(new_n684_), .B2(new_n410_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n582_), .A2(new_n584_), .A3(new_n725_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT107), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n726_), .A2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n250_), .A2(new_n501_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n722_), .B1(new_n731_), .B2(new_n732_), .ZN(G1332gat));
  OR3_X1    g532(.A1(new_n720_), .A2(G64gat), .A3(new_n682_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n409_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(G64gat), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G64gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1333gat));
  INV_X1    g538(.A(new_n720_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(new_n493_), .A3(new_n661_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT49), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n731_), .A2(new_n661_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(G71gat), .ZN(new_n744_));
  AOI211_X1 g543(.A(KEYINPUT49), .B(new_n493_), .C1(new_n731_), .C2(new_n661_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1334gat));
  NAND3_X1  g545(.A1(new_n740_), .A2(new_n495_), .A3(new_n363_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n726_), .A2(new_n730_), .A3(new_n363_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(new_n749_), .A3(G78gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n748_), .B2(G78gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  OAI211_X1 g553(.A(KEYINPUT109), .B(new_n747_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1335gat));
  NOR3_X1   g555(.A1(new_n580_), .A2(new_n477_), .A3(new_n633_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT110), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n686_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759_), .B2(new_n250_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n718_), .A2(new_n724_), .A3(new_n611_), .A4(new_n632_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n643_), .A2(new_n524_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(G1336gat));
  OAI21_X1  g562(.A(G92gat), .B1(new_n759_), .B2(new_n682_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n409_), .A2(new_n525_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n761_), .B2(new_n765_), .ZN(G1337gat));
  NOR2_X1   g565(.A1(new_n759_), .A2(new_n434_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n767_), .A2(new_n510_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n661_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n761_), .A2(new_n769_), .ZN(new_n770_));
  OR3_X1    g569(.A1(new_n768_), .A2(KEYINPUT51), .A3(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT51), .B1(new_n768_), .B2(new_n770_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1338gat));
  NAND3_X1  g572(.A1(new_n686_), .A2(new_n363_), .A3(new_n758_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(G106gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G106gat), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n363_), .A2(new_n511_), .ZN(new_n778_));
  OAI22_X1  g577(.A1(new_n776_), .A2(new_n777_), .B1(new_n761_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT53), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781_));
  OAI221_X1 g580(.A(new_n781_), .B1(new_n761_), .B2(new_n778_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1339gat));
  NAND4_X1  g582(.A1(new_n612_), .A2(new_n633_), .A3(new_n478_), .A4(new_n614_), .ZN(new_n784_));
  AOI211_X1 g583(.A(KEYINPUT54), .B(new_n784_), .C1(new_n577_), .C2(new_n579_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786_));
  INV_X1    g585(.A(new_n784_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n580_), .B2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n477_), .A2(new_n573_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n564_), .A2(KEYINPUT12), .A3(new_n552_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n558_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n488_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n559_), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n488_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT111), .B1(new_n798_), .B2(KEYINPUT55), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n559_), .A2(new_n800_), .A3(new_n796_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n797_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n792_), .B1(new_n802_), .B2(new_n484_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n557_), .A2(new_n487_), .A3(new_n558_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(KEYINPUT55), .B2(new_n798_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n798_), .A2(KEYINPUT111), .A3(KEYINPUT55), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n800_), .B1(new_n559_), .B2(new_n796_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n805_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(KEYINPUT56), .A3(new_n485_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n791_), .B1(new_n803_), .B2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n487_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n793_), .A2(new_n794_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n811_), .A2(new_n486_), .B1(new_n812_), .B2(new_n487_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n484_), .B1(new_n813_), .B2(new_n572_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n483_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n560_), .A2(new_n568_), .A3(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT70), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n569_), .A2(new_n570_), .A3(new_n573_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n586_), .A2(new_n449_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n465_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n451_), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n470_), .B1(new_n453_), .B2(new_n465_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT112), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n821_), .A2(new_n822_), .A3(new_n825_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n824_), .A2(new_n474_), .A3(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n817_), .A2(new_n818_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT113), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n817_), .A2(new_n830_), .A3(new_n818_), .A4(new_n827_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n810_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n790_), .B1(new_n832_), .B2(new_n611_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n810_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n830_), .B1(new_n576_), .B2(new_n827_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n831_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n611_), .A2(new_n790_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n824_), .A2(new_n474_), .A3(new_n826_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT114), .B1(new_n816_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n827_), .A2(new_n842_), .A3(new_n573_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n803_), .A2(new_n809_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(KEYINPUT58), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n615_), .B1(new_n844_), .B2(KEYINPUT58), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n833_), .A2(new_n839_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n789_), .B1(new_n849_), .B2(new_n632_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n682_), .A2(new_n415_), .A3(new_n643_), .A4(new_n661_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(G113gat), .B1(new_n852_), .B2(new_n477_), .ZN(new_n853_));
  XOR2_X1   g652(.A(new_n852_), .B(KEYINPUT59), .Z(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(G113gat), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n477_), .A2(KEYINPUT115), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(G113gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n853_), .B1(new_n855_), .B2(new_n859_), .ZN(G1340gat));
  OAI21_X1  g659(.A(G120gat), .B1(new_n854_), .B2(new_n585_), .ZN(new_n861_));
  INV_X1    g660(.A(G120gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n580_), .B2(KEYINPUT60), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n852_), .B(new_n863_), .C1(KEYINPUT60), .C2(new_n862_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n861_), .A2(new_n864_), .ZN(G1341gat));
  OAI21_X1  g664(.A(G127gat), .B1(new_n854_), .B2(new_n632_), .ZN(new_n866_));
  INV_X1    g665(.A(G127gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n852_), .A2(new_n867_), .A3(new_n633_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1342gat));
  OAI21_X1  g668(.A(G134gat), .B1(new_n854_), .B2(new_n615_), .ZN(new_n870_));
  INV_X1    g669(.A(G134gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n852_), .A2(new_n871_), .A3(new_n611_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(G1343gat));
  NAND4_X1  g672(.A1(new_n682_), .A2(new_n643_), .A3(new_n363_), .A4(new_n434_), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT116), .B1(new_n850_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876_));
  INV_X1    g675(.A(new_n874_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n837_), .A2(new_n838_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n633_), .B1(new_n878_), .B2(new_n833_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n876_), .B(new_n877_), .C1(new_n879_), .C2(new_n789_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n875_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n477_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT117), .B(G141gat), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1344gat));
  NAND2_X1  g683(.A1(new_n881_), .A2(new_n724_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n881_), .B2(new_n633_), .ZN(new_n888_));
  AOI211_X1 g687(.A(KEYINPUT118), .B(new_n632_), .C1(new_n875_), .C2(new_n880_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT61), .B(G155gat), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n888_), .A2(new_n889_), .A3(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT57), .B1(new_n837_), .B2(new_n727_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n838_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n803_), .A2(new_n809_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n841_), .A2(new_n843_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n895_), .A2(KEYINPUT58), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n681_), .ZN(new_n898_));
  OAI22_X1  g697(.A1(new_n832_), .A2(new_n894_), .B1(new_n898_), .B2(new_n845_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n632_), .B1(new_n893_), .B2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n789_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n876_), .B1(new_n902_), .B2(new_n877_), .ZN(new_n903_));
  AOI211_X1 g702(.A(KEYINPUT116), .B(new_n874_), .C1(new_n900_), .C2(new_n901_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n633_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT118), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n881_), .A2(new_n887_), .A3(new_n633_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n890_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n892_), .A2(new_n908_), .ZN(G1346gat));
  NOR2_X1   g708(.A1(new_n903_), .A2(new_n904_), .ZN(new_n910_));
  INV_X1    g709(.A(G162gat), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n910_), .A2(new_n911_), .A3(new_n615_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n910_), .B2(new_n727_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT119), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n915_), .B(new_n911_), .C1(new_n910_), .C2(new_n727_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n912_), .B1(new_n914_), .B2(new_n916_), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n682_), .A2(new_n309_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n918_), .A2(KEYINPUT120), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(KEYINPUT120), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n363_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n902_), .A2(new_n921_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n922_), .A2(new_n369_), .A3(new_n478_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n902_), .A2(new_n921_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n262_), .B1(new_n924_), .B2(new_n477_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n923_), .B1(new_n925_), .B2(KEYINPUT62), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n926_), .B1(KEYINPUT62), .B2(new_n925_), .ZN(G1348gat));
  NAND3_X1  g726(.A1(new_n924_), .A2(new_n263_), .A3(new_n581_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G176gat), .B1(new_n922_), .B2(new_n585_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT121), .ZN(G1349gat));
  NAND3_X1  g730(.A1(new_n924_), .A2(new_n375_), .A3(new_n633_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n252_), .B1(new_n922_), .B2(new_n632_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  XOR2_X1   g733(.A(new_n934_), .B(KEYINPUT122), .Z(G1350gat));
  NAND3_X1  g734(.A1(new_n924_), .A2(new_n376_), .A3(new_n611_), .ZN(new_n936_));
  OAI21_X1  g735(.A(G190gat), .B1(new_n922_), .B2(new_n615_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1351gat));
  NAND2_X1  g737(.A1(new_n434_), .A2(new_n409_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n850_), .A2(new_n432_), .A3(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n477_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n724_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n332_), .A2(KEYINPUT123), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n943_), .B(new_n944_), .ZN(G1353gat));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n946_));
  NAND2_X1  g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n940_), .A2(new_n633_), .A3(new_n947_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(KEYINPUT124), .ZN(new_n951_));
  INV_X1    g750(.A(new_n951_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n946_), .B1(new_n949_), .B2(new_n952_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n948_), .A2(KEYINPUT126), .A3(new_n951_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n949_), .A2(KEYINPUT125), .A3(new_n952_), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT125), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n956_), .B1(new_n948_), .B2(new_n951_), .ZN(new_n957_));
  AOI22_X1  g756(.A1(new_n953_), .A2(new_n954_), .B1(new_n955_), .B2(new_n957_), .ZN(G1354gat));
  AND3_X1   g757(.A1(new_n940_), .A2(G218gat), .A3(new_n681_), .ZN(new_n959_));
  AND2_X1   g758(.A1(new_n940_), .A2(new_n611_), .ZN(new_n960_));
  OR2_X1    g759(.A1(new_n960_), .A2(KEYINPUT127), .ZN(new_n961_));
  AOI21_X1  g760(.A(G218gat), .B1(new_n960_), .B2(KEYINPUT127), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n959_), .B1(new_n961_), .B2(new_n962_), .ZN(G1355gat));
endmodule


