//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n202_));
  NAND3_X1  g001(.A1(new_n202_), .A2(G183gat), .A3(G190gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT81), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G190gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT23), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n203_), .A2(KEYINPUT81), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT24), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  MUX2_X1   g012(.A(new_n212_), .B(KEYINPUT24), .S(new_n213_), .Z(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT26), .B(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT80), .B(G183gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n217_), .B1(new_n218_), .B2(KEYINPUT25), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n209_), .B(new_n214_), .C1(new_n216_), .C2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n207_), .A2(new_n203_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(G190gat), .B2(new_n218_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n210_), .A2(new_n211_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT22), .B(G169gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(new_n211_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(KEYINPUT82), .B(KEYINPUT30), .Z(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G127gat), .B(G134gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(G113gat), .ZN(new_n231_));
  INV_X1    g030(.A(G120gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n229_), .B(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n235_));
  NAND2_X1  g034(.A1(G227gat), .A2(G233gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G15gat), .B(G43gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(G71gat), .B(G99gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n237_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n234_), .B(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT18), .B(G64gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G92gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G8gat), .B(G36gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n245_), .B(new_n246_), .Z(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G226gat), .A2(G233gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n249_), .B(KEYINPUT92), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT19), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT93), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT20), .ZN(new_n254_));
  INV_X1    g053(.A(G204gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  OAI211_X1 g057(.A(KEYINPUT21), .B(new_n256_), .C1(new_n258_), .C2(KEYINPUT87), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n259_), .A2(KEYINPUT88), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(KEYINPUT88), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G211gat), .B(G218gat), .Z(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT89), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT21), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n257_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n264_), .A2(new_n265_), .A3(new_n257_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n209_), .B1(G183gat), .B2(G190gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n225_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT25), .B(G183gat), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n215_), .A2(new_n273_), .B1(new_n207_), .B2(new_n203_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n214_), .A2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n254_), .B1(new_n270_), .B2(new_n277_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n260_), .A2(new_n261_), .B1(new_n265_), .B2(new_n257_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n268_), .B1(new_n279_), .B2(new_n264_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n227_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n253_), .B1(new_n278_), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n251_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n267_), .A2(new_n269_), .A3(new_n276_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT20), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n248_), .B1(new_n283_), .B2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT20), .B1(new_n280_), .B2(new_n276_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n270_), .A2(new_n227_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n252_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n270_), .A2(new_n227_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n292_), .A2(KEYINPUT20), .A3(new_n251_), .A4(new_n285_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n247_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT94), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n288_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT27), .ZN(new_n297_));
  OAI211_X1 g096(.A(KEYINPUT94), .B(new_n248_), .C1(new_n283_), .C2(new_n287_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G78gat), .B(G106gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(G22gat), .B(G50gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT3), .ZN(new_n302_));
  INV_X1    g101(.A(G141gat), .ZN(new_n303_));
  INV_X1    g102(.A(G148gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n305_), .A2(new_n308_), .A3(new_n309_), .A4(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT85), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n318_));
  OR3_X1    g117(.A1(new_n312_), .A2(KEYINPUT84), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n313_), .B1(new_n312_), .B2(new_n318_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT84), .B1(new_n312_), .B2(new_n318_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n303_), .A2(new_n304_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n306_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n317_), .A2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n301_), .B1(new_n325_), .B2(KEYINPUT29), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n328_));
  INV_X1    g127(.A(new_n301_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n317_), .A2(new_n328_), .A3(new_n324_), .A4(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n326_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n327_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n300_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT91), .ZN(new_n335_));
  INV_X1    g134(.A(new_n333_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n335_), .B1(new_n336_), .B2(new_n331_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n334_), .B1(new_n337_), .B2(new_n300_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G228gat), .A2(G233gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n325_), .A2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n340_), .B1(new_n280_), .B2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n340_), .B1(new_n325_), .B2(KEYINPUT29), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n270_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n338_), .A2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n334_), .B(new_n346_), .C1(new_n337_), .C2(new_n300_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n289_), .A2(new_n290_), .A3(new_n252_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT98), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n286_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n285_), .A2(KEYINPUT98), .A3(KEYINPUT20), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n292_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n251_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n351_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(KEYINPUT27), .B(new_n294_), .C1(new_n357_), .C2(new_n247_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n299_), .A2(new_n350_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT99), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n299_), .A2(new_n350_), .A3(new_n358_), .A4(KEYINPUT99), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n243_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n325_), .A2(new_n233_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n325_), .A2(new_n233_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(KEYINPUT4), .A3(new_n365_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n365_), .A2(KEYINPUT4), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n366_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n364_), .A2(new_n368_), .A3(new_n365_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT0), .B(G57gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G85gat), .ZN(new_n374_));
  XOR2_X1   g173(.A(G1gat), .B(G29gat), .Z(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n370_), .A2(new_n371_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n350_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n299_), .A2(new_n381_), .A3(new_n358_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n296_), .A2(new_n298_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n364_), .A2(new_n365_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n376_), .B1(new_n385_), .B2(new_n368_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT96), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n366_), .A2(new_n368_), .A3(new_n367_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT96), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n389_), .B(new_n376_), .C1(new_n385_), .C2(new_n368_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n387_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT97), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT97), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n387_), .A2(new_n393_), .A3(new_n388_), .A4(new_n390_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n370_), .A2(KEYINPUT33), .A3(new_n371_), .A4(new_n378_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT95), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n379_), .A2(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n384_), .A2(new_n395_), .A3(new_n397_), .A4(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n283_), .A2(new_n287_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n247_), .A2(KEYINPUT32), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n377_), .A2(new_n379_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n286_), .A2(new_n352_), .B1(new_n227_), .B2(new_n270_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n251_), .B1(new_n404_), .B2(new_n354_), .ZN(new_n405_));
  OAI211_X1 g204(.A(KEYINPUT32), .B(new_n247_), .C1(new_n405_), .C2(new_n351_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n403_), .A2(new_n406_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n382_), .A2(new_n383_), .B1(new_n400_), .B2(new_n407_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n363_), .A2(new_n381_), .B1(new_n408_), .B2(new_n243_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G15gat), .B(G22gat), .ZN(new_n410_));
  INV_X1    g209(.A(G1gat), .ZN(new_n411_));
  INV_X1    g210(.A(G8gat), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT14), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G8gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G231gat), .A2(G233gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  OR2_X1    g217(.A1(G57gat), .A2(G64gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G57gat), .A2(G64gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT11), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G71gat), .B(G78gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT11), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n419_), .A2(new_n425_), .A3(new_n420_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n421_), .A2(new_n423_), .A3(KEYINPUT11), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n418_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G127gat), .B(G155gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G183gat), .B(G211gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(KEYINPUT75), .A3(KEYINPUT17), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(KEYINPUT17), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT75), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n431_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n441_), .B(KEYINPUT76), .Z(new_n442_));
  AOI21_X1  g241(.A(new_n431_), .B1(KEYINPUT17), .B2(new_n436_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n443_), .B1(KEYINPUT17), .B2(new_n436_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(G29gat), .A2(G36gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G29gat), .A2(G36gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(G43gat), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G29gat), .ZN(new_n450_));
  INV_X1    g249(.A(G36gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G43gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G29gat), .A2(G36gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n449_), .A2(new_n455_), .A3(G50gat), .ZN(new_n456_));
  AOI21_X1  g255(.A(G50gat), .B1(new_n449_), .B2(new_n455_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT70), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G50gat), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n447_), .A2(new_n448_), .A3(G43gat), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n453_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT70), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n449_), .A2(new_n455_), .A3(G50gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT15), .B1(new_n458_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n458_), .A2(new_n465_), .A3(KEYINPUT15), .ZN(new_n468_));
  XOR2_X1   g267(.A(KEYINPUT10), .B(G99gat), .Z(new_n469_));
  INV_X1    g268(.A(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G92gat), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n472_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT65), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n474_), .A2(G92gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(G85gat), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n472_), .A2(G85gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n472_), .A2(G85gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT9), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n471_), .A2(new_n476_), .A3(new_n479_), .A4(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI22_X1  g287(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n488_), .A2(new_n482_), .A3(new_n483_), .A4(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT8), .ZN(new_n491_));
  XOR2_X1   g290(.A(G85gat), .B(G92gat), .Z(new_n492_));
  AND3_X1   g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n491_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n485_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT67), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  OAI211_X1 g296(.A(KEYINPUT67), .B(new_n485_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n467_), .A2(new_n468_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G232gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT69), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT34), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT35), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n462_), .A2(new_n464_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n504_), .B1(new_n495_), .B2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n499_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT71), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n502_), .A2(new_n503_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G190gat), .B(G218gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(G134gat), .ZN(new_n512_));
  INV_X1    g311(.A(G162gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n515_), .A2(KEYINPUT36), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n509_), .A2(new_n508_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT71), .B1(new_n502_), .B2(new_n503_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n518_), .B(new_n519_), .C1(new_n499_), .C2(new_n506_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(KEYINPUT36), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n510_), .A2(new_n517_), .A3(new_n520_), .A4(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n510_), .A2(new_n520_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n516_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT72), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT72), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n524_), .A2(new_n527_), .A3(new_n516_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n523_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(KEYINPUT73), .A3(KEYINPUT37), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT37), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n527_), .B1(new_n524_), .B2(new_n516_), .ZN(new_n532_));
  AOI211_X1 g331(.A(KEYINPUT72), .B(new_n517_), .C1(new_n510_), .C2(new_n520_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n522_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT73), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n531_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n409_), .A2(new_n446_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT77), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n539_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n462_), .A2(KEYINPUT77), .A3(new_n464_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n540_), .A2(new_n416_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n416_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n468_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n416_), .B1(new_n547_), .B2(new_n466_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n540_), .A2(new_n541_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n416_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n545_), .B(KEYINPUT78), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G113gat), .B(G141gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(new_n210_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(G197gat), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n546_), .A2(new_n553_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n546_), .B2(new_n553_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n561_), .A2(KEYINPUT79), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(KEYINPUT79), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n430_), .A2(KEYINPUT12), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n490_), .A2(new_n492_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT8), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT67), .B1(new_n571_), .B2(new_n485_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n498_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n567_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT12), .B1(new_n495_), .B2(new_n430_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n429_), .B(new_n485_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT64), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n574_), .A2(new_n578_), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n429_), .B1(new_n571_), .B2(new_n485_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n580_), .B1(new_n577_), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G120gat), .B(G148gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(new_n255_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT5), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(G176gat), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(G176gat), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n582_), .A2(new_n584_), .A3(new_n588_), .A4(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n582_), .A2(new_n584_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n587_), .B(G176gat), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT68), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n589_), .A2(KEYINPUT68), .A3(new_n588_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n590_), .B1(new_n591_), .B2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT13), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n565_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n538_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n411_), .A3(new_n380_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT38), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n409_), .A2(new_n529_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n599_), .A2(new_n561_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n445_), .A3(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G1gat), .B1(new_n606_), .B2(new_n381_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n607_), .ZN(G1324gat));
  NAND2_X1  g407(.A1(new_n299_), .A2(new_n358_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n601_), .A2(new_n412_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n609_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G8gat), .B1(new_n606_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT39), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT101), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n612_), .A2(new_n618_), .A3(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT40), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(new_n619_), .A3(KEYINPUT40), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(G1325gat));
  OAI21_X1  g423(.A(G15gat), .B1(new_n606_), .B2(new_n243_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT41), .Z(new_n626_));
  INV_X1    g425(.A(G15gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n601_), .A2(new_n627_), .A3(new_n242_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1326gat));
  OAI21_X1  g428(.A(G22gat), .B1(new_n606_), .B2(new_n350_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT42), .ZN(new_n631_));
  INV_X1    g430(.A(G22gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n601_), .A2(new_n632_), .A3(new_n382_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(G1327gat));
  INV_X1    g433(.A(KEYINPUT43), .ZN(new_n635_));
  INV_X1    g434(.A(new_n537_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n409_), .B2(KEYINPUT102), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n361_), .A2(new_n362_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n381_), .A3(new_n242_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n408_), .A2(new_n243_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n635_), .B1(new_n637_), .B2(new_n643_), .ZN(new_n644_));
  AOI211_X1 g443(.A(new_n380_), .B(new_n243_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n383_), .A2(new_n382_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n400_), .A2(new_n407_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n646_), .A2(new_n647_), .A3(new_n243_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n635_), .B(new_n537_), .C1(new_n645_), .C2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT103), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n641_), .A2(new_n651_), .A3(new_n635_), .A4(new_n537_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n446_), .B(new_n605_), .C1(new_n644_), .C2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n639_), .A2(KEYINPUT102), .A3(new_n640_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n537_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n409_), .A2(KEYINPUT102), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT43), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n650_), .A3(new_n652_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n446_), .A4(new_n605_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n656_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n663_), .A2(G29gat), .A3(new_n380_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n641_), .A2(new_n446_), .A3(new_n529_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n600_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n450_), .B1(new_n668_), .B2(new_n381_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n664_), .A2(new_n669_), .ZN(G1328gat));
  NAND3_X1  g469(.A1(new_n667_), .A2(new_n451_), .A3(new_n609_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT45), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n656_), .A2(new_n609_), .A3(new_n662_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n673_), .A2(new_n674_), .A3(G36gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n673_), .B2(G36gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(KEYINPUT46), .B(new_n672_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1329gat));
  NOR3_X1   g480(.A1(new_n668_), .A2(G43gat), .A3(new_n243_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n663_), .A2(new_n242_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n683_), .B2(G43gat), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  AOI211_X1 g485(.A(KEYINPUT47), .B(new_n682_), .C1(new_n683_), .C2(G43gat), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1330gat));
  AOI21_X1  g487(.A(G50gat), .B1(new_n667_), .B2(new_n382_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n350_), .A2(new_n459_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n663_), .B2(new_n690_), .ZN(G1331gat));
  INV_X1    g490(.A(new_n561_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n598_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n538_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G57gat), .B1(new_n695_), .B2(new_n380_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G57gat), .B1(new_n381_), .B2(KEYINPUT105), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n604_), .A2(new_n445_), .A3(new_n599_), .A4(new_n565_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(KEYINPUT105), .A2(G57gat), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n696_), .B1(new_n697_), .B2(new_n700_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT106), .Z(G1332gat));
  OAI21_X1  g501(.A(G64gat), .B1(new_n698_), .B2(new_n613_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT48), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n613_), .A2(G64gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n694_), .B2(new_n705_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT107), .Z(G1333gat));
  OAI21_X1  g506(.A(G71gat), .B1(new_n698_), .B2(new_n243_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT49), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n243_), .A2(G71gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n694_), .B2(new_n710_), .ZN(G1334gat));
  OAI21_X1  g510(.A(G78gat), .B1(new_n698_), .B2(new_n350_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT50), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n350_), .A2(G78gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n694_), .B2(new_n714_), .ZN(G1335gat));
  INV_X1    g514(.A(new_n693_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n665_), .A2(new_n716_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n717_), .A2(KEYINPUT108), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(KEYINPUT108), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n720_), .A2(G85gat), .A3(new_n381_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n661_), .A2(new_n446_), .A3(new_n693_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n380_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n721_), .B1(new_n724_), .B2(G85gat), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT109), .ZN(G1336gat));
  INV_X1    g525(.A(new_n720_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G92gat), .B1(new_n727_), .B2(new_n609_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n475_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n474_), .A2(G92gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n613_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n728_), .B1(new_n723_), .B2(new_n731_), .ZN(G1337gat));
  NAND3_X1  g531(.A1(new_n727_), .A2(new_n242_), .A3(new_n469_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G99gat), .B1(new_n722_), .B2(new_n243_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g535(.A(G106gat), .B1(new_n722_), .B2(new_n350_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT52), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n470_), .B(new_n382_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT110), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT53), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n738_), .A2(new_n743_), .A3(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1339gat));
  NAND2_X1  g544(.A1(new_n363_), .A2(new_n380_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT117), .ZN(new_n747_));
  INV_X1    g546(.A(new_n596_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n576_), .B1(new_n583_), .B2(KEYINPUT12), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n566_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n580_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n580_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(KEYINPUT55), .B2(new_n752_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n574_), .A2(new_n578_), .A3(KEYINPUT55), .A4(new_n581_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n748_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n581_), .B1(new_n574_), .B2(new_n578_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n582_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n754_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(KEYINPUT56), .A3(new_n748_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n758_), .A2(new_n759_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766_));
  INV_X1    g565(.A(new_n552_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n540_), .A2(new_n416_), .A3(new_n541_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n551_), .B2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n766_), .B1(new_n769_), .B2(new_n557_), .ZN(new_n770_));
  OAI211_X1 g569(.A(KEYINPUT112), .B(new_n556_), .C1(new_n544_), .C2(new_n767_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n548_), .A2(new_n551_), .A3(new_n767_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .A4(KEYINPUT113), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n775_), .A2(new_n558_), .A3(new_n590_), .A4(new_n776_), .ZN(new_n777_));
  AOI211_X1 g576(.A(new_n757_), .B(new_n596_), .C1(new_n762_), .C2(new_n754_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(KEYINPUT114), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n765_), .A2(KEYINPUT115), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT58), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT115), .B1(new_n765_), .B2(new_n779_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT116), .B(new_n537_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT56), .B1(new_n763_), .B2(new_n748_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n787_), .A2(new_n778_), .A3(KEYINPUT114), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n775_), .A2(new_n558_), .A3(new_n776_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n789_), .B(new_n590_), .C1(new_n764_), .C2(new_n759_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(new_n781_), .A3(new_n780_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT116), .B1(new_n792_), .B2(new_n537_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n788_), .A2(new_n790_), .A3(new_n781_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n785_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n692_), .B(new_n590_), .C1(new_n787_), .C2(new_n778_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n789_), .A2(new_n597_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n798_), .A2(KEYINPUT57), .A3(new_n534_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT57), .B1(new_n798_), .B2(new_n534_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n747_), .B1(new_n795_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n537_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n794_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n784_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(KEYINPUT117), .A3(new_n801_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n803_), .A2(new_n446_), .A3(new_n809_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n446_), .A2(new_n599_), .A3(new_n564_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT111), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(new_n537_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n746_), .B1(new_n810_), .B2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G113gat), .B1(new_n816_), .B2(new_n692_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n813_), .B(KEYINPUT54), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n445_), .B1(new_n808_), .B2(new_n801_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n820_), .A2(KEYINPUT59), .A3(new_n746_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n746_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n808_), .A2(KEYINPUT117), .A3(new_n801_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT117), .B1(new_n808_), .B2(new_n801_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n445_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n822_), .B1(new_n825_), .B2(new_n818_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(KEYINPUT118), .A3(KEYINPUT59), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n816_), .B2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n821_), .B1(new_n827_), .B2(new_n830_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n831_), .A2(new_n564_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n817_), .B1(new_n832_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n232_), .B1(new_n831_), .B2(new_n599_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n232_), .B1(new_n598_), .B2(KEYINPUT60), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n232_), .A2(KEYINPUT60), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n816_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n834_), .B1(new_n835_), .B2(new_n839_), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n598_), .B(new_n821_), .C1(new_n827_), .C2(new_n830_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT119), .B(new_n838_), .C1(new_n841_), .C2(new_n232_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1341gat));
  AOI21_X1  g642(.A(G127gat), .B1(new_n816_), .B2(new_n445_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n445_), .A2(G127gat), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(KEYINPUT120), .Z(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n831_), .B2(new_n846_), .ZN(G1342gat));
  AOI21_X1  g646(.A(G134gat), .B1(new_n816_), .B2(new_n529_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n537_), .A2(G134gat), .ZN(new_n849_));
  XOR2_X1   g648(.A(new_n849_), .B(KEYINPUT121), .Z(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n831_), .B2(new_n850_), .ZN(G1343gat));
  AOI21_X1  g650(.A(new_n609_), .B1(new_n810_), .B2(new_n815_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n350_), .A2(new_n381_), .A3(new_n242_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n561_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n303_), .ZN(G1344gat));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n598_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(new_n304_), .ZN(G1345gat));
  NOR2_X1   g657(.A1(new_n854_), .A2(new_n446_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT61), .B(G155gat), .Z(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1346gat));
  NOR3_X1   g660(.A1(new_n854_), .A2(new_n513_), .A3(new_n636_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n852_), .A2(new_n529_), .A3(new_n853_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n513_), .B2(new_n863_), .ZN(G1347gat));
  NOR2_X1   g663(.A1(new_n613_), .A2(new_n380_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n242_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n820_), .A2(new_n382_), .A3(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G169gat), .B1(new_n868_), .B2(new_n561_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n869_), .A2(KEYINPUT62), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(KEYINPUT62), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n692_), .A2(new_n224_), .ZN(new_n872_));
  XOR2_X1   g671(.A(new_n872_), .B(KEYINPUT122), .Z(new_n873_));
  OAI22_X1  g672(.A1(new_n870_), .A2(new_n871_), .B1(new_n868_), .B2(new_n873_), .ZN(G1348gat));
  AOI21_X1  g673(.A(G176gat), .B1(new_n867_), .B2(new_n599_), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT123), .Z(new_n876_));
  NAND2_X1  g675(.A1(new_n810_), .A2(new_n815_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n350_), .ZN(new_n878_));
  NOR4_X1   g677(.A1(new_n878_), .A2(new_n211_), .A3(new_n598_), .A4(new_n866_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n876_), .A2(new_n879_), .ZN(G1349gat));
  NAND2_X1  g679(.A1(new_n867_), .A2(new_n445_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n218_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n273_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n881_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(KEYINPUT124), .ZN(G1350gat));
  NAND3_X1  g684(.A1(new_n867_), .A2(new_n215_), .A3(new_n529_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n867_), .A2(new_n537_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n886_), .B1(new_n888_), .B2(new_n206_), .ZN(G1351gat));
  NOR2_X1   g688(.A1(new_n350_), .A2(new_n242_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n877_), .A2(new_n890_), .A3(new_n865_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n692_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT126), .B1(new_n895_), .B2(new_n255_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(KEYINPUT126), .B2(new_n255_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n891_), .A2(new_n598_), .ZN(new_n898_));
  MUX2_X1   g697(.A(new_n896_), .B(new_n897_), .S(new_n898_), .Z(G1353gat));
  NAND2_X1  g698(.A1(new_n892_), .A2(new_n445_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  AND2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n900_), .B2(new_n901_), .ZN(G1354gat));
  OR3_X1    g703(.A1(new_n891_), .A2(G218gat), .A3(new_n534_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G218gat), .B1(new_n891_), .B2(new_n636_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


