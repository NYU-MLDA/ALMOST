//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n204_));
  OAI22_X1  g003(.A1(new_n204_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT7), .ZN(new_n206_));
  INV_X1    g005(.A(G99gat), .ZN(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND4_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .A4(KEYINPUT64), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n203_), .A2(new_n205_), .A3(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G85gat), .B(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT8), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n211_), .ZN(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT10), .B(G99gat), .Z(new_n219_));
  AOI22_X1  g018(.A1(new_n218_), .A2(KEYINPUT9), .B1(new_n219_), .B2(new_n208_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n220_), .B(new_n203_), .C1(KEYINPUT9), .C2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G57gat), .B(G64gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT66), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n225_), .A2(KEYINPUT11), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(KEYINPUT11), .ZN(new_n227_));
  XOR2_X1   g026(.A(G71gat), .B(G78gat), .Z(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n227_), .A2(new_n228_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n231_), .A2(KEYINPUT68), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT12), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(new_n231_), .B2(KEYINPUT68), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n223_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G230gat), .A2(G233gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n215_), .A2(new_n222_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n231_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n231_), .A2(new_n237_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n238_), .B1(new_n233_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n235_), .A2(new_n236_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n239_), .ZN(new_n242_));
  OAI211_X1 g041(.A(G230gat), .B(G233gat), .C1(new_n242_), .C2(new_n238_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G120gat), .B(G148gat), .Z(new_n245_));
  XNOR2_X1  g044(.A(G176gat), .B(G204gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n244_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n241_), .A2(new_n243_), .A3(new_n249_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n254_), .A2(KEYINPUT13), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(KEYINPUT13), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G15gat), .B(G22gat), .ZN(new_n258_));
  INV_X1    g057(.A(G1gat), .ZN(new_n259_));
  INV_X1    g058(.A(G8gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT14), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G1gat), .B(G8gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n262_), .B(new_n263_), .Z(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G29gat), .B(G36gat), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n266_), .A2(KEYINPUT71), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(KEYINPUT71), .ZN(new_n268_));
  XOR2_X1   g067(.A(G43gat), .B(G50gat), .Z(new_n269_));
  OR3_X1    g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n269_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n265_), .B(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G229gat), .A2(G233gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n272_), .B(KEYINPUT15), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n265_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT75), .ZN(new_n278_));
  INV_X1    g077(.A(new_n274_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n272_), .B2(new_n264_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n275_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G113gat), .B(G141gat), .Z(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT77), .ZN(new_n283_));
  XOR2_X1   g082(.A(G169gat), .B(G197gat), .Z(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT76), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n281_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n231_), .B(new_n264_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G231gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G127gat), .B(G155gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT16), .ZN(new_n295_));
  XOR2_X1   g094(.A(G183gat), .B(G211gat), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT17), .ZN(new_n298_));
  OR3_X1    g097(.A1(new_n297_), .A2(KEYINPUT68), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n293_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n297_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(KEYINPUT17), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n292_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n257_), .A2(new_n289_), .A3(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n305_), .B(KEYINPUT100), .Z(new_n306_));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G127gat), .B(G134gat), .Z(new_n309_));
  XOR2_X1   g108(.A(G113gat), .B(G120gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT87), .ZN(new_n313_));
  NOR2_X1   g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  OAI211_X1 g115(.A(KEYINPUT87), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(KEYINPUT86), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT86), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(G141gat), .B2(G148gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n315_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G141gat), .A2(G148gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT2), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n318_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n314_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n323_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n326_), .B1(KEYINPUT1), .B2(new_n328_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n328_), .A2(KEYINPUT1), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n312_), .B(KEYINPUT96), .C1(new_n330_), .C2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n335_), .B1(new_n325_), .B2(new_n329_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(new_n338_), .B2(new_n311_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n338_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n341_), .A2(KEYINPUT96), .A3(new_n337_), .A4(new_n312_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n308_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(G85gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT0), .B(G57gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n346_), .B(new_n347_), .Z(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n341_), .A2(new_n312_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n338_), .A2(new_n311_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n308_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n344_), .A2(new_n349_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n336_), .A2(new_n339_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n307_), .B1(new_n355_), .B2(new_n342_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n348_), .B1(new_n356_), .B2(new_n352_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n357_), .A3(KEYINPUT98), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT98), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n359_), .B(new_n348_), .C1(new_n356_), .C2(new_n352_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G8gat), .B(G36gat), .Z(new_n362_));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT19), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G169gat), .A2(G176gat), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n371_), .A2(KEYINPUT79), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(KEYINPUT79), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G176gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT22), .B(G169gat), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n374_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT93), .ZN(new_n378_));
  INV_X1    g177(.A(G183gat), .ZN(new_n379_));
  INV_X1    g178(.A(G190gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT23), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n381_), .A2(KEYINPUT80), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(KEYINPUT80), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n379_), .A2(new_n380_), .A3(KEYINPUT23), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(G183gat), .A2(G190gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n378_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n385_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n391_), .A2(KEYINPUT93), .A3(new_n388_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n377_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n386_), .A2(new_n381_), .ZN(new_n394_));
  INV_X1    g193(.A(G169gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n375_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n396_), .A2(KEYINPUT24), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT25), .B(G183gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT26), .B(G190gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(KEYINPUT24), .A3(new_n371_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n394_), .A2(new_n397_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n393_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G204gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT90), .B1(new_n404_), .B2(G197gat), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT90), .ZN(new_n406_));
  INV_X1    g205(.A(G197gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(G204gat), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n405_), .A2(new_n408_), .B1(G197gat), .B2(new_n404_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT21), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT89), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n407_), .B2(G204gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n404_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n407_), .A2(G204gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT21), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G211gat), .B(G218gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n411_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT91), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n418_), .A2(new_n410_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n409_), .B2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT20), .B(new_n370_), .C1(new_n403_), .C2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT81), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT22), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n425_), .B1(new_n426_), .B2(G169gat), .ZN(new_n427_));
  AOI21_X1  g226(.A(G176gat), .B1(new_n426_), .B2(G169gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n395_), .A2(KEYINPUT81), .A3(KEYINPUT22), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT82), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n427_), .A2(new_n428_), .A3(new_n432_), .A4(new_n429_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n374_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n388_), .B1(new_n386_), .B2(new_n381_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n374_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n439_), .B1(new_n440_), .B2(KEYINPUT83), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT25), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT78), .B1(new_n443_), .B2(G183gat), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n444_), .B(new_n399_), .C1(new_n398_), .C2(KEYINPUT78), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n372_), .A2(KEYINPUT24), .A3(new_n373_), .A4(new_n396_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(new_n397_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n447_), .A2(new_n391_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT84), .B1(new_n442_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n451_));
  AOI211_X1 g250(.A(new_n451_), .B(new_n448_), .C1(new_n438_), .C2(new_n441_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n423_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT94), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n434_), .A2(KEYINPUT83), .A3(new_n435_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n439_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n440_), .A2(KEYINPUT83), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n449_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n451_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n442_), .A2(KEYINPUT84), .A3(new_n449_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(KEYINPUT94), .A3(new_n423_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n424_), .B1(new_n455_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n466_), .B1(new_n403_), .B2(new_n423_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n422_), .A2(new_n409_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n419_), .A2(new_n420_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n419_), .A2(new_n420_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n461_), .A2(new_n462_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n370_), .B1(new_n467_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n367_), .B1(new_n465_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n424_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT94), .B1(new_n463_), .B2(new_n423_), .ZN(new_n476_));
  AOI211_X1 g275(.A(new_n454_), .B(new_n471_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n473_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(new_n366_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n474_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT27), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n467_), .A2(new_n472_), .A3(new_n370_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT20), .B1(new_n403_), .B2(new_n423_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n487_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n485_), .B1(new_n488_), .B2(new_n369_), .ZN(new_n489_));
  OAI211_X1 g288(.A(KEYINPUT27), .B(new_n480_), .C1(new_n489_), .C2(new_n366_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n483_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G71gat), .B(G99gat), .ZN(new_n492_));
  INV_X1    g291(.A(G43gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G227gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(G15gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT30), .ZN(new_n499_));
  INV_X1    g298(.A(new_n494_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n461_), .A2(new_n462_), .A3(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n495_), .A2(new_n499_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n499_), .B1(new_n495_), .B2(new_n501_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT31), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n495_), .A2(new_n501_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n499_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT31), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(new_n502_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n505_), .A2(new_n312_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n312_), .B1(new_n505_), .B2(new_n510_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n341_), .A2(KEYINPUT29), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n423_), .A2(KEYINPUT88), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G228gat), .A2(G233gat), .ZN(new_n516_));
  INV_X1    g315(.A(G78gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(G106gat), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n519_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OR3_X1    g321(.A1(new_n341_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT28), .B1(new_n341_), .B2(KEYINPUT29), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G22gat), .B(G50gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n523_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n528_), .A2(KEYINPUT92), .A3(new_n529_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n522_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n520_), .A2(new_n531_), .A3(new_n530_), .A4(new_n521_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NOR4_X1   g336(.A1(new_n491_), .A2(new_n513_), .A3(new_n361_), .A4(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n488_), .A2(new_n369_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n484_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n367_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n480_), .A2(KEYINPUT27), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n541_), .A2(new_n542_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n536_), .A2(new_n361_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n340_), .A2(new_n343_), .A3(new_n308_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n350_), .A2(new_n308_), .A3(new_n351_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n546_), .A2(new_n349_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n547_), .B2(KEYINPUT97), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n547_), .A2(KEYINPUT97), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n357_), .A2(KEYINPUT33), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT33), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n551_), .B(new_n348_), .C1(new_n356_), .C2(new_n352_), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n548_), .A2(new_n549_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n474_), .A2(new_n480_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n366_), .A2(KEYINPUT32), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n555_), .B1(new_n539_), .B2(new_n484_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n478_), .A2(new_n479_), .A3(new_n555_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n361_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n554_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n543_), .A2(new_n544_), .B1(new_n559_), .B2(new_n536_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT85), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n561_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n503_), .A2(new_n504_), .A3(KEYINPUT31), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n509_), .B1(new_n508_), .B2(new_n502_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n311_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n505_), .A2(new_n312_), .A3(new_n510_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(KEYINPUT85), .A3(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT99), .B1(new_n560_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n559_), .A2(new_n536_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n483_), .A2(new_n490_), .A3(new_n544_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT99), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n562_), .A2(new_n567_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n538_), .B1(new_n569_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT72), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT36), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT36), .ZN(new_n583_));
  INV_X1    g382(.A(new_n237_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT35), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n584_), .A2(new_n272_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n217_), .A2(new_n222_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n276_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n590_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n589_), .A2(new_n585_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI221_X1 g394(.A(new_n590_), .B1(new_n585_), .B2(new_n589_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n583_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n595_), .A2(new_n596_), .ZN(new_n598_));
  OAI221_X1 g397(.A(new_n582_), .B1(new_n597_), .B2(new_n581_), .C1(KEYINPUT73), .C2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n582_), .B1(new_n597_), .B2(new_n581_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n598_), .A2(KEYINPUT73), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n576_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n306_), .A2(new_n361_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(G1gat), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT101), .Z(new_n607_));
  NOR2_X1   g406(.A1(new_n576_), .A2(new_n288_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n599_), .A2(new_n602_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT74), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT37), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(KEYINPUT37), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n609_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n599_), .A2(new_n610_), .A3(new_n602_), .A4(KEYINPUT37), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n613_), .A2(new_n257_), .A3(new_n304_), .A4(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n608_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n259_), .A3(new_n361_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT38), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n607_), .A2(new_n620_), .ZN(G1324gat));
  NAND3_X1  g420(.A1(new_n618_), .A2(new_n260_), .A3(new_n491_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n306_), .A2(new_n491_), .A3(new_n604_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(G8gat), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n624_), .A2(KEYINPUT39), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(KEYINPUT39), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n622_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n627_), .B(new_n628_), .Z(G1325gat));
  NAND3_X1  g428(.A1(new_n618_), .A2(new_n497_), .A3(new_n568_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n306_), .A2(new_n568_), .A3(new_n604_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n631_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT41), .B1(new_n631_), .B2(G15gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n630_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT103), .Z(G1326gat));
  NAND3_X1  g434(.A1(new_n306_), .A2(new_n537_), .A3(new_n604_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(G22gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT42), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n536_), .A2(G22gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n617_), .B2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT104), .ZN(G1327gat));
  INV_X1    g440(.A(new_n257_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n304_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n603_), .A2(new_n643_), .ZN(new_n644_));
  NOR4_X1   g443(.A1(new_n576_), .A2(new_n288_), .A3(new_n642_), .A4(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(G29gat), .B1(new_n645_), .B2(new_n361_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n613_), .A2(new_n614_), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT43), .B1(new_n576_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n538_), .ZN(new_n649_));
  AOI221_X4 g448(.A(KEYINPUT99), .B1(new_n562_), .B2(new_n567_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n573_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n613_), .A2(new_n614_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n648_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n257_), .A2(new_n289_), .A3(new_n643_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT44), .B1(new_n656_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  AOI211_X1 g459(.A(new_n660_), .B(new_n657_), .C1(new_n648_), .C2(new_n655_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n361_), .A2(G29gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n646_), .B1(new_n662_), .B2(new_n663_), .ZN(G1328gat));
  NOR2_X1   g463(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT107), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n659_), .A2(new_n661_), .A3(new_n543_), .ZN(new_n668_));
  INV_X1    g467(.A(G36gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n667_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n648_), .A2(new_n655_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n660_), .B1(new_n671_), .B2(new_n657_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n656_), .A2(KEYINPUT44), .A3(new_n658_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n491_), .A3(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n674_), .A2(KEYINPUT105), .A3(G36gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n670_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n645_), .A2(new_n669_), .A3(new_n491_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT45), .Z(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n666_), .B1(new_n676_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n666_), .ZN(new_n681_));
  AOI211_X1 g480(.A(new_n681_), .B(new_n678_), .C1(new_n670_), .C2(new_n675_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n680_), .A2(new_n682_), .ZN(G1329gat));
  AOI21_X1  g482(.A(G43gat), .B1(new_n645_), .B2(new_n568_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n513_), .A2(new_n493_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n662_), .B2(new_n685_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g486(.A(G50gat), .B1(new_n645_), .B2(new_n537_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n537_), .A2(G50gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n662_), .B2(new_n689_), .ZN(G1331gat));
  NOR2_X1   g489(.A1(new_n257_), .A2(new_n289_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n576_), .A2(new_n692_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n613_), .A2(new_n304_), .A3(new_n614_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G57gat), .B1(new_n696_), .B2(new_n361_), .ZN(new_n697_));
  NOR4_X1   g496(.A1(new_n576_), .A2(new_n692_), .A3(new_n603_), .A4(new_n643_), .ZN(new_n698_));
  INV_X1    g497(.A(G57gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n361_), .B2(KEYINPUT108), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(KEYINPUT108), .B2(new_n699_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n697_), .B1(new_n698_), .B2(new_n701_), .ZN(G1332gat));
  INV_X1    g501(.A(G64gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n698_), .B2(new_n491_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT48), .Z(new_n705_));
  NAND3_X1  g504(.A1(new_n696_), .A2(new_n703_), .A3(new_n491_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1333gat));
  INV_X1    g506(.A(G71gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n698_), .B2(new_n568_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT49), .Z(new_n710_));
  NAND3_X1  g509(.A1(new_n696_), .A2(new_n708_), .A3(new_n568_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1334gat));
  AOI21_X1  g511(.A(new_n517_), .B1(new_n698_), .B2(new_n537_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT50), .Z(new_n714_));
  NOR2_X1   g513(.A1(new_n536_), .A2(G78gat), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT109), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n714_), .B1(new_n695_), .B2(new_n716_), .ZN(G1335gat));
  NAND2_X1  g516(.A1(new_n671_), .A2(KEYINPUT111), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n656_), .A2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n692_), .A2(new_n304_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n718_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(G85gat), .A3(new_n361_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n644_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n693_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G85gat), .B1(new_n726_), .B2(new_n361_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT110), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n723_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(G1336gat));
  INV_X1    g530(.A(G92gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n726_), .A2(new_n732_), .A3(new_n491_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n722_), .A2(new_n491_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n732_), .ZN(G1337gat));
  NAND4_X1  g534(.A1(new_n718_), .A2(new_n568_), .A3(new_n720_), .A4(new_n721_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G99gat), .ZN(new_n737_));
  INV_X1    g536(.A(new_n513_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n693_), .A2(new_n738_), .A3(new_n219_), .A4(new_n724_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT113), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n741_), .A2(KEYINPUT115), .A3(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(KEYINPUT51), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n745_));
  INV_X1    g544(.A(new_n740_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(G99gat), .B2(new_n736_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n742_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n743_), .B1(new_n744_), .B2(new_n749_), .ZN(G1338gat));
  AND3_X1   g549(.A1(new_n656_), .A2(new_n537_), .A3(new_n721_), .ZN(new_n751_));
  OR3_X1    g550(.A1(new_n751_), .A2(KEYINPUT116), .A3(new_n208_), .ZN(new_n752_));
  OAI21_X1  g551(.A(KEYINPUT116), .B1(new_n751_), .B2(new_n208_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(KEYINPUT52), .A3(new_n753_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n753_), .A2(KEYINPUT52), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n726_), .A2(new_n208_), .A3(new_n537_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n754_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT53), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n754_), .A2(new_n755_), .A3(new_n759_), .A4(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1339gat));
  NAND4_X1  g560(.A1(new_n235_), .A2(KEYINPUT55), .A3(new_n236_), .A4(new_n240_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT117), .B1(new_n241_), .B2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n236_), .B1(new_n235_), .B2(new_n240_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n241_), .A2(KEYINPUT117), .A3(new_n765_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n764_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n250_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT56), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(new_n773_), .A3(new_n250_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n274_), .B1(new_n272_), .B2(new_n264_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n278_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n273_), .A2(new_n279_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n285_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(new_n281_), .B2(new_n285_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(new_n252_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n772_), .A2(new_n774_), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n782_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(new_n654_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT120), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n773_), .A2(KEYINPUT119), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n771_), .A2(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n289_), .A2(new_n252_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n770_), .A2(KEYINPUT119), .A3(new_n773_), .A4(new_n250_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n779_), .A2(new_n253_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n603_), .B1(KEYINPUT121), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n794_), .A2(KEYINPUT121), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n797_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n793_), .A2(new_n795_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n783_), .A2(new_n802_), .A3(new_n654_), .A4(new_n784_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n786_), .A2(new_n801_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n643_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n694_), .A2(new_n806_), .A3(new_n288_), .A4(new_n257_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT54), .B1(new_n615_), .B2(new_n289_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n805_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n361_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n491_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n814_), .A2(new_n537_), .A3(new_n513_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n811_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT59), .ZN(new_n817_));
  INV_X1    g616(.A(new_n800_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n799_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n785_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n809_), .B1(new_n820_), .B2(new_n643_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT59), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n815_), .A2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT122), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  OR3_X1    g623(.A1(new_n821_), .A2(KEYINPUT122), .A3(new_n823_), .ZN(new_n825_));
  INV_X1    g624(.A(G113gat), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n288_), .A2(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT123), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n817_), .A2(new_n824_), .A3(new_n825_), .A4(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n826_), .B1(new_n816_), .B2(new_n288_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1340gat));
  NAND4_X1  g630(.A1(new_n817_), .A2(new_n824_), .A3(new_n825_), .A4(new_n642_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(G120gat), .ZN(new_n833_));
  INV_X1    g632(.A(new_n816_), .ZN(new_n834_));
  INV_X1    g633(.A(G120gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n257_), .B2(KEYINPUT60), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n834_), .B(new_n836_), .C1(KEYINPUT60), .C2(new_n835_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n833_), .A2(new_n837_), .ZN(G1341gat));
  NAND4_X1  g637(.A1(new_n817_), .A2(new_n824_), .A3(new_n825_), .A4(new_n304_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(G127gat), .ZN(new_n840_));
  OR3_X1    g639(.A1(new_n816_), .A2(G127gat), .A3(new_n643_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1342gat));
  NAND4_X1  g641(.A1(new_n817_), .A2(new_n824_), .A3(new_n825_), .A4(new_n654_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(G134gat), .ZN(new_n844_));
  OR3_X1    g643(.A1(new_n816_), .A2(G134gat), .A3(new_n609_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1343gat));
  AOI21_X1  g645(.A(new_n809_), .B1(new_n804_), .B2(new_n643_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n568_), .A2(new_n536_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n847_), .A2(new_n814_), .A3(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n289_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n642_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g653(.A1(new_n850_), .A2(new_n304_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT61), .B(G155gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1346gat));
  NOR4_X1   g656(.A1(new_n847_), .A2(new_n609_), .A3(new_n814_), .A4(new_n849_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT124), .ZN(new_n859_));
  OR3_X1    g658(.A1(new_n858_), .A2(new_n859_), .A3(G162gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n858_), .B2(G162gat), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n654_), .A2(G162gat), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n860_), .A2(new_n861_), .B1(new_n850_), .B2(new_n862_), .ZN(G1347gat));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n543_), .A2(new_n361_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n568_), .A2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n537_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n864_), .B1(new_n821_), .B2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n304_), .B1(new_n801_), .B2(new_n785_), .ZN(new_n870_));
  OAI211_X1 g669(.A(KEYINPUT125), .B(new_n867_), .C1(new_n870_), .C2(new_n809_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n376_), .A3(new_n289_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n289_), .B(new_n867_), .C1(new_n870_), .C2(new_n809_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n874_), .A2(new_n875_), .A3(G169gat), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n874_), .B2(G169gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n873_), .B1(new_n876_), .B2(new_n877_), .ZN(G1348gat));
  AOI21_X1  g677(.A(G176gat), .B1(new_n872_), .B2(new_n642_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n847_), .A2(new_n537_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n866_), .A2(new_n257_), .A3(new_n375_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(G1349gat));
  NAND4_X1  g681(.A1(new_n880_), .A2(new_n568_), .A3(new_n304_), .A4(new_n865_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n643_), .A2(new_n398_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n883_), .A2(new_n379_), .B1(new_n872_), .B2(new_n884_), .ZN(G1350gat));
  AOI21_X1  g684(.A(new_n380_), .B1(new_n872_), .B2(new_n654_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n603_), .A2(new_n399_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT126), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n887_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n872_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n647_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n891_), .B(new_n892_), .C1(new_n380_), .C2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n889_), .A2(new_n894_), .ZN(G1351gat));
  NOR2_X1   g694(.A1(new_n847_), .A2(new_n849_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n289_), .A3(new_n865_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n642_), .A3(new_n865_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n404_), .A2(KEYINPUT127), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1353gat));
  NAND3_X1  g700(.A1(new_n896_), .A2(new_n304_), .A3(new_n865_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  AND2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n902_), .A2(new_n903_), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n902_), .B2(new_n903_), .ZN(G1354gat));
  NAND2_X1  g705(.A1(new_n896_), .A2(new_n865_), .ZN(new_n907_));
  OAI21_X1  g706(.A(G218gat), .B1(new_n907_), .B2(new_n647_), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n609_), .A2(G218gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n907_), .B2(new_n909_), .ZN(G1355gat));
endmodule


