//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n880_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT88), .ZN(new_n203_));
  INV_X1    g002(.A(G204gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G197gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT87), .ZN(new_n206_));
  INV_X1    g005(.A(G197gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G204gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n203_), .A2(new_n209_), .A3(KEYINPUT21), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT89), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n209_), .A2(KEYINPUT21), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT85), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(new_n205_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n208_), .A2(new_n213_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT21), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n217_), .A2(KEYINPUT86), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(KEYINPUT86), .ZN(new_n219_));
  INV_X1    g018(.A(new_n203_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n212_), .A2(new_n218_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n211_), .A2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT83), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n223_), .B1(new_n226_), .B2(KEYINPUT1), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(KEYINPUT1), .B2(new_n226_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G141gat), .A2(G148gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G141gat), .A2(G148gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n230_), .B(KEYINPUT3), .Z(new_n233_));
  XOR2_X1   g032(.A(new_n229_), .B(KEYINPUT2), .Z(new_n234_));
  OAI221_X1 g033(.A(new_n226_), .B1(G155gat), .B2(G162gat), .C1(new_n233_), .C2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT29), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n222_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G228gat), .A2(G233gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n222_), .A2(new_n239_), .A3(new_n237_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G78gat), .B(G106gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n241_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n236_), .A2(KEYINPUT29), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n246_), .A2(new_n247_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G22gat), .B(G50gat), .Z(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OR3_X1    g050(.A1(new_n248_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n251_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n241_), .A2(new_n242_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n243_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n245_), .A2(KEYINPUT90), .ZN(new_n257_));
  AND4_X1   g056(.A1(new_n245_), .A2(new_n254_), .A3(new_n256_), .A4(new_n257_), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n254_), .A2(new_n257_), .B1(new_n256_), .B2(new_n245_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(G169gat), .ZN(new_n261_));
  INV_X1    g060(.A(G176gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(KEYINPUT24), .A3(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G190gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT80), .ZN(new_n267_));
  INV_X1    g066(.A(G183gat), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n268_), .A2(KEYINPUT25), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n266_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT25), .B(G183gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(KEYINPUT80), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT23), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(KEYINPUT24), .B2(new_n263_), .ZN(new_n275_));
  OAI221_X1 g074(.A(new_n265_), .B1(new_n270_), .B2(new_n272_), .C1(new_n275_), .C2(KEYINPUT81), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n275_), .A2(KEYINPUT81), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n274_), .B1(G183gat), .B2(G190gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n280_));
  OR3_X1    g079(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G71gat), .B(G99gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(G43gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n283_), .B(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G127gat), .B(G134gat), .Z(new_n287_));
  XOR2_X1   g086(.A(G113gat), .B(G120gat), .Z(new_n288_));
  XOR2_X1   g087(.A(new_n287_), .B(new_n288_), .Z(new_n289_));
  XNOR2_X1  g088(.A(new_n286_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G227gat), .A2(G233gat), .ZN(new_n291_));
  INV_X1    g090(.A(G15gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT30), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT31), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n290_), .B(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n236_), .A2(new_n289_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n289_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n232_), .A2(new_n298_), .A3(new_n235_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(KEYINPUT4), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n236_), .A2(new_n301_), .A3(new_n289_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT99), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n236_), .A2(KEYINPUT99), .A3(new_n301_), .A4(new_n289_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n300_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n297_), .A2(new_n299_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n310_), .A2(new_n308_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G1gat), .B(G29gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(G57gat), .B(G85gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n315_), .B(new_n316_), .Z(new_n317_));
  NOR2_X1   g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n296_), .A2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(G64gat), .B(G92gat), .Z(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT97), .ZN(new_n325_));
  XOR2_X1   g124(.A(G8gat), .B(G36gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT95), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n211_), .A2(new_n278_), .A3(new_n221_), .A4(new_n282_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT20), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n271_), .B(KEYINPUT92), .ZN(new_n338_));
  INV_X1    g137(.A(new_n266_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n265_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT93), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n275_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n342_), .B1(new_n341_), .B2(new_n340_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G169gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT94), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n264_), .B(new_n279_), .C1(new_n345_), .C2(G176gat), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n343_), .A2(new_n346_), .B1(new_n211_), .B2(new_n221_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n331_), .B(new_n335_), .C1(new_n337_), .C2(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n343_), .A2(new_n346_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n222_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT20), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(new_n222_), .B2(new_n283_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n334_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n348_), .A2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(KEYINPUT20), .B(new_n336_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n331_), .B1(new_n356_), .B2(new_n335_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n330_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT98), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n337_), .A2(new_n347_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT95), .B1(new_n360_), .B2(new_n334_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n361_), .A2(new_n329_), .A3(new_n354_), .A4(new_n348_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT27), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n354_), .A3(new_n348_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(KEYINPUT98), .A3(new_n330_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n356_), .A2(new_n335_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n334_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n330_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n362_), .A2(new_n370_), .A3(KEYINPUT27), .ZN(new_n371_));
  AND4_X1   g170(.A1(new_n260_), .A2(new_n323_), .A3(new_n367_), .A4(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n312_), .A2(new_n317_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n373_), .A2(KEYINPUT33), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n306_), .A2(new_n308_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n310_), .A2(new_n308_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n319_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n373_), .B(KEYINPUT33), .C1(new_n375_), .C2(new_n377_), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n363_), .A2(new_n366_), .B1(new_n374_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n329_), .A2(KEYINPUT32), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n368_), .A2(new_n369_), .A3(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n381_), .B1(new_n365_), .B2(KEYINPUT101), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT101), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n380_), .B1(new_n365_), .B2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n321_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n260_), .B1(new_n379_), .B2(new_n385_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n322_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n296_), .B(KEYINPUT82), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n372_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G15gat), .B(G22gat), .ZN(new_n394_));
  INV_X1    g193(.A(G1gat), .ZN(new_n395_));
  INV_X1    g194(.A(G8gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT14), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G1gat), .B(G8gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G29gat), .B(G36gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G43gat), .B(G50gat), .Z(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G43gat), .B(G50gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n393_), .B1(new_n400_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n404_), .A2(new_n406_), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n398_), .A2(new_n399_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n398_), .A2(new_n399_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(KEYINPUT79), .A4(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(G229gat), .A2(G233gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n400_), .A2(new_n407_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G113gat), .B(G141gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G169gat), .B(G197gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n417_), .B(new_n418_), .Z(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n409_), .B(KEYINPUT15), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n400_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n422_), .A2(new_n413_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n416_), .B(new_n420_), .C1(new_n423_), .C2(new_n414_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n416_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n414_), .B1(new_n422_), .B2(new_n413_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n419_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n392_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G57gat), .B(G64gat), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n430_), .A2(KEYINPUT11), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(KEYINPUT11), .ZN(new_n432_));
  XOR2_X1   g231(.A(G71gat), .B(G78gat), .Z(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n432_), .A2(new_n433_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  OAI22_X1  g236(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(G99gat), .A2(G106gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(G99gat), .B2(G106gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G99gat), .A2(G106gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n444_), .A2(KEYINPUT6), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n438_), .B(new_n441_), .C1(new_n443_), .C2(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(G85gat), .A2(G92gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G85gat), .A2(G92gat), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n446_), .A2(KEYINPUT66), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT66), .B1(new_n446_), .B2(new_n449_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT8), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n443_), .A2(new_n445_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n441_), .A2(new_n438_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n449_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT66), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(new_n452_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n444_), .A2(KEYINPUT6), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n442_), .A2(G99gat), .A3(G106gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G92gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(KEYINPUT9), .ZN(new_n463_));
  AND2_X1   g262(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n447_), .A2(KEYINPUT9), .A3(new_n448_), .ZN(new_n467_));
  OR2_X1    g266(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n468_));
  INV_X1    g267(.A(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  AND4_X1   g270(.A1(new_n461_), .A2(new_n466_), .A3(new_n467_), .A4(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n458_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n437_), .B1(new_n453_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT12), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n476_), .A2(KEYINPUT68), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G230gat), .A2(G233gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n456_), .A2(new_n457_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n446_), .A2(KEYINPUT66), .A3(new_n449_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(KEYINPUT8), .A3(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n472_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n436_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n483_), .A2(new_n484_), .A3(new_n436_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n479_), .A2(new_n480_), .A3(new_n488_), .A4(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT67), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n475_), .A2(new_n491_), .A3(new_n489_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n480_), .B1(new_n485_), .B2(KEYINPUT67), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G120gat), .B(G148gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT5), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G176gat), .B(G204gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n490_), .A2(new_n494_), .A3(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT70), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT70), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n490_), .A2(new_n494_), .A3(new_n501_), .A4(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n498_), .B(KEYINPUT69), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT71), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT71), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n503_), .A2(new_n510_), .A3(new_n507_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(KEYINPUT13), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT13), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n510_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n514_));
  AOI211_X1 g313(.A(KEYINPUT71), .B(new_n506_), .C1(new_n500_), .C2(new_n502_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n513_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n512_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT76), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n421_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n453_), .A2(new_n474_), .A3(new_n409_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n524_), .A2(new_n525_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n521_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n521_), .A2(new_n526_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT73), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n521_), .A2(KEYINPUT73), .A3(new_n526_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n528_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G134gat), .B(G162gat), .Z(new_n534_));
  XNOR2_X1  g333(.A(G190gat), .B(G218gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(KEYINPUT77), .B(KEYINPUT36), .Z(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n518_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT37), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT74), .B(KEYINPUT36), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n542_), .B(KEYINPUT75), .Z(new_n543_));
  AND2_X1   g342(.A1(new_n533_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n533_), .A2(new_n538_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n540_), .A2(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(KEYINPUT37), .B(new_n539_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n436_), .B(new_n400_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554_));
  XOR2_X1   g353(.A(G127gat), .B(G155gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT16), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G183gat), .B(G211gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  OR3_X1    g357(.A1(new_n553_), .A2(new_n554_), .A3(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(KEYINPUT17), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n553_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n549_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT78), .Z(new_n565_));
  AND3_X1   g364(.A1(new_n429_), .A2(new_n517_), .A3(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n566_), .A2(new_n395_), .A3(new_n322_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT38), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n392_), .A2(new_n546_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n517_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n571_), .A2(new_n428_), .A3(new_n562_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(G1gat), .B1(new_n573_), .B2(new_n321_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n567_), .A2(new_n568_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n569_), .A2(new_n574_), .A3(new_n575_), .ZN(G1324gat));
  NAND2_X1  g375(.A1(new_n367_), .A2(new_n371_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n566_), .A2(new_n396_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT102), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(KEYINPUT39), .ZN(new_n580_));
  INV_X1    g379(.A(new_n573_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n577_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n396_), .B1(new_n579_), .B2(KEYINPUT39), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n580_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n577_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n580_), .B(new_n583_), .C1(new_n573_), .C2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n578_), .B1(new_n584_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT40), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n578_), .B(KEYINPUT40), .C1(new_n584_), .C2(new_n587_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(G1325gat));
  AOI21_X1  g391(.A(new_n292_), .B1(new_n581_), .B2(new_n390_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT41), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n566_), .A2(new_n292_), .A3(new_n390_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT103), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n593_), .A2(new_n594_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n597_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n595_), .A2(new_n598_), .A3(new_n599_), .A4(new_n600_), .ZN(G1326gat));
  OAI21_X1  g400(.A(G22gat), .B1(new_n573_), .B2(new_n260_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT42), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n260_), .A2(G22gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT104), .Z(new_n605_));
  NAND2_X1  g404(.A1(new_n566_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(G1327gat));
  NAND2_X1  g406(.A1(new_n546_), .A2(new_n562_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n571_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n429_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(G29gat), .B1(new_n611_), .B2(new_n322_), .ZN(new_n612_));
  OAI21_X1  g411(.A(KEYINPUT43), .B1(new_n392_), .B2(new_n549_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT43), .ZN(new_n614_));
  INV_X1    g413(.A(new_n549_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n390_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n614_), .B(new_n615_), .C1(new_n616_), .C2(new_n372_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n613_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n428_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n517_), .A2(new_n619_), .A3(new_n562_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT44), .B1(new_n618_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT44), .ZN(new_n623_));
  AOI211_X1 g422(.A(new_n623_), .B(new_n620_), .C1(new_n613_), .C2(new_n617_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n322_), .A2(G29gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n612_), .B1(new_n625_), .B2(new_n626_), .ZN(G1328gat));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(KEYINPUT46), .ZN(new_n629_));
  INV_X1    g428(.A(G36gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n625_), .B2(new_n577_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n585_), .A2(G36gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OR3_X1    g432(.A1(new_n610_), .A2(KEYINPUT45), .A3(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT45), .B1(new_n610_), .B2(new_n633_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n629_), .B1(new_n631_), .B2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n622_), .A2(new_n624_), .A3(new_n585_), .ZN(new_n639_));
  OAI221_X1 g438(.A(new_n636_), .B1(new_n628_), .B2(KEYINPUT46), .C1(new_n639_), .C2(new_n630_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(G1329gat));
  INV_X1    g440(.A(new_n296_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(G43gat), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n622_), .A2(new_n624_), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(G43gat), .B1(new_n611_), .B2(new_n390_), .ZN(new_n645_));
  OR3_X1    g444(.A1(new_n644_), .A2(KEYINPUT47), .A3(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT47), .B1(new_n644_), .B2(new_n645_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1330gat));
  INV_X1    g447(.A(new_n260_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(G50gat), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n622_), .A2(new_n624_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652_));
  AOI21_X1  g451(.A(G50gat), .B1(new_n611_), .B2(new_n649_), .ZN(new_n653_));
  OR3_X1    g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n652_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1331gat));
  NAND2_X1  g455(.A1(new_n565_), .A2(new_n571_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n657_), .A2(KEYINPUT107), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(KEYINPUT107), .ZN(new_n659_));
  NOR4_X1   g458(.A1(new_n658_), .A2(new_n659_), .A3(new_n392_), .A4(new_n619_), .ZN(new_n660_));
  INV_X1    g459(.A(G57gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n322_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n570_), .A2(new_n428_), .A3(new_n571_), .A4(new_n563_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G57gat), .B1(new_n663_), .B2(new_n321_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1332gat));
  OAI21_X1  g464(.A(G64gat), .B1(new_n663_), .B2(new_n585_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT48), .ZN(new_n667_));
  INV_X1    g466(.A(G64gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n660_), .A2(new_n668_), .A3(new_n577_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1333gat));
  OAI21_X1  g469(.A(G71gat), .B1(new_n663_), .B2(new_n391_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(G71gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n660_), .A2(new_n674_), .A3(new_n390_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1334gat));
  OAI21_X1  g475(.A(G78gat), .B1(new_n663_), .B2(new_n260_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT50), .ZN(new_n678_));
  INV_X1    g477(.A(G78gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n660_), .A2(new_n679_), .A3(new_n649_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1335gat));
  INV_X1    g480(.A(new_n392_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n517_), .A2(new_n608_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n428_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G85gat), .B1(new_n685_), .B2(new_n322_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n563_), .A2(new_n619_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n618_), .A2(new_n571_), .A3(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n322_), .B1(new_n465_), .B2(new_n464_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT109), .Z(new_n690_));
  AOI21_X1  g489(.A(new_n686_), .B1(new_n688_), .B2(new_n690_), .ZN(G1336gat));
  AOI21_X1  g490(.A(new_n462_), .B1(new_n688_), .B2(new_n577_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n684_), .A2(G92gat), .A3(new_n585_), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n692_), .A2(KEYINPUT110), .A3(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT110), .B1(new_n692_), .B2(new_n693_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1337gat));
  INV_X1    g495(.A(G99gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n688_), .B2(new_n390_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT51), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(KEYINPUT111), .ZN(new_n700_));
  AND4_X1   g499(.A1(new_n642_), .A2(new_n685_), .A3(new_n468_), .A4(new_n470_), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n698_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n700_), .B1(new_n698_), .B2(new_n701_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1338gat));
  NAND4_X1  g503(.A1(new_n618_), .A2(new_n649_), .A3(new_n571_), .A4(new_n687_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n469_), .B1(KEYINPUT113), .B2(KEYINPUT52), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n649_), .A2(new_n469_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n684_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n705_), .B(new_n706_), .C1(KEYINPUT113), .C2(KEYINPUT52), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n709_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT53), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT53), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n709_), .A2(new_n713_), .A3(new_n717_), .A4(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1339gat));
  NOR2_X1   g518(.A1(new_n577_), .A2(new_n649_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n296_), .A2(new_n321_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT117), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n423_), .A2(new_n414_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n413_), .A2(new_n415_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n724_), .B(new_n420_), .C1(new_n414_), .C2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n427_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n503_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT115), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT56), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n489_), .B1(new_n485_), .B2(new_n477_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n480_), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n436_), .B(new_n486_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(KEYINPUT55), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT55), .ZN(new_n738_));
  NOR4_X1   g537(.A1(new_n732_), .A2(new_n734_), .A3(new_n738_), .A4(new_n733_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n731_), .B(new_n504_), .C1(new_n737_), .C2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n503_), .A2(new_n728_), .A3(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n504_), .B1(new_n737_), .B2(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT56), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n730_), .A2(new_n740_), .A3(new_n742_), .A4(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT58), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(KEYINPUT116), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(KEYINPUT116), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n549_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT57), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n728_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n736_), .A2(KEYINPUT55), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n490_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n739_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n505_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n731_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n743_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n428_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n757_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n751_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n546_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n750_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  AOI211_X1 g564(.A(KEYINPUT57), .B(new_n546_), .C1(new_n751_), .C2(new_n762_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n723_), .B1(new_n749_), .B2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n727_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n761_), .B1(new_n755_), .B2(new_n758_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n740_), .A2(KEYINPUT114), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n764_), .B1(new_n769_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT57), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n763_), .A2(new_n750_), .A3(new_n764_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n745_), .A2(KEYINPUT116), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT58), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n745_), .A2(KEYINPUT116), .A3(new_n746_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n615_), .A3(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n776_), .A2(new_n780_), .A3(KEYINPUT117), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n768_), .A2(new_n562_), .A3(new_n781_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n517_), .A2(new_n428_), .A3(new_n563_), .A4(new_n549_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n722_), .B1(new_n782_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(G113gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n619_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n563_), .B1(new_n776_), .B2(new_n780_), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n785_), .A2(new_n790_), .ZN(new_n791_));
  XOR2_X1   g590(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n792_));
  NOR2_X1   g591(.A1(new_n722_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT59), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n787_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n619_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n789_), .B1(new_n799_), .B2(new_n788_), .ZN(G1340gat));
  INV_X1    g599(.A(G120gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n517_), .B2(KEYINPUT60), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n787_), .B(new_n802_), .C1(KEYINPUT60), .C2(new_n801_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n797_), .A2(new_n571_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n805_), .B2(new_n801_), .ZN(G1341gat));
  OAI21_X1  g605(.A(G127gat), .B1(new_n796_), .B2(new_n562_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n787_), .ZN(new_n808_));
  OR3_X1    g607(.A1(new_n808_), .A2(G127gat), .A3(new_n562_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n807_), .A2(new_n809_), .A3(KEYINPUT119), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(G1342gat));
  INV_X1    g613(.A(G134gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n808_), .B2(new_n764_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n816_), .A2(KEYINPUT120), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(KEYINPUT120), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n549_), .A2(new_n815_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n817_), .A2(new_n818_), .B1(new_n797_), .B2(new_n819_), .ZN(G1343gat));
  NAND2_X1  g619(.A1(new_n776_), .A2(new_n780_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n563_), .B1(new_n821_), .B2(new_n723_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n785_), .B1(new_n822_), .B2(new_n781_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n391_), .A2(new_n585_), .A3(new_n322_), .A4(new_n649_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT121), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n782_), .A2(new_n786_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n827_));
  INV_X1    g626(.A(new_n824_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n825_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n619_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT122), .B(G141gat), .Z(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(G1344gat));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n571_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g634(.A(KEYINPUT61), .B(G155gat), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT123), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n830_), .B2(new_n563_), .ZN(new_n839_));
  AOI211_X1 g638(.A(KEYINPUT123), .B(new_n562_), .C1(new_n825_), .C2(new_n829_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n837_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n827_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n842_));
  AOI211_X1 g641(.A(KEYINPUT121), .B(new_n824_), .C1(new_n782_), .C2(new_n786_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n563_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT123), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n830_), .A2(new_n838_), .A3(new_n563_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n836_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n841_), .A2(new_n847_), .ZN(G1346gat));
  INV_X1    g647(.A(new_n830_), .ZN(new_n849_));
  OR3_X1    g648(.A1(new_n849_), .A2(G162gat), .A3(new_n764_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G162gat), .B1(new_n849_), .B2(new_n549_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1347gat));
  NOR2_X1   g651(.A1(new_n785_), .A2(new_n790_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n391_), .A2(new_n585_), .A3(new_n322_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n260_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n857_), .A2(new_n345_), .A3(new_n428_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n261_), .B1(new_n856_), .B2(new_n619_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(KEYINPUT124), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n858_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n859_), .A2(KEYINPUT124), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT62), .B1(new_n859_), .B2(KEYINPUT124), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(G1348gat));
  INV_X1    g664(.A(new_n854_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n826_), .A2(new_n260_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(KEYINPUT125), .ZN(new_n868_));
  OR3_X1    g667(.A1(new_n823_), .A2(KEYINPUT125), .A3(new_n649_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n517_), .A2(new_n262_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n868_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT126), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT126), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n868_), .A2(new_n869_), .A3(new_n873_), .A4(new_n870_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n262_), .B1(new_n857_), .B2(new_n517_), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n872_), .A2(new_n874_), .A3(new_n875_), .ZN(G1349gat));
  AND3_X1   g675(.A1(new_n856_), .A2(new_n338_), .A3(new_n563_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n868_), .A2(new_n563_), .A3(new_n869_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n268_), .ZN(G1350gat));
  NAND2_X1  g678(.A1(new_n856_), .A2(new_n615_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n764_), .A2(new_n339_), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n880_), .A2(G190gat), .B1(new_n856_), .B2(new_n881_), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(KEYINPUT127), .Z(G1351gat));
  AND4_X1   g682(.A1(new_n387_), .A2(new_n826_), .A3(new_n577_), .A4(new_n391_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n619_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n571_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g687(.A1(new_n884_), .A2(new_n563_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT63), .B(G211gat), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n889_), .B2(new_n892_), .ZN(G1354gat));
  INV_X1    g692(.A(G218gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n884_), .A2(new_n894_), .A3(new_n546_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n884_), .A2(new_n615_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n894_), .ZN(G1355gat));
endmodule


