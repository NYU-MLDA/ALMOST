//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n964_, new_n965_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n202_));
  NAND3_X1  g001(.A1(new_n202_), .A2(G183gat), .A3(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT76), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT76), .ZN(new_n205_));
  NAND4_X1  g004(.A1(new_n205_), .A2(new_n202_), .A3(G183gat), .A4(G190gat), .ZN(new_n206_));
  INV_X1    g005(.A(G183gat), .ZN(new_n207_));
  INV_X1    g006(.A(G190gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT23), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n204_), .A2(new_n206_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT26), .B(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n210_), .A2(new_n215_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n209_), .A2(KEYINPUT78), .A3(new_n203_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n207_), .A2(new_n208_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT78), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n223_), .A2(new_n202_), .A3(G183gat), .A4(G190gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n221_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n211_), .A2(KEYINPUT22), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G169gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n229_), .A3(new_n212_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT77), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G169gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT77), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n212_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n234_), .A3(new_n214_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n220_), .B1(new_n226_), .B2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G71gat), .B(G99gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(G43gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n236_), .B(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G113gat), .B(G120gat), .Z(new_n244_));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT80), .B1(new_n242_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT79), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n242_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n249_), .B1(new_n242_), .B2(new_n247_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n246_), .B(new_n248_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G227gat), .A2(G233gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(G15gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT30), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n252_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n241_), .B(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G141gat), .ZN(new_n258_));
  INV_X1    g057(.A(G148gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(KEYINPUT3), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(G141gat), .B2(G148gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT83), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G141gat), .A2(G148gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT2), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n264_), .A2(new_n265_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(KEYINPUT83), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n263_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G155gat), .ZN(new_n271_));
  INV_X1    g070(.A(G162gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT82), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT82), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(G155gat), .B2(G162gat), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n273_), .A2(new_n275_), .B1(G155gat), .B2(G162gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n270_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G155gat), .A2(G162gat), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(KEYINPUT1), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(KEYINPUT1), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT82), .B1(new_n271_), .B2(new_n272_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n274_), .A2(G155gat), .A3(G162gat), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n279_), .B(new_n280_), .C1(new_n281_), .C2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G141gat), .B(G148gat), .Z(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n277_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT29), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT89), .ZN(new_n288_));
  INV_X1    g087(.A(G204gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n288_), .B1(G197gat), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT88), .B(G204gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(G197gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(KEYINPUT88), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT88), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(G204gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G197gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n288_), .A3(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n292_), .A2(new_n298_), .A3(KEYINPUT21), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n293_), .A2(new_n295_), .A3(G197gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT21), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n297_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT90), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(new_n289_), .B2(G197gat), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .A4(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n299_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n300_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n306_), .A2(new_n301_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n307_), .A2(KEYINPUT92), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT92), .B1(new_n307_), .B2(new_n310_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n287_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G228gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT86), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT87), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n316_), .B(new_n319_), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n270_), .A2(new_n276_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n320_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n305_), .A2(new_n306_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n324_), .A2(new_n299_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT91), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n292_), .A2(new_n298_), .A3(KEYINPUT21), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n305_), .A2(new_n306_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n310_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT91), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n287_), .A2(new_n329_), .A3(new_n330_), .A4(new_n320_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n326_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G78gat), .B(G106gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n318_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n335_), .A2(KEYINPUT95), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n321_), .A2(new_n322_), .ZN(new_n337_));
  XOR2_X1   g136(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT85), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n337_), .B(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G22gat), .B(G50gat), .Z(new_n341_));
  XOR2_X1   g140(.A(new_n340_), .B(new_n341_), .Z(new_n342_));
  NAND2_X1  g141(.A1(new_n335_), .A2(KEYINPUT95), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT92), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n329_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n311_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n316_), .B1(new_n346_), .B2(new_n287_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n326_), .A2(new_n331_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n333_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n336_), .A2(new_n342_), .A3(new_n343_), .A4(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n334_), .B1(new_n318_), .B2(new_n332_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n335_), .B1(new_n351_), .B2(KEYINPUT93), .ZN(new_n352_));
  NOR4_X1   g151(.A1(new_n347_), .A2(new_n348_), .A3(KEYINPUT93), .A4(new_n333_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n342_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT94), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n350_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  AOI211_X1 g156(.A(KEYINPUT94), .B(new_n342_), .C1(new_n352_), .C2(new_n354_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT98), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n231_), .A2(new_n234_), .A3(new_n214_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n218_), .A2(new_n215_), .A3(new_n219_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n361_), .A2(new_n225_), .B1(new_n362_), .B2(new_n210_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n360_), .B1(new_n325_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT19), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT96), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n230_), .A2(new_n367_), .A3(new_n214_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n230_), .B2(new_n214_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n210_), .A2(new_n222_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n221_), .A2(new_n224_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n370_), .A2(new_n371_), .B1(new_n362_), .B2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n366_), .B1(new_n325_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n329_), .A2(new_n236_), .A3(KEYINPUT98), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n364_), .A2(new_n374_), .A3(KEYINPUT20), .A4(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT20), .B1(new_n329_), .B2(new_n236_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT97), .B1(new_n325_), .B2(new_n373_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n362_), .A2(new_n372_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n369_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n230_), .A2(new_n367_), .A3(new_n214_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n371_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT97), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n329_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n377_), .B1(new_n378_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n366_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n376_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G8gat), .B(G36gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT18), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G64gat), .B(G92gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G1gat), .B(G29gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G57gat), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n250_), .A2(new_n251_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n246_), .A2(new_n248_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n286_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n243_), .A2(new_n244_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n242_), .A2(new_n247_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n277_), .A2(new_n405_), .A3(new_n285_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n407_), .A2(KEYINPUT103), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT100), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n407_), .B2(KEYINPUT103), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n399_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n406_), .B(KEYINPUT4), .C1(new_n321_), .C2(new_n252_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT99), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n402_), .A2(KEYINPUT99), .A3(KEYINPUT4), .A4(new_n406_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n411_), .B1(new_n402_), .B2(KEYINPUT4), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n413_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n376_), .B(new_n392_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n394_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT101), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n410_), .B1(new_n402_), .B2(KEYINPUT4), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n423_), .B1(new_n418_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n402_), .A2(new_n406_), .A3(new_n411_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n424_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n428_), .B2(KEYINPUT101), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n425_), .A2(new_n429_), .A3(new_n399_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT33), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n425_), .A2(new_n429_), .A3(new_n432_), .A4(new_n399_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n422_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT104), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n364_), .A2(KEYINPUT20), .A3(new_n375_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n312_), .A2(new_n313_), .A3(new_n383_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n366_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n386_), .A2(new_n387_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n392_), .A2(KEYINPUT32), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n376_), .B(new_n443_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT105), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n442_), .A2(new_n444_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n445_), .A2(new_n446_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n430_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n399_), .B1(new_n425_), .B2(new_n429_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n447_), .B(new_n448_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n359_), .B1(new_n437_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n442_), .A2(new_n393_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT106), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(KEYINPUT27), .A4(new_n421_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n421_), .A2(KEYINPUT27), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n392_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT106), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n394_), .A2(new_n421_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT27), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n456_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n449_), .A2(new_n450_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n463_), .B(new_n465_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n257_), .B1(new_n453_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n359_), .A2(new_n463_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n257_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G29gat), .B(G36gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G43gat), .B(G50gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT15), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G15gat), .B(G22gat), .ZN(new_n476_));
  INV_X1    g275(.A(G1gat), .ZN(new_n477_));
  INV_X1    g276(.A(G8gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT14), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G8gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n475_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n482_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(new_n474_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n474_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n474_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n482_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n483_), .A2(new_n487_), .B1(new_n491_), .B2(new_n485_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G113gat), .B(G141gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(G169gat), .B(G197gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n492_), .B(new_n495_), .Z(new_n496_));
  NOR2_X1   g295(.A1(new_n471_), .A2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(KEYINPUT10), .B(G99gat), .Z(new_n498_));
  INV_X1    g297(.A(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G85gat), .B(G92gat), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT9), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT6), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(G99gat), .A3(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(G85gat), .ZN(new_n508_));
  INV_X1    g307(.A(G92gat), .ZN(new_n509_));
  OR3_X1    g308(.A1(new_n508_), .A2(new_n509_), .A3(KEYINPUT9), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n500_), .A2(new_n502_), .A3(new_n507_), .A4(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT68), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n504_), .A2(new_n506_), .A3(KEYINPUT65), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT65), .B1(new_n504_), .B2(new_n506_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT7), .ZN(new_n515_));
  INV_X1    g314(.A(G99gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n516_), .A3(new_n499_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n513_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n501_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT8), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n519_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT8), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT64), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n524_), .A2(KEYINPUT64), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n501_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n512_), .B1(new_n522_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT65), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n507_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n519_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n504_), .A2(new_n506_), .A3(KEYINPUT65), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n524_), .B1(new_n535_), .B2(new_n501_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n536_), .A2(KEYINPUT68), .A3(new_n528_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n511_), .B1(new_n530_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n475_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT71), .ZN(new_n541_));
  XOR2_X1   g340(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT35), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT72), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(new_n543_), .B2(KEYINPUT35), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n511_), .B1(new_n536_), .B2(new_n528_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n547_), .B1(new_n548_), .B2(new_n489_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n539_), .A2(new_n544_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n544_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n475_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n522_), .A2(new_n512_), .A3(new_n529_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT68), .B1(new_n536_), .B2(new_n528_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n553_), .B1(new_n556_), .B2(new_n511_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n552_), .B1(new_n557_), .B2(new_n549_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(KEYINPUT36), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n551_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n561_), .B(KEYINPUT36), .Z(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n551_), .B2(new_n558_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT37), .B1(new_n563_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT73), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT73), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n569_), .B(KEYINPUT37), .C1(new_n563_), .C2(new_n566_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n544_), .B1(new_n539_), .B2(new_n550_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n557_), .A2(new_n552_), .A3(new_n549_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n564_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT37), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n551_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT74), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n574_), .A2(KEYINPUT74), .A3(new_n575_), .A4(new_n576_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n571_), .A2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G127gat), .B(G155gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590_));
  NOR2_X1   g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G57gat), .B(G64gat), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n592_), .B1(new_n593_), .B2(KEYINPUT11), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT66), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n593_), .B2(KEYINPUT11), .ZN(new_n596_));
  INV_X1    g395(.A(G64gat), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(G57gat), .ZN(new_n598_));
  INV_X1    g397(.A(G57gat), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(G64gat), .ZN(new_n600_));
  AND4_X1   g399(.A1(new_n595_), .A2(new_n598_), .A3(new_n600_), .A4(KEYINPUT11), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n594_), .B1(new_n596_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n598_), .A2(new_n600_), .A3(KEYINPUT11), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT66), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n600_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT11), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n598_), .A2(new_n600_), .A3(new_n595_), .A4(KEYINPUT11), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n604_), .A2(new_n607_), .A3(new_n592_), .A4(new_n608_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n602_), .A2(new_n609_), .A3(KEYINPUT67), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT67), .B1(new_n602_), .B2(new_n609_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n482_), .B(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n589_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n602_), .A2(new_n609_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n620_), .A2(new_n588_), .A3(new_n587_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n619_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n622_), .B2(new_n615_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n618_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n582_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT12), .ZN(new_n627_));
  INV_X1    g426(.A(new_n511_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n522_), .B2(new_n529_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n627_), .B1(new_n612_), .B2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n612_), .B2(new_n629_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n628_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n619_), .A2(new_n627_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n630_), .B(new_n632_), .C1(new_n633_), .C2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n612_), .A2(new_n629_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n548_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n631_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(G120gat), .B(G148gat), .Z(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n636_), .A2(new_n639_), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n645_), .B1(new_n636_), .B2(new_n639_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(KEYINPUT13), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(KEYINPUT13), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n626_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n497_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(new_n477_), .A3(new_n464_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT38), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n653_), .A2(new_n496_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n625_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n257_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n342_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n347_), .A2(new_n333_), .A3(new_n348_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT93), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(new_n349_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n662_), .B1(new_n665_), .B2(new_n353_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT94), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n355_), .A2(new_n356_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n350_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n431_), .A2(new_n433_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n422_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n447_), .A2(new_n448_), .ZN(new_n673_));
  AOI22_X1  g472(.A1(new_n672_), .A2(KEYINPUT104), .B1(new_n464_), .B2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n669_), .B1(new_n674_), .B2(new_n436_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n466_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n661_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n470_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n563_), .A2(new_n566_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT107), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT108), .B1(new_n679_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(KEYINPUT108), .B(new_n681_), .C1(new_n467_), .C2(new_n470_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n660_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(new_n464_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n658_), .B1(new_n477_), .B2(new_n686_), .ZN(G1324gat));
  INV_X1    g486(.A(new_n463_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n656_), .A2(new_n478_), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n660_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n684_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n688_), .B(new_n690_), .C1(new_n682_), .C2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT109), .B(KEYINPUT39), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(G8gat), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n692_), .B2(G8gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n689_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT40), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT40), .B(new_n689_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1325gat));
  OR3_X1    g499(.A1(new_n655_), .A2(G15gat), .A3(new_n661_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n685_), .A2(new_n257_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n702_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT41), .B1(new_n702_), .B2(G15gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n701_), .B1(new_n703_), .B2(new_n704_), .ZN(G1326gat));
  OR3_X1    g504(.A1(new_n655_), .A2(G22gat), .A3(new_n359_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n685_), .A2(new_n669_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(G22gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n707_), .B2(G22gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(G1327gat));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n582_), .B(KEYINPUT110), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n713_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n582_), .A2(KEYINPUT43), .ZN(new_n715_));
  AOI22_X1  g514(.A1(KEYINPUT43), .A2(new_n714_), .B1(new_n679_), .B2(new_n715_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n653_), .A2(new_n496_), .A3(new_n625_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n712_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n679_), .B2(new_n713_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n715_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n471_), .A2(new_n722_), .ZN(new_n723_));
  OAI211_X1 g522(.A(KEYINPUT44), .B(new_n717_), .C1(new_n721_), .C2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n719_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(G29gat), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n465_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n496_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n680_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(new_n625_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n652_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n679_), .A2(new_n728_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n679_), .A2(KEYINPUT111), .A3(new_n728_), .A4(new_n731_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(new_n464_), .A3(new_n735_), .ZN(new_n736_));
  AOI22_X1  g535(.A1(new_n725_), .A2(new_n727_), .B1(new_n726_), .B2(new_n736_), .ZN(G1328gat));
  NAND3_X1  g536(.A1(new_n719_), .A2(new_n688_), .A3(new_n724_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G36gat), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n463_), .A2(G36gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n734_), .A2(new_n735_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT45), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n734_), .A2(new_n743_), .A3(new_n735_), .A4(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n739_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT46), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n739_), .A2(KEYINPUT46), .A3(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1329gat));
  NAND4_X1  g549(.A1(new_n719_), .A2(G43gat), .A3(new_n724_), .A4(new_n257_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n734_), .A2(new_n257_), .A3(new_n735_), .ZN(new_n752_));
  INV_X1    g551(.A(G43gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n751_), .A2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g555(.A(G50gat), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n359_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n734_), .A2(new_n669_), .A3(new_n735_), .ZN(new_n759_));
  AOI22_X1  g558(.A1(new_n725_), .A2(new_n758_), .B1(new_n757_), .B2(new_n759_), .ZN(G1331gat));
  NOR2_X1   g559(.A1(new_n652_), .A2(new_n728_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n679_), .A2(new_n761_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(new_n626_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n599_), .A3(new_n464_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n761_), .A2(new_n625_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(new_n464_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n765_), .B1(new_n768_), .B2(new_n599_), .ZN(G1332gat));
  NAND3_X1  g568(.A1(new_n764_), .A2(new_n597_), .A3(new_n688_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT48), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n767_), .A2(new_n688_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(G64gat), .ZN(new_n773_));
  AOI211_X1 g572(.A(KEYINPUT48), .B(new_n597_), .C1(new_n767_), .C2(new_n688_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(G1333gat));
  INV_X1    g574(.A(G71gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n764_), .A2(new_n776_), .A3(new_n257_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n767_), .A2(new_n257_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(G71gat), .ZN(new_n780_));
  AOI211_X1 g579(.A(KEYINPUT49), .B(new_n776_), .C1(new_n767_), .C2(new_n257_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(G1334gat));
  OR3_X1    g581(.A1(new_n763_), .A2(G78gat), .A3(new_n359_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n767_), .A2(new_n669_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(G78gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G78gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(G1335gat));
  NAND2_X1  g587(.A1(new_n714_), .A2(KEYINPUT43), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n679_), .A2(new_n715_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n789_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n761_), .A2(new_n624_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n791_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(G85gat), .B1(new_n797_), .B2(new_n465_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n679_), .A2(new_n730_), .A3(new_n761_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(new_n508_), .A3(new_n464_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(new_n801_), .ZN(G1336gat));
  OAI21_X1  g601(.A(G92gat), .B1(new_n797_), .B2(new_n463_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(new_n509_), .A3(new_n688_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1337gat));
  NAND3_X1  g604(.A1(new_n800_), .A2(new_n257_), .A3(new_n498_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n795_), .A2(new_n661_), .A3(new_n796_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n516_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT51), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n810_), .B(new_n806_), .C1(new_n807_), .C2(new_n516_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1338gat));
  NAND3_X1  g611(.A1(new_n800_), .A2(new_n499_), .A3(new_n669_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n789_), .A2(new_n790_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n793_), .A2(new_n359_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n814_), .B1(new_n817_), .B2(G106gat), .ZN(new_n818_));
  AOI211_X1 g617(.A(KEYINPUT52), .B(new_n499_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n813_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT53), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(new_n813_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1339gat));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825_));
  INV_X1    g624(.A(G113gat), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n496_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n468_), .A2(new_n465_), .A3(new_n661_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n729_), .A2(KEYINPUT57), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n495_), .B1(new_n491_), .B2(new_n484_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n483_), .A2(new_n488_), .A3(new_n485_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n492_), .A2(new_n495_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n728_), .A2(new_n646_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n612_), .A2(new_n629_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n630_), .B(new_n839_), .C1(new_n633_), .C2(new_n635_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n631_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n636_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n538_), .A2(new_n634_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n844_), .A2(KEYINPUT55), .A3(new_n630_), .A4(new_n632_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(new_n843_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n644_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT113), .B(KEYINPUT56), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n846_), .A2(KEYINPUT56), .A3(new_n644_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n838_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n837_), .B1(new_n852_), .B2(KEYINPUT114), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n496_), .A2(new_n647_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n846_), .A2(KEYINPUT56), .A3(new_n644_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n848_), .B1(new_n846_), .B2(new_n644_), .ZN(new_n856_));
  OAI211_X1 g655(.A(KEYINPUT114), .B(new_n854_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n833_), .B1(new_n853_), .B2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n646_), .A2(new_n836_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n646_), .A2(KEYINPUT116), .A3(new_n836_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT56), .B1(new_n846_), .B2(new_n644_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n855_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n568_), .A2(new_n570_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n864_), .B(KEYINPUT58), .C1(new_n855_), .C2(new_n865_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n868_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n859_), .A2(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n837_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n854_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT114), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n857_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n874_), .B1(new_n879_), .B2(new_n729_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n624_), .B1(new_n872_), .B2(new_n880_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n582_), .A2(new_n652_), .A3(new_n496_), .A4(new_n625_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT54), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n831_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n829_), .B1(new_n884_), .B2(KEYINPUT117), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n832_), .B1(new_n878_), .B2(new_n857_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n868_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n729_), .B1(new_n853_), .B2(new_n858_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n873_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n625_), .B1(new_n889_), .B2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n882_), .B(new_n893_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n886_), .B(new_n830_), .C1(new_n892_), .C2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n885_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n895_), .A2(new_n896_), .A3(new_n829_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n828_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G113gat), .B1(new_n884_), .B2(new_n728_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n825_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(KEYINPUT117), .B1(new_n884_), .B2(new_n886_), .ZN(new_n903_));
  OAI211_X1 g702(.A(KEYINPUT117), .B(new_n830_), .C1(new_n892_), .C2(new_n894_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT59), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n899_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n827_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n901_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n907_), .A2(KEYINPUT119), .A3(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n902_), .A2(new_n909_), .ZN(G1340gat));
  INV_X1    g709(.A(G120gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n911_), .B1(new_n652_), .B2(KEYINPUT60), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n884_), .B(new_n912_), .C1(KEYINPUT60), .C2(new_n911_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n652_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n911_), .ZN(G1341gat));
  INV_X1    g714(.A(G127gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n884_), .A2(new_n916_), .A3(new_n625_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n624_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n916_), .ZN(G1342gat));
  INV_X1    g718(.A(new_n681_), .ZN(new_n920_));
  AOI21_X1  g719(.A(G134gat), .B1(new_n884_), .B2(new_n920_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(KEYINPUT120), .Z(new_n922_));
  INV_X1    g721(.A(G134gat), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n582_), .A2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n906_), .B2(new_n924_), .ZN(G1343gat));
  AOI21_X1  g724(.A(new_n257_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n359_), .A2(new_n688_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n926_), .A2(new_n464_), .A3(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n496_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(new_n258_), .ZN(G1344gat));
  NOR2_X1   g729(.A1(new_n928_), .A2(new_n652_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(new_n259_), .ZN(G1345gat));
  INV_X1    g731(.A(new_n928_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n933_), .A2(new_n934_), .A3(new_n625_), .ZN(new_n935_));
  OAI21_X1  g734(.A(KEYINPUT121), .B1(new_n928_), .B2(new_n624_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT61), .B(G155gat), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n937_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1346gat));
  NAND3_X1  g739(.A1(new_n933_), .A2(G162gat), .A3(new_n713_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n272_), .B1(new_n928_), .B2(new_n681_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n941_), .A2(KEYINPUT122), .A3(new_n942_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(G1347gat));
  NOR3_X1   g746(.A1(new_n469_), .A2(new_n669_), .A3(new_n463_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n948_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n949_));
  OAI21_X1  g748(.A(G169gat), .B1(new_n949_), .B2(new_n496_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n950_), .A2(KEYINPUT62), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(KEYINPUT62), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n728_), .A2(new_n232_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(KEYINPUT123), .ZN(new_n954_));
  OAI22_X1  g753(.A1(new_n951_), .A2(new_n952_), .B1(new_n949_), .B2(new_n954_), .ZN(G1348gat));
  NOR2_X1   g754(.A1(new_n949_), .A2(new_n652_), .ZN(new_n956_));
  XOR2_X1   g755(.A(KEYINPUT124), .B(G176gat), .Z(new_n957_));
  XNOR2_X1  g756(.A(new_n956_), .B(new_n957_), .ZN(G1349gat));
  NOR2_X1   g757(.A1(new_n949_), .A2(new_n624_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n207_), .A2(KEYINPUT125), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n959_), .A2(new_n216_), .A3(new_n960_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(KEYINPUT125), .A2(G183gat), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n961_), .B1(new_n959_), .B2(new_n962_), .ZN(G1350gat));
  OAI21_X1  g762(.A(G190gat), .B1(new_n949_), .B2(new_n582_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n920_), .A2(new_n217_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n964_), .B1(new_n949_), .B2(new_n965_), .ZN(G1351gat));
  NOR3_X1   g765(.A1(new_n359_), .A2(new_n464_), .A3(new_n463_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n926_), .A2(new_n967_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n968_), .A2(new_n496_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(KEYINPUT126), .B(G197gat), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n969_), .B(new_n970_), .ZN(G1352gat));
  NOR2_X1   g770(.A1(new_n968_), .A2(new_n652_), .ZN(new_n972_));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n972_), .B1(new_n973_), .B2(G204gat), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n291_), .B1(KEYINPUT127), .B2(G204gat), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n974_), .B1(new_n972_), .B2(new_n975_), .ZN(G1353gat));
  NOR2_X1   g775(.A1(new_n968_), .A2(new_n624_), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n977_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n978_));
  XOR2_X1   g777(.A(KEYINPUT63), .B(G211gat), .Z(new_n979_));
  AOI21_X1  g778(.A(new_n978_), .B1(new_n977_), .B2(new_n979_), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n968_), .B2(new_n582_), .ZN(new_n981_));
  OR2_X1    g780(.A1(new_n681_), .A2(G218gat), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n981_), .B1(new_n968_), .B2(new_n982_), .ZN(G1355gat));
endmodule


