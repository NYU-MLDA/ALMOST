//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G29gat), .B(G36gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n208_), .B(new_n211_), .Z(new_n212_));
  NAND2_X1  g011(.A1(G229gat), .A2(G233gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n211_), .B(KEYINPUT15), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(new_n208_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n208_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n214_), .B1(new_n217_), .B2(new_n211_), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n212_), .A2(new_n214_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(G113gat), .B(G141gat), .Z(new_n220_));
  XNOR2_X1  g019(.A(G169gat), .B(G197gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n219_), .B(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT96), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G225gat), .A2(G233gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT4), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G113gat), .B(G120gat), .ZN(new_n229_));
  XOR2_X1   g028(.A(G127gat), .B(G134gat), .Z(new_n230_));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT76), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n229_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n234_), .A3(new_n229_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(G155gat), .A2(G162gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G155gat), .A2(G162gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n242_));
  INV_X1    g041(.A(G141gat), .ZN(new_n243_));
  INV_X1    g042(.A(G148gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT78), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n243_), .B(new_n244_), .C1(new_n245_), .C2(KEYINPUT3), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n247_), .B(KEYINPUT78), .C1(G141gat), .C2(G148gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G141gat), .A2(G148gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT2), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT79), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n250_), .A2(new_n255_), .A3(new_n251_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n255_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n242_), .B1(new_n254_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n250_), .A2(new_n251_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT79), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n250_), .A2(new_n255_), .A3(new_n251_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n252_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT80), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n241_), .B1(new_n259_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT77), .ZN(new_n267_));
  OR3_X1    g066(.A1(new_n240_), .A2(new_n267_), .A3(KEYINPUT1), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n267_), .B1(new_n240_), .B2(KEYINPUT1), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n240_), .A2(KEYINPUT1), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n268_), .A2(new_n239_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n243_), .A2(new_n244_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n250_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n238_), .B1(new_n266_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n241_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT80), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT80), .B1(new_n263_), .B2(new_n264_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n232_), .A2(new_n234_), .A3(new_n229_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n280_), .A2(new_n235_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n281_), .A3(new_n273_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n275_), .A2(KEYINPUT91), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n273_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT91), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n285_), .A3(new_n238_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n228_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n275_), .A2(KEYINPUT4), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n227_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n283_), .A2(new_n226_), .A3(new_n286_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G1gat), .B(G29gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(G85gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT0), .B(G57gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n292_), .B(new_n293_), .Z(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n289_), .A2(new_n290_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n295_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n225_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n289_), .A2(new_n290_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n294_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(KEYINPUT96), .A3(new_n296_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT23), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OR3_X1    g107(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT25), .B(G183gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT26), .B(G190gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(KEYINPUT74), .A2(G169gat), .A3(G176gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n313_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n310_), .B1(new_n321_), .B2(KEYINPUT75), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n313_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT22), .B(G169gat), .ZN(new_n326_));
  INV_X1    g125(.A(G176gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n306_), .B(new_n307_), .C1(G183gat), .C2(G190gat), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n318_), .A2(new_n319_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n325_), .A2(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G71gat), .B(G99gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(G43gat), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n334_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n281_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G227gat), .A2(G233gat), .ZN(new_n339_));
  INV_X1    g138(.A(G15gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT30), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT31), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n335_), .A2(new_n238_), .A3(new_n336_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n338_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n343_), .B1(new_n338_), .B2(new_n344_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G211gat), .B(G218gat), .Z(new_n348_));
  INV_X1    g147(.A(G197gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G204gat), .ZN(new_n350_));
  INV_X1    g149(.A(G204gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G197gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n348_), .A2(KEYINPUT21), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT83), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n350_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT21), .B1(new_n350_), .B2(new_n356_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT84), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT21), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n351_), .A2(G197gat), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(KEYINPUT83), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT84), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n350_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n359_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n350_), .A2(new_n352_), .A3(new_n360_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT85), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT85), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n350_), .A2(new_n352_), .A3(new_n369_), .A4(new_n360_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n348_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n355_), .B1(new_n366_), .B2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n372_), .B1(new_n284_), .B2(KEYINPUT29), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT28), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n279_), .A2(new_n375_), .A3(new_n376_), .A4(new_n273_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT28), .B1(new_n284_), .B2(KEYINPUT29), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n374_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n377_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n373_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(KEYINPUT81), .A2(G233gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(KEYINPUT81), .A2(G233gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(G228gat), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n385_), .B(KEYINPUT82), .Z(new_n386_));
  OAI21_X1  g185(.A(new_n386_), .B1(new_n372_), .B2(KEYINPUT86), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G78gat), .ZN(new_n388_));
  INV_X1    g187(.A(G78gat), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n389_), .B(new_n386_), .C1(new_n372_), .C2(KEYINPUT86), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G106gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n388_), .A2(G106gat), .A3(new_n390_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G22gat), .B(G50gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n393_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n396_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n382_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n393_), .A2(new_n394_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n395_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n382_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n397_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n347_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT18), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n407_), .B(new_n408_), .Z(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT20), .ZN(new_n411_));
  INV_X1    g210(.A(new_n331_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n411_), .B1(new_n413_), .B2(new_n372_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n365_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n363_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n371_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n354_), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n326_), .A2(KEYINPUT88), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n326_), .A2(KEYINPUT88), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n327_), .A3(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n329_), .A2(new_n330_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n308_), .A2(new_n309_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n311_), .A2(new_n312_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT89), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n418_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n421_), .A2(new_n422_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT89), .B1(new_n372_), .B2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n414_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G226gat), .A2(G233gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(KEYINPUT90), .A3(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT20), .B1(new_n418_), .B2(new_n427_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n413_), .A2(new_n372_), .ZN(new_n439_));
  OR3_X1    g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n436_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT90), .B1(new_n432_), .B2(new_n436_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n410_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n432_), .A2(new_n436_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT90), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n446_), .A2(new_n409_), .A3(new_n440_), .A4(new_n437_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT27), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n436_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n450_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n449_), .B1(new_n451_), .B2(new_n410_), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n448_), .A2(new_n449_), .B1(new_n447_), .B2(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n303_), .A2(new_n405_), .A3(new_n453_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n297_), .A2(new_n298_), .A3(new_n225_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT96), .B1(new_n301_), .B2(new_n296_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n453_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n400_), .A2(new_n404_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n347_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n409_), .A2(KEYINPUT32), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n301_), .A2(new_n296_), .B1(new_n461_), .B2(new_n451_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n446_), .A2(new_n440_), .A3(new_n437_), .A4(new_n460_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT95), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n458_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT92), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT33), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n301_), .B2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n298_), .A2(KEYINPUT92), .A3(KEYINPUT33), .ZN(new_n470_));
  INV_X1    g269(.A(new_n448_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n283_), .A2(new_n286_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n294_), .B1(new_n472_), .B2(new_n227_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT94), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  OR3_X1    g274(.A1(new_n287_), .A2(new_n227_), .A3(new_n288_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n474_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .A4(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT93), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n301_), .B2(new_n468_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n298_), .A2(KEYINPUT93), .A3(KEYINPUT33), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n466_), .B1(new_n479_), .B2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n454_), .B1(new_n459_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(KEYINPUT10), .B(G99gat), .Z(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n392_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G85gat), .B(G92gat), .Z(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT9), .ZN(new_n493_));
  INV_X1    g292(.A(G85gat), .ZN(new_n494_));
  INV_X1    g293(.A(G92gat), .ZN(new_n495_));
  OR3_X1    g294(.A1(new_n494_), .A2(new_n495_), .A3(KEYINPUT9), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n489_), .A2(new_n491_), .A3(new_n493_), .A4(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT8), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n488_), .A2(new_n500_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT64), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT65), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n492_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n498_), .B1(new_n504_), .B2(new_n507_), .ZN(new_n508_));
  AOI211_X1 g307(.A(KEYINPUT8), .B(new_n506_), .C1(new_n501_), .C2(new_n503_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n497_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT66), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n513_));
  XOR2_X1   g312(.A(G71gat), .B(G78gat), .Z(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n513_), .A2(new_n514_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT12), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT66), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n522_), .B(new_n497_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n511_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n510_), .A2(new_n519_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT12), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G230gat), .A2(G233gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n517_), .A2(new_n518_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n497_), .B(new_n529_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n524_), .A2(new_n527_), .A3(new_n528_), .A4(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n525_), .A2(new_n530_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(G230gat), .A3(G233gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G120gat), .B(G148gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(G176gat), .B(G204gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n534_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n531_), .A2(new_n533_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT13), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n540_), .A2(KEYINPUT13), .A3(new_n542_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT37), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT34), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT35), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT68), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n551_), .A2(KEYINPUT35), .ZN(new_n555_));
  INV_X1    g354(.A(new_n497_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n504_), .A2(new_n507_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT8), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n504_), .A2(new_n498_), .A3(new_n507_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n556_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  AOI211_X1 g359(.A(new_n554_), .B(new_n555_), .C1(new_n560_), .C2(new_n211_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n552_), .A2(new_n553_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n511_), .A2(new_n215_), .A3(new_n523_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n562_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G190gat), .B(G218gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n569_), .A2(KEYINPUT36), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(KEYINPUT36), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n566_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n570_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n549_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n573_), .A2(new_n549_), .A3(new_n574_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n208_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(new_n519_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT72), .ZN(new_n582_));
  XOR2_X1   g381(.A(G127gat), .B(G155gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT70), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT71), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n584_), .B(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(KEYINPUT69), .B(KEYINPUT16), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT17), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n582_), .B(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n589_), .A2(KEYINPUT17), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n591_), .B1(new_n581_), .B2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT73), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n578_), .A2(new_n594_), .ZN(new_n595_));
  OR4_X1    g394(.A1(new_n224_), .A2(new_n485_), .A3(new_n548_), .A4(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT97), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n303_), .B(KEYINPUT98), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(new_n203_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT38), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n594_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n573_), .A2(new_n574_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n485_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n548_), .A2(new_n224_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G1gat), .B1(new_n607_), .B2(new_n303_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n599_), .A2(new_n600_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n601_), .A2(new_n608_), .A3(new_n609_), .ZN(G1324gat));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n611_));
  OAI221_X1 g410(.A(G8gat), .B1(KEYINPUT99), .B2(new_n611_), .C1(new_n607_), .C2(new_n453_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(KEYINPUT99), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n453_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n597_), .A2(new_n204_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(G1325gat));
  NAND3_X1  g418(.A1(new_n605_), .A2(new_n347_), .A3(new_n606_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(G15gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT41), .Z(new_n622_));
  NAND2_X1  g421(.A1(new_n347_), .A2(new_n340_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n622_), .B1(new_n596_), .B2(new_n623_), .ZN(G1326gat));
  INV_X1    g423(.A(new_n458_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G22gat), .B1(new_n607_), .B2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT42), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n625_), .A2(G22gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n627_), .B1(new_n596_), .B2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT101), .Z(G1327gat));
  NAND2_X1  g429(.A1(new_n602_), .A2(new_n604_), .ZN(new_n631_));
  NOR4_X1   g430(.A1(new_n485_), .A2(new_n631_), .A3(new_n224_), .A4(new_n548_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n303_), .A2(G29gat), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n548_), .A2(new_n594_), .A3(new_n224_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT43), .B1(new_n485_), .B2(new_n578_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n485_), .A2(KEYINPUT43), .A3(new_n578_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n636_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NOR4_X1   g438(.A1(new_n485_), .A2(KEYINPUT102), .A3(KEYINPUT43), .A4(new_n578_), .ZN(new_n640_));
  OAI211_X1 g439(.A(KEYINPUT44), .B(new_n635_), .C1(new_n639_), .C2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n644_));
  INV_X1    g443(.A(new_n577_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n575_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n459_), .A2(new_n484_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n644_), .B(new_n646_), .C1(new_n647_), .C2(new_n454_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT102), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n637_), .A2(new_n638_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n636_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n651_), .A2(KEYINPUT105), .A3(KEYINPUT44), .A4(new_n635_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n643_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n635_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT104), .B1(new_n654_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n658_));
  AOI211_X1 g457(.A(new_n658_), .B(new_n655_), .C1(new_n651_), .C2(new_n635_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n653_), .B(new_n598_), .C1(new_n657_), .C2(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT106), .B1(new_n660_), .B2(G29gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n634_), .B1(new_n661_), .B2(new_n662_), .ZN(G1328gat));
  INV_X1    g462(.A(G36gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n632_), .A2(new_n664_), .A3(new_n615_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT45), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n653_), .B(new_n615_), .C1(new_n657_), .C2(new_n659_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G36gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G36gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI211_X1 g472(.A(KEYINPUT46), .B(new_n666_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1329gat));
  NOR2_X1   g474(.A1(new_n657_), .A2(new_n659_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n643_), .B2(new_n652_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n347_), .A2(G43gat), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n632_), .A2(new_n347_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT108), .B(G43gat), .ZN(new_n680_));
  AOI22_X1  g479(.A1(new_n677_), .A2(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(G1330gat));
  AOI21_X1  g482(.A(G50gat), .B1(new_n632_), .B2(new_n458_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n458_), .A2(G50gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n677_), .B2(new_n685_), .ZN(G1331gat));
  NOR2_X1   g485(.A1(new_n547_), .A2(new_n223_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n605_), .A2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT110), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G57gat), .B1(new_n690_), .B2(new_n303_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n485_), .A2(new_n223_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n692_), .A2(new_n548_), .A3(new_n594_), .A4(new_n578_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n598_), .ZN(new_n694_));
  OR3_X1    g493(.A1(new_n693_), .A2(G57gat), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n691_), .A2(new_n695_), .ZN(G1332gat));
  INV_X1    g495(.A(G64gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n689_), .B2(new_n615_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT48), .Z(new_n699_));
  INV_X1    g498(.A(new_n693_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(new_n697_), .A3(new_n615_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1333gat));
  INV_X1    g501(.A(G71gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n689_), .B2(new_n347_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT49), .Z(new_n705_));
  NAND3_X1  g504(.A1(new_n700_), .A2(new_n703_), .A3(new_n347_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1334gat));
  AOI21_X1  g506(.A(new_n389_), .B1(new_n689_), .B2(new_n458_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT50), .Z(new_n709_));
  NAND3_X1  g508(.A1(new_n700_), .A2(new_n389_), .A3(new_n458_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1335gat));
  NOR2_X1   g510(.A1(new_n631_), .A2(new_n547_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n692_), .A2(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n494_), .B1(new_n713_), .B2(new_n694_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT111), .ZN(new_n715_));
  INV_X1    g514(.A(new_n651_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n716_), .A2(KEYINPUT112), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(KEYINPUT112), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n602_), .A2(new_n687_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n717_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n303_), .A2(new_n494_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n715_), .B1(new_n720_), .B2(new_n721_), .ZN(G1336gat));
  INV_X1    g521(.A(new_n713_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G92gat), .B1(new_n723_), .B2(new_n615_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n453_), .A2(new_n495_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT113), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n720_), .B2(new_n726_), .ZN(G1337gat));
  NAND2_X1  g526(.A1(new_n720_), .A2(new_n347_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(G99gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n723_), .A2(new_n347_), .A3(new_n490_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g531(.A1(new_n602_), .A2(new_n687_), .A3(new_n458_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G106gat), .B1(new_n716_), .B2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT52), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n723_), .A2(new_n392_), .A3(new_n458_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g537(.A(KEYINPUT59), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT57), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n542_), .A2(new_n223_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n530_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n526_), .B2(new_n525_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n528_), .B1(new_n743_), .B2(new_n524_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT55), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n531_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n743_), .A2(KEYINPUT55), .A3(new_n528_), .A4(new_n524_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n541_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT56), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n741_), .B1(new_n750_), .B2(KEYINPUT114), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n749_), .B1(new_n748_), .B2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n222_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n213_), .B1(new_n217_), .B2(new_n211_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n216_), .A2(new_n755_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n219_), .A2(new_n222_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n751_), .A2(new_n753_), .B1(new_n543_), .B2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n740_), .B1(new_n758_), .B2(new_n604_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n741_), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n748_), .A2(new_n749_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n753_), .B(new_n760_), .C1(new_n761_), .C2(new_n752_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n543_), .A2(new_n757_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(KEYINPUT57), .A3(new_n603_), .ZN(new_n765_));
  AOI211_X1 g564(.A(KEYINPUT56), .B(new_n541_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n542_), .A2(KEYINPUT115), .A3(new_n757_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT115), .B1(new_n542_), .B2(new_n757_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n750_), .A2(new_n766_), .A3(new_n769_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n646_), .B(KEYINPUT116), .C1(new_n770_), .C2(KEYINPUT58), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(KEYINPUT58), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n769_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n748_), .A2(new_n749_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n761_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT58), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT116), .B1(new_n778_), .B2(new_n646_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n759_), .B(new_n765_), .C1(new_n773_), .C2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n750_), .A2(new_n766_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT58), .B1(new_n784_), .B2(new_n774_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n783_), .B1(new_n785_), .B2(new_n578_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(new_n772_), .A3(new_n771_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n787_), .A2(KEYINPUT117), .A3(new_n759_), .A4(new_n765_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n782_), .A2(new_n788_), .A3(new_n602_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n578_), .A2(new_n594_), .A3(new_n224_), .A4(new_n547_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n790_), .B(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n694_), .A2(new_n615_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n405_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n739_), .B1(new_n794_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n796_), .A2(KEYINPUT59), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n759_), .A2(new_n765_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n594_), .B1(new_n801_), .B2(new_n787_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n799_), .B(new_n800_), .C1(new_n802_), .C2(new_n792_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n792_), .B1(new_n780_), .B2(new_n602_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n797_), .A2(new_n739_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT118), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT119), .B1(new_n798_), .B2(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n803_), .A2(new_n806_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n594_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n792_), .B1(new_n811_), .B2(new_n788_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT59), .B1(new_n812_), .B2(new_n796_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n809_), .A2(new_n810_), .A3(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n808_), .A2(new_n223_), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(G113gat), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n812_), .A2(new_n796_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  OR3_X1    g617(.A1(new_n818_), .A2(G113gat), .A3(new_n224_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n816_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n816_), .A2(KEYINPUT120), .A3(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1340gat));
  NAND3_X1  g623(.A1(new_n809_), .A2(new_n548_), .A3(new_n813_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT121), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n547_), .A2(G120gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n817_), .B1(KEYINPUT60), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n825_), .A2(KEYINPUT121), .ZN(new_n830_));
  OAI21_X1  g629(.A(G120gat), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(KEYINPUT60), .B2(new_n828_), .ZN(G1341gat));
  NAND3_X1  g631(.A1(new_n808_), .A2(new_n594_), .A3(new_n814_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G127gat), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n602_), .A2(G127gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n818_), .B2(new_n835_), .ZN(G1342gat));
  AOI21_X1  g635(.A(G134gat), .B1(new_n817_), .B2(new_n604_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n808_), .A2(new_n814_), .A3(G134gat), .A4(new_n646_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT123), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n839_), .A2(new_n843_), .A3(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1343gat));
  NOR3_X1   g644(.A1(new_n812_), .A2(new_n625_), .A3(new_n347_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n795_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n224_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(new_n243_), .ZN(G1344gat));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n547_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(new_n244_), .ZN(G1345gat));
  NOR2_X1   g650(.A1(new_n847_), .A2(new_n602_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT61), .B(G155gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1346gat));
  INV_X1    g653(.A(G162gat), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n847_), .A2(new_n855_), .A3(new_n578_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n847_), .B2(new_n603_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n857_), .A2(KEYINPUT124), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(KEYINPUT124), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n856_), .B1(new_n858_), .B2(new_n859_), .ZN(G1347gat));
  NAND2_X1  g659(.A1(new_n615_), .A2(new_n347_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n598_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n804_), .A2(new_n458_), .A3(new_n863_), .ZN(new_n864_));
  AND4_X1   g663(.A1(new_n223_), .A2(new_n864_), .A3(new_n419_), .A4(new_n420_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n223_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n866_), .A2(KEYINPUT125), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(KEYINPUT125), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(G169gat), .A3(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n865_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n870_), .B2(new_n869_), .ZN(G1348gat));
  AOI21_X1  g671(.A(G176gat), .B1(new_n864_), .B2(new_n548_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n812_), .A2(new_n458_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n863_), .A2(new_n327_), .A3(new_n547_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(G1349gat));
  NAND3_X1  g675(.A1(new_n874_), .A2(new_n594_), .A3(new_n862_), .ZN(new_n877_));
  INV_X1    g676(.A(G183gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n602_), .A2(new_n311_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n877_), .A2(new_n878_), .B1(new_n864_), .B2(new_n879_), .ZN(G1350gat));
  NAND2_X1  g679(.A1(new_n864_), .A2(new_n646_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(G190gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n864_), .A2(new_n312_), .A3(new_n604_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1351gat));
  AND3_X1   g683(.A1(new_n846_), .A2(new_n303_), .A3(new_n615_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n223_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n548_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n351_), .A2(KEYINPUT127), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1353gat));
  NAND2_X1  g689(.A1(new_n885_), .A2(new_n594_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  AND2_X1   g691(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n891_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n891_), .B2(new_n892_), .ZN(G1354gat));
  INV_X1    g694(.A(G218gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n885_), .A2(new_n896_), .A3(new_n604_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n885_), .A2(new_n646_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n896_), .ZN(G1355gat));
endmodule


