//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(G225gat), .A2(G233gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(G127gat), .B(G134gat), .Z(new_n210_));
  INV_X1    g009(.A(KEYINPUT85), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G127gat), .B(G134gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(KEYINPUT85), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n209_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n211_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(KEYINPUT85), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(new_n208_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225_));
  AND2_X1   g024(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n226_));
  NOR2_X1   g025(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT87), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT88), .B1(new_n225_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT88), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n232_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G141gat), .ZN(new_n235_));
  INV_X1    g034(.A(G148gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT89), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT2), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(KEYINPUT89), .A2(KEYINPUT2), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n237_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  OAI22_X1  g041(.A1(new_n238_), .A2(new_n239_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n234_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n224_), .B1(new_n229_), .B2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n222_), .B1(KEYINPUT1), .B2(new_n220_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n220_), .A2(KEYINPUT1), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NOR3_X1   g047(.A1(new_n248_), .A2(new_n225_), .A3(new_n237_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n219_), .B1(new_n245_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT87), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n228_), .B(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n234_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n223_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n249_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n215_), .A2(new_n218_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n250_), .A2(KEYINPUT97), .A3(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n245_), .A2(new_n249_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT97), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(new_n260_), .A3(new_n256_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n207_), .B1(new_n258_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT98), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n258_), .A2(KEYINPUT4), .A3(new_n261_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n250_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n207_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n205_), .B1(new_n264_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n258_), .A2(new_n261_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n206_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n263_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n262_), .A2(KEYINPUT98), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n269_), .A2(new_n273_), .A3(new_n205_), .A4(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n270_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G197gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT91), .B1(new_n278_), .B2(G204gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT91), .ZN(new_n280_));
  INV_X1    g079(.A(G204gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(G197gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n278_), .A2(G204gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G211gat), .B(G218gat), .Z(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(KEYINPUT21), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(G197gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n283_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT21), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G211gat), .B(G218gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n284_), .A2(KEYINPUT21), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n286_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT29), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n293_), .B1(new_n259_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G228gat), .ZN(new_n296_));
  INV_X1    g095(.A(G233gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT92), .B1(new_n295_), .B2(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n284_), .A2(KEYINPUT21), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n285_), .B1(KEYINPUT21), .B2(new_n288_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n285_), .A2(KEYINPUT21), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n300_), .A2(new_n301_), .B1(new_n302_), .B2(new_n284_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n254_), .A2(new_n255_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n304_), .B2(KEYINPUT29), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT92), .ZN(new_n306_));
  INV_X1    g105(.A(new_n298_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n299_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT93), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n295_), .A2(new_n310_), .A3(new_n298_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT93), .B1(new_n305_), .B2(new_n307_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n309_), .A2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n259_), .A2(new_n294_), .A3(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n304_), .B2(KEYINPUT29), .ZN(new_n318_));
  XOR2_X1   g117(.A(G22gat), .B(G50gat), .Z(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n317_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G78gat), .B(G106gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n320_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n322_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(KEYINPUT94), .ZN(new_n326_));
  INV_X1    g125(.A(new_n324_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(new_n321_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n314_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n309_), .A2(new_n313_), .ZN(new_n330_));
  OAI211_X1 g129(.A(KEYINPUT94), .B(new_n323_), .C1(new_n322_), .C2(new_n324_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n327_), .A2(new_n321_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n330_), .B(new_n331_), .C1(new_n323_), .C2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT20), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT22), .B(G169gat), .ZN(new_n336_));
  INV_X1    g135(.A(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n338_), .B(new_n339_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT25), .B(G183gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT26), .B(G190gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n340_), .B(KEYINPUT23), .ZN(new_n348_));
  INV_X1    g147(.A(G169gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n337_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n350_), .A2(KEYINPUT24), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(KEYINPUT24), .A3(new_n339_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n347_), .A2(new_n348_), .A3(new_n351_), .A4(new_n352_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n344_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n335_), .B1(new_n354_), .B2(new_n303_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT22), .B1(new_n349_), .B2(KEYINPUT84), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT22), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G169gat), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n356_), .B(new_n337_), .C1(KEYINPUT84), .C2(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n359_), .B(new_n339_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n353_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT95), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n361_), .A2(new_n293_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n361_), .B2(new_n293_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n355_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT19), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n300_), .A2(new_n301_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n369_), .A2(new_n360_), .A3(new_n353_), .A4(new_n286_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n344_), .A2(new_n353_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n293_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n372_), .A3(KEYINPUT20), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n373_), .A2(new_n367_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G8gat), .B(G36gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n375_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n367_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n355_), .B(new_n382_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n373_), .A2(new_n367_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n380_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n381_), .A2(KEYINPUT99), .A3(KEYINPUT27), .A4(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT99), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(KEYINPUT27), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n385_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT27), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n383_), .A2(new_n385_), .A3(new_n384_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n385_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n392_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n387_), .A2(new_n391_), .A3(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n277_), .A2(new_n334_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n269_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n205_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n275_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n383_), .A2(new_n384_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n385_), .A2(KEYINPUT32), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n403_), .B2(new_n375_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n393_), .A2(new_n394_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n271_), .A2(new_n207_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n399_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n207_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n406_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n410_), .B1(new_n275_), .B2(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n264_), .A2(KEYINPUT33), .A3(new_n205_), .A4(new_n269_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n401_), .A2(new_n405_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n397_), .B1(new_n414_), .B2(new_n334_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G71gat), .B(G99gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(G43gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n361_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(new_n256_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G227gat), .A2(G233gat), .ZN(new_n420_));
  INV_X1    g219(.A(G15gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT30), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT31), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n419_), .B(new_n424_), .Z(new_n425_));
  INV_X1    g224(.A(new_n396_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(new_n334_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n401_), .A2(new_n425_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n415_), .A2(new_n425_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT68), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT67), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT8), .ZN(new_n432_));
  NOR2_X1   g231(.A1(G99gat), .A2(G106gat), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT7), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(G99gat), .B2(G106gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G99gat), .A2(G106gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n439_), .A2(KEYINPUT6), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n435_), .B(new_n436_), .C1(new_n438_), .C2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G85gat), .ZN(new_n442_));
  INV_X1    g241(.A(G92gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G85gat), .A2(G92gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n432_), .B1(new_n441_), .B2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n446_), .A2(KEYINPUT8), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n435_), .A2(new_n436_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n439_), .A2(KEYINPUT6), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n437_), .A2(G99gat), .A3(G106gat), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n452_), .A2(new_n453_), .A3(KEYINPUT65), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT65), .B1(new_n452_), .B2(new_n453_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n451_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT66), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n450_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n451_), .B(KEYINPUT66), .C1(new_n454_), .C2(new_n455_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n448_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT9), .ZN(new_n461_));
  INV_X1    g260(.A(new_n445_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n461_), .B(new_n444_), .C1(new_n462_), .C2(KEYINPUT64), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT64), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n444_), .A2(new_n464_), .A3(KEYINPUT9), .A4(new_n445_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT10), .B(G99gat), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n463_), .B(new_n465_), .C1(G106gat), .C2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n454_), .A2(new_n455_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n431_), .B1(new_n460_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n448_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n435_), .A2(new_n436_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT65), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n473_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n452_), .A2(new_n453_), .A3(KEYINPUT65), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n472_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n449_), .B1(new_n476_), .B2(KEYINPUT66), .ZN(new_n477_));
  INV_X1    g276(.A(new_n459_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n471_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n469_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(KEYINPUT67), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G57gat), .B(G64gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT11), .ZN(new_n483_));
  XOR2_X1   g282(.A(G71gat), .B(G78gat), .Z(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n482_), .A2(KEYINPUT11), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n483_), .A2(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n470_), .A2(new_n481_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n479_), .A2(new_n480_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n489_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(KEYINPUT12), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n489_), .B1(new_n470_), .B2(new_n481_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n490_), .B(new_n493_), .C1(new_n494_), .C2(KEYINPUT12), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G230gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n430_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT67), .B1(new_n479_), .B2(new_n480_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n456_), .A2(new_n457_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(new_n459_), .A3(new_n449_), .ZN(new_n501_));
  AOI211_X1 g300(.A(new_n431_), .B(new_n469_), .C1(new_n501_), .C2(new_n471_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n492_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n490_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n497_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n490_), .A2(new_n493_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT12), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n506_), .A2(new_n508_), .A3(KEYINPUT68), .A4(new_n496_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n498_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G120gat), .B(G148gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT5), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G176gat), .B(G204gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n514_), .B(KEYINPUT69), .Z(new_n515_));
  NAND2_X1  g314(.A1(new_n510_), .A2(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n498_), .A2(new_n509_), .A3(new_n505_), .A4(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n518_), .A2(KEYINPUT13), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT13), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT76), .B(G1gat), .ZN(new_n523_));
  INV_X1    g322(.A(G8gat), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT14), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G1gat), .B(G8gat), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n527_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G29gat), .B(G36gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G43gat), .B(G50gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n530_), .B(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n537_), .A2(KEYINPUT80), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n530_), .A2(new_n533_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT15), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n533_), .B(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n539_), .B1(new_n541_), .B2(new_n530_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n537_), .B(KEYINPUT80), .C1(new_n536_), .C2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G113gat), .B(G141gat), .Z(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT82), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G169gat), .B(G197gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n544_), .A2(KEYINPUT81), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n544_), .B1(KEYINPUT81), .B2(new_n549_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n552_), .A2(KEYINPUT83), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(KEYINPUT83), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NOR3_X1   g354(.A1(new_n429_), .A2(new_n522_), .A3(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G190gat), .B(G218gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G134gat), .B(G162gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n559_), .B(KEYINPUT36), .Z(new_n560_));
  NAND2_X1  g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT34), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT35), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n469_), .B1(new_n501_), .B2(new_n471_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT70), .B1(new_n564_), .B2(new_n541_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n533_), .B(KEYINPUT15), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT70), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n566_), .B(new_n567_), .C1(new_n460_), .C2(new_n469_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n565_), .A2(KEYINPUT71), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT71), .B1(new_n565_), .B2(new_n568_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n470_), .A2(new_n481_), .A3(new_n533_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n470_), .A2(new_n481_), .A3(KEYINPUT72), .A4(new_n533_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n563_), .B1(new_n571_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n563_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n562_), .A2(KEYINPUT35), .ZN(new_n579_));
  AOI211_X1 g378(.A(new_n578_), .B(new_n579_), .C1(new_n565_), .C2(new_n568_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n560_), .B1(new_n577_), .B2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n574_), .A2(new_n575_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT71), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n567_), .B1(new_n491_), .B2(new_n566_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n564_), .A2(KEYINPUT70), .A3(new_n541_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n565_), .A2(KEYINPUT71), .A3(new_n568_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n578_), .B1(new_n584_), .B2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n559_), .A2(KEYINPUT36), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n581_), .A3(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n583_), .A2(new_n593_), .A3(KEYINPUT73), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT74), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT73), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n591_), .A2(new_n596_), .A3(new_n581_), .A4(new_n592_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n594_), .A2(new_n595_), .A3(KEYINPUT37), .A4(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(KEYINPUT75), .B1(new_n577_), .B2(new_n582_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT75), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n591_), .A2(new_n600_), .A3(new_n581_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n599_), .A2(new_n601_), .A3(new_n560_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n603_), .A3(new_n593_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n597_), .A2(KEYINPUT37), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n595_), .B1(new_n607_), .B2(new_n594_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT77), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n489_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(new_n530_), .ZN(new_n613_));
  XOR2_X1   g412(.A(G127gat), .B(G155gat), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT16), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT17), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n613_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT79), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n613_), .A2(new_n621_), .A3(new_n617_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT78), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n620_), .B(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n609_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n556_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n523_), .A3(new_n401_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n522_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n625_), .A3(new_n552_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n602_), .A2(new_n593_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n429_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G1gat), .B1(new_n639_), .B2(new_n277_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n630_), .A2(new_n631_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n632_), .A2(new_n640_), .A3(new_n641_), .ZN(G1324gat));
  NAND3_X1  g441(.A1(new_n629_), .A2(new_n524_), .A3(new_n426_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n639_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n426_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  AND4_X1   g445(.A1(KEYINPUT100), .A2(new_n645_), .A3(new_n646_), .A4(G8gat), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n524_), .B1(new_n648_), .B2(KEYINPUT39), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n645_), .A2(new_n649_), .B1(KEYINPUT100), .B2(new_n646_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n643_), .B1(new_n647_), .B2(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g451(.A(G15gat), .B1(new_n639_), .B2(new_n425_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT41), .Z(new_n654_));
  INV_X1    g453(.A(new_n425_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n629_), .A2(new_n421_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1326gat));
  INV_X1    g456(.A(new_n334_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G22gat), .B1(new_n639_), .B2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n658_), .A2(G22gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n661_), .B1(new_n628_), .B2(new_n662_), .ZN(G1327gat));
  NOR2_X1   g462(.A1(new_n636_), .A2(new_n625_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n556_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G29gat), .B1(new_n665_), .B2(new_n401_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n583_), .A2(new_n593_), .A3(KEYINPUT73), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT74), .B1(new_n667_), .B2(new_n606_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(new_n604_), .A3(new_n598_), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT43), .B1(new_n429_), .B2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n405_), .B1(new_n270_), .B2(new_n276_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n275_), .A2(new_n411_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n410_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n413_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n334_), .B1(new_n671_), .B2(new_n674_), .ZN(new_n675_));
  AND4_X1   g474(.A1(new_n275_), .A2(new_n334_), .A3(new_n396_), .A4(new_n400_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n425_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n427_), .A2(new_n428_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n609_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n670_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n633_), .A2(new_n626_), .A3(new_n552_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(KEYINPUT102), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n683_), .B1(new_n670_), .B2(new_n681_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(KEYINPUT44), .ZN(new_n690_));
  AOI22_X1  g489(.A1(new_n687_), .A2(new_n690_), .B1(KEYINPUT44), .B2(new_n689_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n401_), .A2(G29gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n666_), .B1(new_n691_), .B2(new_n692_), .ZN(G1328gat));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT105), .B1(new_n694_), .B2(KEYINPUT46), .ZN(new_n695_));
  NOR2_X1   g494(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n696_));
  INV_X1    g495(.A(new_n665_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n396_), .A2(G36gat), .ZN(new_n698_));
  OR3_X1    g497(.A1(new_n697_), .A2(KEYINPUT45), .A3(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT45), .B1(new_n697_), .B2(new_n698_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n687_), .A2(new_n690_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n396_), .B1(new_n689_), .B2(KEYINPUT44), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n702_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n703_), .B1(new_n702_), .B2(new_n704_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n695_), .B(new_n701_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT102), .B1(new_n685_), .B2(new_n686_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n689_), .A2(new_n688_), .A3(KEYINPUT44), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n704_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT103), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(G36gat), .A3(new_n705_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n695_), .B1(new_n714_), .B2(new_n701_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n709_), .A2(new_n715_), .ZN(G1329gat));
  NAND3_X1  g515(.A1(new_n691_), .A2(G43gat), .A3(new_n655_), .ZN(new_n717_));
  INV_X1    g516(.A(G43gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n697_), .B2(new_n425_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1330gat));
  OR3_X1    g521(.A1(new_n697_), .A2(G50gat), .A3(new_n658_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n691_), .A2(new_n334_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(KEYINPUT107), .ZN(new_n725_));
  OAI21_X1  g524(.A(G50gat), .B1(new_n724_), .B2(KEYINPUT107), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n723_), .B1(new_n725_), .B2(new_n726_), .ZN(G1331gat));
  NAND4_X1  g526(.A1(new_n638_), .A2(new_n625_), .A3(new_n522_), .A4(new_n555_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G57gat), .B1(new_n728_), .B2(new_n277_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n552_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n522_), .A2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n429_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n627_), .A2(new_n732_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n277_), .A2(G57gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n733_), .B2(new_n734_), .ZN(G1332gat));
  OAI21_X1  g534(.A(G64gat), .B1(new_n728_), .B2(new_n396_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT48), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n396_), .A2(G64gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n733_), .B2(new_n738_), .ZN(G1333gat));
  OAI21_X1  g538(.A(G71gat), .B1(new_n728_), .B2(new_n425_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT49), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n425_), .A2(G71gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n733_), .B2(new_n742_), .ZN(G1334gat));
  OAI21_X1  g542(.A(G78gat), .B1(new_n728_), .B2(new_n658_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n658_), .A2(G78gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n733_), .B2(new_n747_), .ZN(G1335gat));
  NAND2_X1  g547(.A1(new_n732_), .A2(new_n664_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G85gat), .B1(new_n750_), .B2(new_n401_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n522_), .A2(new_n626_), .A3(new_n730_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n682_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT109), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n682_), .A2(new_n753_), .A3(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n401_), .A2(G85gat), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT110), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n751_), .B1(new_n758_), .B2(new_n760_), .ZN(G1336gat));
  NAND3_X1  g560(.A1(new_n750_), .A2(new_n443_), .A3(new_n426_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n396_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n443_), .ZN(G1337gat));
  NOR3_X1   g563(.A1(new_n749_), .A2(new_n466_), .A3(new_n425_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n756_), .B1(new_n682_), .B2(new_n753_), .ZN(new_n766_));
  AOI211_X1 g565(.A(KEYINPUT109), .B(new_n752_), .C1(new_n670_), .C2(new_n681_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n655_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n765_), .B1(new_n768_), .B2(G99gat), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT112), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT51), .B1(new_n769_), .B2(KEYINPUT111), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n773_), .B(new_n765_), .C1(new_n768_), .C2(G99gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n771_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n765_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n425_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n777_));
  INV_X1    g576(.A(G99gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n776_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n773_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n769_), .A2(KEYINPUT111), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n780_), .A2(KEYINPUT112), .A3(new_n781_), .A4(KEYINPUT51), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n775_), .A2(new_n782_), .ZN(G1338gat));
  OAI21_X1  g582(.A(G106gat), .B1(new_n754_), .B2(new_n658_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT52), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n658_), .A2(G106gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n749_), .B2(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g587(.A1(new_n427_), .A2(new_n655_), .A3(new_n401_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n535_), .B1(new_n542_), .B2(KEYINPUT118), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(KEYINPUT118), .B2(new_n542_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n548_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n790_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n792_), .A2(new_n790_), .A3(new_n793_), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n794_), .B(new_n795_), .C1(new_n548_), .C2(new_n544_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n518_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n552_), .A2(new_n517_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n506_), .A2(new_n508_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n470_), .A2(new_n481_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT12), .B1(new_n801_), .B2(new_n492_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n490_), .A2(new_n493_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT115), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n800_), .A2(new_n804_), .A3(new_n497_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n506_), .A2(new_n508_), .A3(KEYINPUT55), .A4(new_n496_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT116), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n802_), .A2(new_n803_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(KEYINPUT55), .A4(new_n496_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n805_), .A2(new_n807_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n498_), .A2(new_n812_), .A3(new_n509_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n515_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n498_), .A2(new_n812_), .A3(new_n509_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n817_), .A2(new_n810_), .A3(new_n805_), .A4(new_n807_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(KEYINPUT56), .A3(new_n515_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n798_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n797_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  AOI211_X1 g621(.A(KEYINPUT117), .B(new_n798_), .C1(new_n816_), .C2(new_n819_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n636_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(KEYINPUT57), .B(new_n636_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n816_), .A2(new_n819_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n796_), .A2(new_n517_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n830_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n828_), .B1(new_n833_), .B2(new_n669_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(KEYINPUT58), .A3(new_n832_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n818_), .A2(KEYINPUT56), .A3(new_n515_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT56), .B1(new_n818_), .B2(new_n515_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n832_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n829_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n609_), .A3(KEYINPUT121), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n834_), .A2(new_n835_), .A3(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n826_), .A2(new_n827_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n626_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n553_), .A2(new_n625_), .A3(new_n554_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n522_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n846_), .B2(new_n669_), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n847_), .A2(KEYINPUT114), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(new_n669_), .A3(new_n844_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n849_), .A2(KEYINPUT113), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(KEYINPUT114), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(KEYINPUT113), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n848_), .A2(new_n850_), .A3(new_n851_), .A4(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n789_), .B1(new_n843_), .B2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(G113gat), .B1(new_n854_), .B2(new_n552_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n843_), .A2(new_n853_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n789_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n860_));
  NAND3_X1  g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n854_), .A2(KEYINPUT123), .A3(new_n860_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n857_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(G113gat), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n555_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n855_), .B1(new_n865_), .B2(new_n867_), .ZN(G1340gat));
  INV_X1    g667(.A(G120gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n633_), .B2(KEYINPUT60), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n854_), .B(new_n870_), .C1(KEYINPUT60), .C2(new_n869_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n522_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n873_), .B2(new_n869_), .ZN(G1341gat));
  AOI21_X1  g673(.A(G127gat), .B1(new_n854_), .B2(new_n625_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n625_), .A2(G127gat), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n865_), .B2(new_n876_), .ZN(G1342gat));
  AOI21_X1  g676(.A(G134gat), .B1(new_n854_), .B2(new_n637_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n609_), .A2(G134gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n865_), .B2(new_n879_), .ZN(G1343gat));
  NOR3_X1   g679(.A1(new_n658_), .A2(new_n277_), .A3(new_n655_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n858_), .A2(new_n396_), .A3(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n730_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n235_), .ZN(G1344gat));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n633_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n236_), .ZN(G1345gat));
  NOR2_X1   g685(.A1(new_n882_), .A2(new_n626_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT61), .B(G155gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  OAI21_X1  g688(.A(G162gat), .B1(new_n882_), .B2(new_n669_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n636_), .A2(G162gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n882_), .B2(new_n891_), .ZN(G1347gat));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n428_), .A2(new_n658_), .A3(new_n426_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n843_), .B2(new_n853_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n552_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n893_), .B1(new_n896_), .B2(G169gat), .ZN(new_n897_));
  AOI211_X1 g696(.A(KEYINPUT62), .B(new_n349_), .C1(new_n895_), .C2(new_n552_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n895_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n552_), .A2(new_n336_), .ZN(new_n900_));
  XOR2_X1   g699(.A(new_n900_), .B(KEYINPUT124), .Z(new_n901_));
  OAI22_X1  g700(.A1(new_n897_), .A2(new_n898_), .B1(new_n899_), .B2(new_n901_), .ZN(G1348gat));
  XNOR2_X1  g701(.A(KEYINPUT125), .B(G176gat), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n337_), .A2(KEYINPUT125), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n895_), .A2(new_n522_), .ZN(new_n905_));
  MUX2_X1   g704(.A(new_n903_), .B(new_n904_), .S(new_n905_), .Z(G1349gat));
  NAND2_X1  g705(.A1(new_n895_), .A2(new_n625_), .ZN(new_n907_));
  MUX2_X1   g706(.A(new_n345_), .B(G183gat), .S(new_n907_), .Z(G1350gat));
  NAND3_X1  g707(.A1(new_n895_), .A2(new_n637_), .A3(new_n346_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(G190gat), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(new_n895_), .B2(new_n609_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT126), .B1(new_n910_), .B2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n912_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n914_), .A2(new_n915_), .A3(new_n909_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n913_), .A2(new_n916_), .ZN(G1351gat));
  NOR4_X1   g716(.A1(new_n658_), .A2(new_n401_), .A3(new_n655_), .A4(new_n396_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n858_), .A2(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G197gat), .B1(new_n919_), .B2(new_n552_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n858_), .A2(G197gat), .A3(new_n552_), .A4(new_n918_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n921_), .A2(KEYINPUT127), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n921_), .A2(KEYINPUT127), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n920_), .A2(new_n922_), .A3(new_n923_), .ZN(G1352gat));
  NAND2_X1  g723(.A1(new_n919_), .A2(new_n522_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g725(.A(KEYINPUT63), .B(G211gat), .C1(new_n919_), .C2(new_n625_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT63), .B(G211gat), .Z(new_n928_));
  AND3_X1   g727(.A1(new_n919_), .A2(new_n625_), .A3(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1354gat));
  INV_X1    g729(.A(G218gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n919_), .A2(new_n931_), .A3(new_n637_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n919_), .A2(new_n609_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(new_n931_), .ZN(G1355gat));
endmodule


