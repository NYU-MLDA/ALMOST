//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT26), .B(G190gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT90), .Z(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT25), .B(G183gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT79), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT24), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n208_), .B(KEYINPUT79), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT23), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n207_), .A2(new_n212_), .A3(new_n215_), .A4(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n217_), .B1(G183gat), .B2(G190gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT22), .B(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n219_), .A2(new_n214_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G204gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT83), .B1(new_n224_), .B2(G197gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT83), .ZN(new_n226_));
  INV_X1    g025(.A(G197gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(G204gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT21), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n224_), .A2(G197gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n225_), .A2(new_n228_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n224_), .A2(G197gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n227_), .A2(G204gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT21), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G218gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G211gat), .ZN(new_n236_));
  INV_X1    g035(.A(G211gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G218gat), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n231_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n225_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n229_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n218_), .A2(new_n223_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n245_));
  INV_X1    g044(.A(G169gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT22), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n246_), .A2(KEYINPUT22), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n221_), .B(new_n247_), .C1(new_n248_), .C2(new_n245_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n219_), .A2(new_n214_), .A3(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n215_), .A2(new_n212_), .A3(new_n217_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT78), .ZN(new_n252_));
  INV_X1    g051(.A(G183gat), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n253_), .A2(KEYINPUT25), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n204_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n206_), .A2(KEYINPUT78), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n250_), .B1(new_n251_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n240_), .A2(new_n243_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT20), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n203_), .B1(new_n244_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT20), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n262_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n203_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n218_), .A2(new_n223_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n263_), .B(new_n264_), .C1(new_n265_), .C2(new_n259_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G8gat), .B(G36gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G64gat), .B(G92gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n261_), .A2(new_n266_), .A3(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n272_), .A2(KEYINPUT27), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n244_), .A2(new_n260_), .A3(new_n203_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT85), .B1(new_n240_), .B2(new_n243_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n240_), .A2(new_n243_), .A3(KEYINPUT85), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n218_), .A2(new_n276_), .A3(new_n277_), .A4(new_n223_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n264_), .B1(new_n278_), .B2(new_n263_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n271_), .B(KEYINPUT95), .Z(new_n281_));
  OAI211_X1 g080(.A(new_n273_), .B(KEYINPUT96), .C1(new_n280_), .C2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G225gat), .A2(G233gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n285_));
  XOR2_X1   g084(.A(G127gat), .B(G134gat), .Z(new_n286_));
  XOR2_X1   g085(.A(G113gat), .B(G120gat), .Z(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G127gat), .B(G134gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G113gat), .B(G120gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT81), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n288_), .A2(KEYINPUT81), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT3), .ZN(new_n296_));
  INV_X1    g095(.A(G141gat), .ZN(new_n297_));
  INV_X1    g096(.A(G148gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT2), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n299_), .A2(new_n302_), .A3(new_n303_), .A4(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(KEYINPUT1), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(G155gat), .A3(G162gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n312_), .A3(new_n306_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G141gat), .B(G148gat), .Z(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n294_), .A2(new_n295_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n292_), .A2(KEYINPUT93), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n305_), .A2(new_n308_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT93), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n288_), .A2(new_n320_), .A3(new_n291_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n285_), .B1(new_n317_), .B2(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n317_), .A2(new_n285_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n284_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n317_), .A2(new_n322_), .A3(new_n283_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G1gat), .B(G29gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(G85gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT0), .B(G57gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n331_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(KEYINPUT27), .B(new_n272_), .C1(new_n280_), .C2(new_n281_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT96), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT27), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n261_), .A2(new_n266_), .A3(new_n271_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n271_), .B1(new_n261_), .B2(new_n266_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n282_), .A2(new_n335_), .A3(new_n338_), .A4(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G78gat), .B(G106gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G228gat), .A2(G233gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT82), .Z(new_n346_));
  INV_X1    g145(.A(KEYINPUT84), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n316_), .A2(new_n347_), .A3(KEYINPUT29), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT84), .B1(new_n319_), .B2(new_n349_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n276_), .A2(new_n277_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n346_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n259_), .A2(new_n346_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n319_), .A2(new_n349_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n344_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n357_));
  OR3_X1    g156(.A1(new_n316_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT28), .B1(new_n316_), .B2(KEYINPUT29), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G22gat), .B(G50gat), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n277_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n350_), .B(new_n348_), .C1(new_n364_), .C2(new_n275_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n346_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n344_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n356_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n357_), .A2(new_n363_), .A3(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT89), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  OAI211_X1 g173(.A(KEYINPUT87), .B(new_n344_), .C1(new_n353_), .C2(new_n356_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT87), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n356_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n376_), .B1(new_n377_), .B2(new_n368_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(KEYINPUT86), .A3(new_n368_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n374_), .A2(new_n375_), .A3(new_n378_), .A4(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n381_));
  INV_X1    g180(.A(new_n363_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n372_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G71gat), .B(G99gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(G43gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n258_), .B(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n294_), .A2(new_n295_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G227gat), .A2(G233gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n391_), .B(G15gat), .Z(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT30), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT31), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n388_), .A2(new_n389_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n390_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n394_), .B1(new_n390_), .B2(new_n395_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n385_), .A2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n372_), .B(new_n398_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n343_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n327_), .B2(new_n331_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n325_), .A2(KEYINPUT33), .A3(new_n326_), .A4(new_n333_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n317_), .A2(new_n322_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT94), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n283_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n407_), .B2(new_n406_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n283_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n331_), .A3(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n404_), .A2(new_n405_), .A3(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT92), .B1(new_n340_), .B2(new_n341_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n261_), .A2(new_n266_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n271_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT92), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(new_n272_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n412_), .B1(new_n413_), .B2(new_n418_), .ZN(new_n419_));
  OAI211_X1 g218(.A(KEYINPUT32), .B(new_n271_), .C1(new_n274_), .C2(new_n279_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n271_), .A2(KEYINPUT32), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n261_), .A2(new_n266_), .A3(new_n421_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n420_), .B(new_n422_), .C1(new_n332_), .C2(new_n334_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n399_), .B1(new_n419_), .B2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(new_n385_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n402_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G57gat), .B(G64gat), .ZN(new_n428_));
  INV_X1    g227(.A(G78gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(G71gat), .ZN(new_n430_));
  INV_X1    g229(.A(G71gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(G78gat), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n428_), .A2(KEYINPUT11), .A3(new_n430_), .A4(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(G64gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(G57gat), .ZN(new_n435_));
  INV_X1    g234(.A(G57gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G64gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n437_), .A3(KEYINPUT11), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n430_), .A2(new_n432_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n428_), .A2(KEYINPUT11), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n433_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n443_));
  INV_X1    g242(.A(G106gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT65), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G99gat), .A2(G106gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT9), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(G85gat), .A3(G92gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n450_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G85gat), .ZN(new_n455_));
  INV_X1    g254(.A(G92gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G85gat), .A2(G92gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(KEYINPUT9), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT65), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n443_), .A2(new_n460_), .A3(new_n444_), .A4(new_n445_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n447_), .A2(new_n454_), .A3(new_n459_), .A4(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT7), .ZN(new_n463_));
  INV_X1    g262(.A(G99gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(new_n444_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n465_), .A2(new_n450_), .A3(new_n453_), .A4(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT8), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n457_), .A2(new_n458_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n468_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n442_), .B(new_n462_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT66), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n467_), .A2(new_n469_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT8), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT66), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(new_n462_), .A4(new_n442_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n462_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n442_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n473_), .A2(new_n479_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G230gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT64), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT67), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n480_), .A2(new_n487_), .ZN(new_n488_));
  OAI211_X1 g287(.A(KEYINPUT67), .B(new_n462_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n489_));
  OAI211_X1 g288(.A(KEYINPUT12), .B(new_n433_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n488_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT12), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n482_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n485_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n472_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n492_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G120gat), .B(G148gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT5), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G176gat), .B(G204gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n486_), .A2(new_n497_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT68), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n486_), .A2(new_n497_), .A3(KEYINPUT68), .A4(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n486_), .A2(new_n497_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n501_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT13), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n506_), .A2(KEYINPUT13), .A3(new_n509_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G113gat), .B(G141gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G169gat), .B(G197gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT72), .B(G8gat), .ZN(new_n519_));
  INV_X1    g318(.A(G1gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT14), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G1gat), .B(G8gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n521_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G29gat), .B(G36gat), .Z(new_n529_));
  INV_X1    g328(.A(G50gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(G43gat), .ZN(new_n531_));
  INV_X1    g330(.A(G43gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(G50gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n529_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G29gat), .B(G36gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G43gat), .B(G50gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT15), .B1(new_n535_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n535_), .A2(new_n538_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT15), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n528_), .A2(new_n539_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n527_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n524_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n535_), .A2(KEYINPUT75), .A3(new_n538_), .ZN(new_n546_));
  AOI21_X1  g345(.A(KEYINPUT75), .B1(new_n535_), .B2(new_n538_), .ZN(new_n547_));
  OAI22_X1  g346(.A1(new_n544_), .A2(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n543_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n547_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n535_), .A2(KEYINPUT75), .A3(new_n538_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n553_), .A2(new_n526_), .A3(new_n527_), .A4(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n548_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n551_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT76), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n556_), .A2(KEYINPUT76), .A3(new_n551_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n552_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT77), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n518_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n543_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(new_n548_), .A3(new_n550_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT76), .B1(new_n556_), .B2(new_n551_), .ZN(new_n566_));
  AOI211_X1 g365(.A(new_n558_), .B(new_n550_), .C1(new_n548_), .C2(new_n555_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(KEYINPUT77), .A3(new_n517_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n563_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n514_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n427_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT97), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT37), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n542_), .A2(new_n539_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n488_), .A2(new_n576_), .A3(new_n489_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT34), .Z(new_n579_));
  INV_X1    g378(.A(KEYINPUT35), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT69), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n540_), .B(new_n462_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n580_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n577_), .A2(new_n582_), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n582_), .B1(new_n577_), .B2(new_n585_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(KEYINPUT36), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n591_), .B(KEYINPUT36), .Z(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n575_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT37), .B1(new_n588_), .B2(new_n592_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(KEYINPUT70), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT70), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n599_), .B(new_n594_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n597_), .A2(new_n598_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT71), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT71), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n597_), .A2(new_n598_), .A3(new_n603_), .A4(new_n600_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n596_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G127gat), .B(G155gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT16), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT73), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n528_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n442_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n544_), .A2(new_n545_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n611_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n528_), .A2(new_n612_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n481_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OAI211_X1 g420(.A(KEYINPUT17), .B(new_n609_), .C1(new_n621_), .C2(KEYINPUT74), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT17), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n609_), .B1(new_n615_), .B2(new_n619_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT74), .B1(new_n615_), .B2(new_n619_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n609_), .ZN(new_n626_));
  OAI22_X1  g425(.A1(new_n623_), .A2(new_n624_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n622_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n605_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n573_), .A2(new_n574_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n343_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n380_), .A2(new_n382_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT88), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n398_), .B1(new_n636_), .B2(new_n372_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n401_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n632_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n385_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n640_), .B(new_n399_), .C1(new_n424_), .C2(new_n419_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(new_n630_), .A3(new_n571_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT97), .ZN(new_n644_));
  INV_X1    g443(.A(new_n335_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n631_), .A2(new_n644_), .A3(new_n520_), .A4(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT38), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT99), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n598_), .A2(new_n600_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n593_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT98), .B1(new_n427_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT98), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n642_), .A2(new_n654_), .A3(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n571_), .A2(new_n628_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(new_n645_), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G1gat), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n649_), .B(new_n660_), .C1(new_n647_), .C2(new_n646_), .ZN(G1324gat));
  AND2_X1   g460(.A1(new_n338_), .A2(new_n342_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n282_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n656_), .A2(new_n663_), .A3(new_n658_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G8gat), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT39), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n664_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n631_), .A2(new_n644_), .A3(new_n519_), .A4(new_n663_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(KEYINPUT100), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(KEYINPUT100), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n667_), .B(new_n668_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(G1325gat));
  NAND3_X1  g473(.A1(new_n656_), .A2(new_n398_), .A3(new_n658_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n675_), .A2(G15gat), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n675_), .B2(G15gat), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n643_), .A2(G15gat), .A3(new_n399_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT104), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n680_), .A2(new_n681_), .A3(new_n683_), .ZN(G1326gat));
  OR3_X1    g483(.A1(new_n643_), .A2(G22gat), .A3(new_n640_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n656_), .A2(new_n385_), .A3(new_n658_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(new_n687_), .A3(G22gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(G22gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(G1327gat));
  NOR2_X1   g489(.A1(new_n651_), .A2(new_n628_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n573_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n645_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n571_), .A2(new_n629_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n605_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT43), .B1(new_n427_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n698_), .B(new_n605_), .C1(new_n402_), .C2(new_n426_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n695_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT44), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n701_), .A2(G29gat), .A3(new_n645_), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n700_), .A2(KEYINPUT44), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n694_), .B1(new_n702_), .B2(new_n703_), .ZN(G1328gat));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT105), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n705_), .A2(KEYINPUT105), .ZN(new_n707_));
  INV_X1    g506(.A(new_n663_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n692_), .A2(G36gat), .A3(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT45), .ZN(new_n710_));
  INV_X1    g509(.A(G36gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n708_), .B1(new_n700_), .B2(KEYINPUT44), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n703_), .B2(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n706_), .B(new_n707_), .C1(new_n710_), .C2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n703_), .A2(new_n712_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G36gat), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n709_), .B(new_n717_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n716_), .A2(new_n718_), .A3(KEYINPUT105), .A4(new_n705_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n714_), .A2(new_n719_), .ZN(G1329gat));
  XOR2_X1   g519(.A(KEYINPUT106), .B(G43gat), .Z(new_n721_));
  OAI21_X1  g520(.A(new_n721_), .B1(new_n692_), .B2(new_n399_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n703_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n701_), .A2(G43gat), .A3(new_n398_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  XOR2_X1   g524(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n693_), .B2(new_n385_), .ZN(new_n728_));
  AOI211_X1 g527(.A(new_n530_), .B(new_n640_), .C1(new_n700_), .C2(KEYINPUT44), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n703_), .ZN(G1331gat));
  INV_X1    g529(.A(new_n514_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n570_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n642_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n630_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT108), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n436_), .A3(new_n645_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n733_), .A2(new_n628_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(new_n645_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n737_), .B1(new_n740_), .B2(new_n436_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n737_), .B(KEYINPUT109), .C1(new_n436_), .C2(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1332gat));
  NAND3_X1  g544(.A1(new_n736_), .A2(new_n434_), .A3(new_n663_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n739_), .A2(new_n663_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G64gat), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT48), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(KEYINPUT48), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(G1333gat));
  NAND3_X1  g550(.A1(new_n736_), .A2(new_n431_), .A3(new_n398_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n739_), .A2(new_n398_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G71gat), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(KEYINPUT49), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(KEYINPUT49), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(G1334gat));
  NAND3_X1  g556(.A1(new_n736_), .A2(new_n429_), .A3(new_n385_), .ZN(new_n758_));
  AOI211_X1 g557(.A(KEYINPUT50), .B(new_n429_), .C1(new_n739_), .C2(new_n385_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n739_), .A2(new_n385_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(G78gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n758_), .B(KEYINPUT110), .C1(new_n762_), .C2(new_n759_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1335gat));
  NAND2_X1  g566(.A1(new_n734_), .A2(new_n691_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n455_), .A3(new_n645_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n733_), .A2(new_n629_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(new_n645_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n770_), .B1(new_n773_), .B2(new_n455_), .ZN(G1336gat));
  NAND3_X1  g573(.A1(new_n769_), .A2(new_n456_), .A3(new_n663_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n772_), .A2(new_n663_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n456_), .ZN(G1337gat));
  AOI21_X1  g576(.A(new_n464_), .B1(new_n772_), .B2(new_n398_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n398_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n769_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT51), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n780_), .B(new_n782_), .ZN(G1338gat));
  NAND3_X1  g582(.A1(new_n769_), .A2(new_n444_), .A3(new_n385_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  INV_X1    g584(.A(new_n771_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n698_), .B1(new_n642_), .B2(new_n605_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n699_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n385_), .B(new_n786_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n772_), .A2(KEYINPUT112), .A3(new_n385_), .ZN(new_n792_));
  AND4_X1   g591(.A1(new_n785_), .A2(new_n791_), .A3(new_n792_), .A4(G106gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n444_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n785_), .B1(new_n794_), .B2(new_n792_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n784_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT53), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n798_), .B(new_n784_), .C1(new_n793_), .C2(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1339gat));
  AOI22_X1  g599(.A1(new_n563_), .A2(new_n569_), .B1(new_n627_), .B2(new_n622_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n512_), .A2(new_n513_), .A3(new_n801_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n605_), .A2(new_n802_), .A3(KEYINPUT54), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT54), .B1(new_n605_), .B2(new_n802_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(KEYINPUT113), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n806_), .B(KEYINPUT54), .C1(new_n605_), .C2(new_n802_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n543_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n551_), .B1(new_n548_), .B2(new_n555_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n518_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n568_), .A2(new_n517_), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n506_), .A2(new_n509_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n492_), .A2(new_n494_), .A3(new_n473_), .A4(new_n479_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n485_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n492_), .A2(new_n494_), .A3(KEYINPUT55), .A4(new_n496_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n497_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n816_), .A2(new_n817_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n508_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(KEYINPUT56), .A3(new_n508_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n563_), .A2(new_n506_), .A3(new_n569_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n814_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n809_), .B1(new_n827_), .B2(new_n652_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n563_), .A2(new_n506_), .A3(new_n569_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT57), .B(new_n651_), .C1(new_n830_), .C2(new_n814_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n813_), .A2(new_n812_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n820_), .A2(KEYINPUT56), .A3(new_n508_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT56), .B1(new_n820_), .B2(new_n508_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(KEYINPUT58), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n837_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n825_), .A2(new_n832_), .A3(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n605_), .A2(new_n838_), .A3(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n828_), .A2(new_n831_), .A3(new_n841_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n805_), .A2(new_n807_), .B1(new_n629_), .B2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n663_), .A2(new_n335_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n638_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT116), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n804_), .A2(KEYINPUT113), .ZN(new_n847_));
  INV_X1    g646(.A(new_n803_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n807_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n842_), .A2(new_n629_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n638_), .A4(new_n844_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n846_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G113gat), .B1(new_n855_), .B2(new_n732_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n845_), .A2(KEYINPUT59), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n828_), .A2(new_n841_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n827_), .A2(new_n652_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n858_), .A2(new_n859_), .B1(KEYINPUT57), .B2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n828_), .A2(new_n841_), .A3(KEYINPUT117), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n628_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n849_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n857_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT59), .B1(new_n843_), .B2(new_n845_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n732_), .A2(G113gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT118), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n856_), .B1(new_n868_), .B2(new_n870_), .ZN(G1340gat));
  NAND3_X1  g670(.A1(new_n868_), .A2(KEYINPUT120), .A3(new_n514_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT119), .B(G120gat), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n867_), .B2(new_n731_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n872_), .A2(new_n874_), .A3(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n873_), .B1(new_n731_), .B2(KEYINPUT60), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(KEYINPUT60), .B2(new_n873_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n877_), .B1(new_n854_), .B2(new_n879_), .ZN(G1341gat));
  OAI21_X1  g679(.A(G127gat), .B1(new_n867_), .B2(new_n629_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n629_), .A2(G127gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n854_), .B2(new_n882_), .ZN(G1342gat));
  NAND4_X1  g682(.A1(new_n865_), .A2(G134gat), .A3(new_n605_), .A4(new_n866_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n846_), .A2(new_n652_), .A3(new_n853_), .ZN(new_n885_));
  INV_X1    g684(.A(G134gat), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n885_), .A2(KEYINPUT121), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(KEYINPUT121), .B1(new_n885_), .B2(new_n886_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n884_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT122), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n891_), .B(new_n884_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1343gat));
  NOR2_X1   g692(.A1(new_n843_), .A2(new_n400_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n844_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n570_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT123), .B(G141gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1344gat));
  NOR2_X1   g697(.A1(new_n895_), .A2(new_n731_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n298_), .ZN(G1345gat));
  NOR2_X1   g699(.A1(new_n895_), .A2(new_n629_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT61), .B(G155gat), .Z(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  OAI21_X1  g702(.A(G162gat), .B1(new_n895_), .B2(new_n696_), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n651_), .A2(G162gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n895_), .B2(new_n905_), .ZN(G1347gat));
  OR2_X1    g705(.A1(new_n863_), .A2(new_n864_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n708_), .A2(new_n399_), .A3(new_n645_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n385_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n907_), .A2(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(G169gat), .B1(new_n911_), .B2(new_n570_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n911_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n915_), .A2(new_n732_), .A3(new_n220_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n912_), .A2(new_n913_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n914_), .A2(new_n916_), .A3(new_n917_), .ZN(G1348gat));
  AOI21_X1  g717(.A(G176gat), .B1(new_n915_), .B2(new_n514_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n851_), .A2(new_n640_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT124), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n909_), .A2(new_n221_), .A3(new_n731_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n919_), .B1(new_n921_), .B2(new_n922_), .ZN(G1349gat));
  NOR3_X1   g722(.A1(new_n911_), .A2(new_n629_), .A3(new_n206_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n921_), .A2(new_n628_), .A3(new_n908_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n253_), .B2(new_n925_), .ZN(G1350gat));
  OAI211_X1 g725(.A(new_n605_), .B(new_n910_), .C1(new_n863_), .C2(new_n864_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n927_), .A2(new_n928_), .A3(G190gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(G190gat), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n652_), .A2(new_n205_), .ZN(new_n931_));
  OAI22_X1  g730(.A1(new_n929_), .A2(new_n930_), .B1(new_n911_), .B2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(KEYINPUT126), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934_));
  OAI221_X1 g733(.A(new_n934_), .B1(new_n911_), .B2(new_n931_), .C1(new_n929_), .C2(new_n930_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1351gat));
  NOR2_X1   g735(.A1(new_n708_), .A2(new_n645_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n894_), .A2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n570_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(new_n227_), .ZN(G1352gat));
  NOR2_X1   g739(.A1(new_n938_), .A2(new_n731_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(new_n224_), .ZN(G1353gat));
  INV_X1    g741(.A(new_n938_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n629_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(KEYINPUT127), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  XOR2_X1   g746(.A(new_n946_), .B(new_n947_), .Z(G1354gat));
  OAI21_X1  g747(.A(G218gat), .B1(new_n938_), .B2(new_n696_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n652_), .A2(new_n235_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n938_), .B2(new_n950_), .ZN(G1355gat));
endmodule


