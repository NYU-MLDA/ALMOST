//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n954_, new_n956_, new_n957_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_;
  INV_X1    g000(.A(KEYINPUT103), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT85), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204_));
  OAI21_X1  g003(.A(G169gat), .B1(new_n204_), .B2(KEYINPUT82), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n205_), .B(new_n206_), .C1(KEYINPUT82), .C2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT83), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n209_), .A2(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT23), .ZN(new_n213_));
  OR2_X1    g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n213_), .A2(KEYINPUT84), .A3(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT84), .B1(new_n213_), .B2(new_n214_), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n210_), .B(new_n211_), .C1(new_n215_), .C2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  INV_X1    g017(.A(G190gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT80), .B1(new_n219_), .B2(KEYINPUT26), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n218_), .B(new_n220_), .C1(new_n221_), .C2(KEYINPUT80), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT81), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n225_), .A2(KEYINPUT24), .A3(new_n226_), .A4(new_n230_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n222_), .A2(new_n229_), .A3(new_n213_), .A4(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n203_), .B1(new_n217_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT97), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT21), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G197gat), .A2(G204gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT95), .B(G204gat), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n238_), .B1(new_n239_), .B2(G197gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n236_), .B1(new_n237_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT96), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n239_), .A2(G197gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n237_), .B1(G197gat), .B2(G204gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n243_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(KEYINPUT96), .B(new_n245_), .C1(new_n239_), .C2(G197gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT97), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n235_), .B(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(new_n237_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n242_), .A2(new_n249_), .B1(new_n252_), .B2(new_n240_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n217_), .A2(new_n203_), .A3(new_n232_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n234_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT20), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n213_), .A2(new_n214_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT22), .B(G169gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n206_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n230_), .A3(new_n259_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n221_), .A2(new_n218_), .B1(new_n228_), .B2(new_n223_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(new_n213_), .A3(new_n231_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n262_), .A2(KEYINPUT98), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(KEYINPUT98), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n260_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n241_), .A2(new_n237_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n249_), .A2(new_n251_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n252_), .A2(new_n240_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n256_), .B1(new_n265_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n255_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G226gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT19), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G8gat), .B(G36gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT18), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G64gat), .B(G92gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n273_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT20), .ZN(new_n280_));
  INV_X1    g079(.A(new_n265_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n280_), .B1(new_n281_), .B2(new_n253_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n254_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n269_), .B1(new_n283_), .B2(new_n233_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n274_), .A2(new_n278_), .A3(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n278_), .B(KEYINPUT101), .Z(new_n287_));
  AOI21_X1  g086(.A(new_n253_), .B1(new_n234_), .B2(new_n254_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n260_), .A2(new_n262_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n253_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT20), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n273_), .B1(new_n288_), .B2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n255_), .A2(new_n270_), .A3(new_n279_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n287_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n286_), .B(KEYINPUT27), .C1(new_n294_), .C2(KEYINPUT102), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n294_), .A2(KEYINPUT102), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n202_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n294_), .A2(KEYINPUT102), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(KEYINPUT102), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT27), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n271_), .A2(new_n273_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n300_), .B1(new_n301_), .B2(new_n278_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n298_), .A2(KEYINPUT103), .A3(new_n299_), .A4(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT99), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n286_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n301_), .A2(KEYINPUT99), .A3(new_n278_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n305_), .B(new_n306_), .C1(new_n278_), .C2(new_n301_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n297_), .A2(new_n303_), .B1(new_n300_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  OR3_X1    g108(.A1(new_n309_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n310_));
  INV_X1    g109(.A(G141gat), .ZN(new_n311_));
  INV_X1    g110(.A(G148gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n309_), .A2(KEYINPUT1), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(G155gat), .A3(G162gat), .ZN(new_n317_));
  OR2_X1    g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n315_), .A2(new_n317_), .A3(new_n318_), .A4(KEYINPUT89), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G141gat), .A2(G148gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT88), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT88), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(G141gat), .A3(G148gat), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n314_), .A2(KEYINPUT90), .A3(new_n319_), .A4(new_n324_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n319_), .A2(new_n324_), .A3(new_n310_), .A4(new_n313_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT90), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n320_), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n329_), .A2(KEYINPUT2), .B1(new_n313_), .B2(KEYINPUT3), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n321_), .A2(new_n323_), .ZN(new_n331_));
  OAI221_X1 g130(.A(new_n330_), .B1(KEYINPUT3), .B2(new_n313_), .C1(KEYINPUT2), .C2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n318_), .A2(new_n309_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT91), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n325_), .A2(new_n328_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G127gat), .B(G134gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G113gat), .B(G120gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT87), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n340_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n339_), .B(KEYINPUT4), .C1(new_n335_), .C2(new_n343_), .ZN(new_n344_));
  OR3_X1    g143(.A1(new_n343_), .A2(new_n335_), .A3(KEYINPUT4), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n344_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n343_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n332_), .A2(new_n334_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n326_), .A2(new_n327_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n326_), .A2(new_n327_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(new_n339_), .A3(new_n346_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n348_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G1gat), .B(G29gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G85gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT0), .B(G57gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n348_), .B2(new_n355_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT30), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n283_), .B2(new_n233_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n234_), .A2(KEYINPUT30), .A3(new_n254_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT86), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G71gat), .B(G99gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(G43gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G15gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n372_), .B(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n370_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n367_), .A2(new_n368_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT86), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n343_), .A2(KEYINPUT31), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT31), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n383_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n378_), .A2(KEYINPUT86), .A3(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n377_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  AOI211_X1 g186(.A(new_n369_), .B(new_n383_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n385_), .B1(new_n378_), .B2(KEYINPUT86), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n376_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G22gat), .B(G50gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n350_), .B(new_n394_), .C1(new_n351_), .C2(new_n352_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT92), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT92), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n335_), .A2(new_n397_), .A3(new_n394_), .ZN(new_n398_));
  XOR2_X1   g197(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n396_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n393_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n396_), .A2(new_n398_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n399_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n396_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n392_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n403_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT94), .B1(new_n267_), .B2(new_n268_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(G106gat), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G106gat), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n413_), .B(new_n410_), .C1(new_n253_), .C2(KEYINPUT94), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n353_), .A2(KEYINPUT29), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n269_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(G78gat), .ZN(new_n418_));
  INV_X1    g217(.A(G78gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n416_), .A2(new_n419_), .A3(new_n269_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n415_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n416_), .A2(new_n419_), .A3(new_n269_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n419_), .B1(new_n416_), .B2(new_n269_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n414_), .B(new_n412_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n408_), .A2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n407_), .A2(new_n403_), .A3(new_n421_), .A4(new_n424_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n391_), .A2(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n387_), .A2(new_n426_), .A3(new_n390_), .A4(new_n427_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n365_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n308_), .A2(new_n431_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n354_), .A2(new_n339_), .A3(new_n347_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n361_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT33), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(new_n356_), .B2(new_n361_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n348_), .A2(KEYINPUT33), .A3(new_n355_), .A4(new_n360_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT100), .ZN(new_n439_));
  OR2_X1    g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n439_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n437_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n278_), .A2(KEYINPUT32), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n301_), .A2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n292_), .A2(new_n293_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n444_), .B1(new_n445_), .B2(new_n443_), .ZN(new_n446_));
  OAI22_X1  g245(.A1(new_n307_), .A2(new_n442_), .B1(new_n364_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n391_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n448_), .A2(new_n428_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n432_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT104), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G113gat), .B(G141gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT79), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G169gat), .B(G197gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT77), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G29gat), .B(G36gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G43gat), .B(G50gat), .Z(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G43gat), .B(G50gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n459_), .A2(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G15gat), .B(G22gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G1gat), .A2(G8gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT14), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(G1gat), .A2(G8gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n467_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n466_), .A2(new_n467_), .A3(new_n470_), .A4(new_n468_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n458_), .B1(new_n465_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n462_), .A2(new_n464_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n476_), .A2(KEYINPUT77), .A3(new_n472_), .A4(new_n473_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n465_), .A2(KEYINPUT15), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT15), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n474_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G229gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT78), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n478_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n465_), .A2(new_n474_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n483_), .B1(new_n478_), .B2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n457_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n478_), .A2(new_n487_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n485_), .B(new_n456_), .C1(new_n490_), .C2(new_n483_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n451_), .A2(new_n452_), .A3(new_n493_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n308_), .A2(new_n431_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT104), .B1(new_n495_), .B2(new_n492_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G232gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT34), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT35), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n501_), .A2(KEYINPUT73), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT7), .ZN(new_n503_));
  INV_X1    g302(.A(G99gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n504_), .A3(new_n413_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n505_), .A2(new_n508_), .A3(new_n509_), .A4(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(G85gat), .ZN(new_n512_));
  INV_X1    g311(.A(G92gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G85gat), .A2(G92gat), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n514_), .A2(KEYINPUT67), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT8), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT8), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n511_), .A2(new_n516_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT10), .B(G99gat), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n508_), .B(new_n509_), .C1(new_n522_), .C2(G106gat), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT66), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT9), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n515_), .A2(new_n525_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n524_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n515_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(G85gat), .A2(G92gat), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT9), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(KEYINPUT66), .A3(new_n527_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n523_), .B1(new_n529_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT70), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  AOI211_X1 g335(.A(KEYINPUT70), .B(new_n523_), .C1(new_n533_), .C2(new_n529_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n521_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n479_), .A2(new_n481_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n499_), .A2(KEYINPUT35), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n529_), .A2(new_n533_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n523_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n542_), .A2(new_n543_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n541_), .B1(new_n544_), .B2(new_n476_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n502_), .B1(new_n540_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT73), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n546_), .B1(new_n547_), .B2(new_n500_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G190gat), .B(G218gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n551_), .A2(KEYINPUT36), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n540_), .A2(new_n545_), .A3(KEYINPUT73), .A4(new_n501_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(KEYINPUT36), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n548_), .A2(new_n553_), .A3(new_n554_), .A4(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT74), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n548_), .A2(new_n554_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n557_), .B1(new_n558_), .B2(new_n552_), .ZN(new_n559_));
  AOI211_X1 g358(.A(KEYINPUT74), .B(new_n553_), .C1(new_n548_), .C2(new_n554_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n556_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT37), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(G127gat), .B(G155gat), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT16), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G183gat), .B(G211gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT17), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n474_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(G64gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(G57gat), .ZN(new_n572_));
  INV_X1    g371(.A(G57gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(G64gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT11), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT69), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT69), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n572_), .A2(new_n574_), .A3(new_n578_), .A4(KEYINPUT11), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(new_n576_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT68), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(G71gat), .ZN(new_n583_));
  INV_X1    g382(.A(G71gat), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT68), .ZN(new_n585_));
  OAI21_X1  g384(.A(G78gat), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(KEYINPUT68), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n582_), .A2(G71gat), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n419_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n581_), .A2(new_n586_), .A3(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n580_), .A2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT11), .B1(new_n572_), .B2(new_n574_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n419_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n594_), .A2(new_n589_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n570_), .B(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n568_), .A2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT76), .Z(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n597_), .A2(new_n567_), .A3(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n556_), .B(KEYINPUT37), .C1(new_n559_), .C2(new_n560_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n563_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT12), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n596_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n538_), .A2(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n526_), .A2(new_n528_), .A3(new_n524_), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT66), .B1(new_n532_), .B2(new_n527_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n543_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n580_), .A2(new_n590_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n594_), .A2(new_n577_), .A3(new_n579_), .A4(new_n589_), .ZN(new_n612_));
  AND4_X1   g411(.A1(new_n521_), .A2(new_n610_), .A3(new_n611_), .A4(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n613_), .A2(new_n617_), .ZN(new_n618_));
  AOI22_X1  g417(.A1(new_n521_), .A2(new_n610_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT71), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n619_), .A2(new_n620_), .A3(KEYINPUT12), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n511_), .A2(new_n516_), .A3(new_n519_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n519_), .B1(new_n511_), .B2(new_n516_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OAI22_X1  g423(.A1(new_n624_), .A2(new_n534_), .B1(new_n591_), .B2(new_n595_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT71), .B1(new_n625_), .B2(new_n605_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n607_), .B(new_n618_), .C1(new_n621_), .C2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n613_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n616_), .B1(new_n628_), .B2(new_n625_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT5), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n632_), .B(new_n633_), .Z(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n627_), .A2(new_n630_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT72), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n627_), .A2(new_n630_), .A3(KEYINPUT72), .A4(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n627_), .A2(new_n630_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n634_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT13), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(KEYINPUT13), .A3(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n604_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n497_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n497_), .A2(KEYINPUT105), .A3(new_n649_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n364_), .B(KEYINPUT106), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(G1gat), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT38), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n654_), .A2(KEYINPUT38), .A3(new_n656_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n647_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n561_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n602_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n451_), .A2(new_n493_), .A3(new_n661_), .A4(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G1gat), .B1(new_n665_), .B2(new_n364_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n659_), .A2(new_n660_), .A3(new_n666_), .ZN(G1324gat));
  INV_X1    g466(.A(G8gat), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n297_), .A2(new_n303_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n307_), .A2(new_n300_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n654_), .A2(new_n668_), .A3(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G8gat), .B1(new_n665_), .B2(new_n308_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT39), .Z(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n672_), .A2(KEYINPUT40), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n677_));
  NOR4_X1   g476(.A1(new_n652_), .A2(new_n653_), .A3(G8gat), .A4(new_n308_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(new_n678_), .B2(new_n674_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(G1325gat));
  INV_X1    g479(.A(G15gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n654_), .A2(new_n681_), .A3(new_n448_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G15gat), .B1(new_n665_), .B2(new_n391_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT41), .Z(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1326gat));
  INV_X1    g484(.A(G22gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n654_), .A2(new_n686_), .A3(new_n428_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n428_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G22gat), .B1(new_n665_), .B2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT42), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(G1327gat));
  NAND2_X1  g490(.A1(new_n662_), .A2(new_n663_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(new_n661_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n365_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n563_), .A2(new_n603_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n451_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n698_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT43), .B1(new_n495_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n661_), .A2(new_n493_), .A3(new_n663_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(G29gat), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n655_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(new_n706_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n696_), .B1(new_n709_), .B2(new_n710_), .ZN(G1328gat));
  AOI21_X1  g510(.A(new_n703_), .B1(new_n699_), .B2(new_n701_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n308_), .B1(new_n712_), .B2(KEYINPUT44), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G36gat), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n308_), .A2(G36gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n695_), .A2(KEYINPUT45), .A3(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT45), .B1(new_n695_), .B2(new_n716_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n715_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT46), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(G36gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n713_), .B2(new_n710_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n695_), .A2(new_n716_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n717_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n722_), .B(KEYINPUT46), .C1(new_n725_), .C2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n723_), .A2(new_n731_), .ZN(G1329gat));
  INV_X1    g531(.A(new_n710_), .ZN(new_n733_));
  OAI211_X1 g532(.A(G43gat), .B(new_n448_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n695_), .A2(new_n448_), .ZN(new_n735_));
  OAI22_X1  g534(.A1(new_n733_), .A2(new_n734_), .B1(G43gat), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g536(.A(G50gat), .B1(new_n695_), .B2(new_n428_), .ZN(new_n738_));
  INV_X1    g537(.A(G50gat), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n707_), .A2(new_n739_), .A3(new_n688_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n740_), .B2(new_n710_), .ZN(G1331gat));
  NOR3_X1   g540(.A1(new_n495_), .A2(new_n493_), .A3(new_n661_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n664_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT108), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n742_), .A2(new_n745_), .A3(new_n664_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n573_), .B1(new_n747_), .B2(new_n365_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n604_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n742_), .A2(new_n749_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n750_), .A2(G57gat), .A3(new_n655_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1332gat));
  NAND2_X1  g551(.A1(new_n747_), .A2(new_n671_), .ZN(new_n753_));
  XOR2_X1   g552(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(G64gat), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n753_), .B2(G64gat), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n671_), .A2(new_n571_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT110), .ZN(new_n758_));
  OAI22_X1  g557(.A1(new_n755_), .A2(new_n756_), .B1(new_n750_), .B2(new_n758_), .ZN(G1333gat));
  INV_X1    g558(.A(new_n750_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(new_n584_), .A3(new_n448_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n744_), .A2(new_n448_), .A3(new_n746_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G71gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G71gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  OAI211_X1 g567(.A(KEYINPUT111), .B(new_n761_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1334gat));
  NAND2_X1  g569(.A1(new_n428_), .A2(new_n419_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT112), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n760_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n744_), .A2(new_n428_), .A3(new_n746_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(G78gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G78gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT113), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n773_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1335gat));
  NAND2_X1  g581(.A1(new_n742_), .A2(new_n693_), .ZN(new_n783_));
  OR3_X1    g582(.A1(new_n783_), .A2(G85gat), .A3(new_n655_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n661_), .A2(new_n493_), .A3(new_n602_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n702_), .A2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(new_n365_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n784_), .B1(new_n787_), .B2(new_n512_), .ZN(G1336gat));
  INV_X1    g587(.A(new_n783_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(new_n513_), .A3(new_n671_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n786_), .A2(new_n671_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n513_), .ZN(G1337gat));
  AOI21_X1  g591(.A(new_n504_), .B1(new_n786_), .B2(new_n448_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n783_), .A2(new_n391_), .A3(new_n522_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795_));
  OAI22_X1  g594(.A1(new_n793_), .A2(new_n794_), .B1(new_n795_), .B2(KEYINPUT51), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(KEYINPUT51), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n796_), .B(new_n797_), .ZN(G1338gat));
  NAND3_X1  g597(.A1(new_n789_), .A2(new_n413_), .A3(new_n428_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n697_), .B1(new_n451_), .B2(new_n698_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n495_), .A2(KEYINPUT43), .A3(new_n700_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n428_), .B(new_n785_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n702_), .A2(KEYINPUT115), .A3(new_n428_), .A4(new_n785_), .ZN(new_n806_));
  AND4_X1   g605(.A1(new_n800_), .A2(new_n805_), .A3(G106gat), .A4(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n413_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n800_), .B1(new_n808_), .B2(new_n806_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n799_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT53), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n812_), .B(new_n799_), .C1(new_n807_), .C2(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1339gat));
  INV_X1    g613(.A(G113gat), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n627_), .A2(KEYINPUT55), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n620_), .B1(new_n619_), .B2(KEYINPUT12), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n625_), .A2(KEYINPUT71), .A3(new_n605_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n818_), .A2(new_n819_), .B1(new_n538_), .B2(new_n606_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n618_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n817_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n628_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n617_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n635_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(KEYINPUT117), .A3(new_n828_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n817_), .A2(new_n822_), .B1(new_n824_), .B2(new_n617_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n827_), .B1(new_n830_), .B2(new_n635_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  INV_X1    g631(.A(new_n828_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n829_), .A2(new_n831_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n640_), .B2(new_n493_), .ZN(new_n837_));
  AOI211_X1 g636(.A(KEYINPUT116), .B(new_n492_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n816_), .B1(new_n835_), .B2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n829_), .A2(new_n831_), .A3(new_n834_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n841_), .B(KEYINPUT118), .C1(new_n837_), .C2(new_n838_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n484_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n478_), .A2(new_n482_), .A3(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n457_), .B(new_n844_), .C1(new_n490_), .C2(new_n843_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n491_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n643_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n840_), .A2(new_n842_), .A3(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n561_), .A2(KEYINPUT57), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n640_), .A2(new_n846_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT56), .B1(new_n826_), .B2(new_n634_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n830_), .A2(new_n833_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n851_), .B(KEYINPUT58), .C1(new_n852_), .C2(new_n853_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n856_), .A2(new_n698_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n850_), .A2(new_n859_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(new_n848_), .B2(new_n561_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n663_), .B1(new_n860_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n648_), .B2(new_n492_), .ZN(new_n866_));
  NOR4_X1   g665(.A1(new_n604_), .A2(new_n647_), .A3(KEYINPUT54), .A4(new_n493_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n864_), .A2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n671_), .A2(new_n655_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n430_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n870_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n815_), .B1(new_n875_), .B2(new_n492_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT120), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n878_), .B(new_n815_), .C1(new_n875_), .C2(new_n492_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n847_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n841_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n816_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n662_), .B1(new_n882_), .B2(new_n842_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n850_), .B(new_n859_), .C1(new_n883_), .C2(new_n862_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n868_), .B1(new_n884_), .B2(new_n663_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n886_));
  OAI22_X1  g685(.A1(new_n885_), .A2(new_n873_), .B1(new_n886_), .B2(KEYINPUT59), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n888_));
  NAND3_X1  g687(.A1(new_n870_), .A2(new_n874_), .A3(new_n888_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n492_), .A2(new_n815_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n877_), .A2(new_n879_), .B1(new_n890_), .B2(new_n891_), .ZN(G1340gat));
  INV_X1    g691(.A(new_n875_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT122), .B(G120gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n894_), .B1(new_n661_), .B2(KEYINPUT60), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n893_), .B(new_n895_), .C1(KEYINPUT60), .C2(new_n894_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n887_), .A2(new_n889_), .A3(new_n647_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n894_), .ZN(G1341gat));
  NAND3_X1  g697(.A1(new_n887_), .A2(new_n889_), .A3(new_n602_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G127gat), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n663_), .A2(G127gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n875_), .B2(new_n901_), .ZN(G1342gat));
  AOI21_X1  g701(.A(G134gat), .B1(new_n893_), .B2(new_n662_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n698_), .A2(G134gat), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n904_), .B(KEYINPUT123), .Z(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n890_), .B2(new_n905_), .ZN(G1343gat));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n429_), .B1(new_n864_), .B2(new_n869_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n871_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n871_), .ZN(new_n910_));
  NOR4_X1   g709(.A1(new_n885_), .A2(KEYINPUT124), .A3(new_n429_), .A4(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n493_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(G141gat), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n311_), .B(new_n493_), .C1(new_n909_), .C2(new_n911_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1344gat));
  OAI21_X1  g714(.A(new_n647_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT125), .B(G148gat), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n647_), .B(new_n917_), .C1(new_n909_), .C2(new_n911_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1345gat));
  OAI21_X1  g720(.A(new_n602_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT61), .B(G155gat), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n923_), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n602_), .B(new_n925_), .C1(new_n909_), .C2(new_n911_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1346gat));
  INV_X1    g726(.A(G162gat), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n928_), .B(new_n662_), .C1(new_n909_), .C2(new_n911_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n908_), .A2(new_n871_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(KEYINPUT124), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n908_), .A2(new_n907_), .A3(new_n871_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n700_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n929_), .B1(new_n933_), .B2(new_n928_), .ZN(G1347gat));
  AND3_X1   g733(.A1(new_n671_), .A2(new_n655_), .A3(new_n872_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n848_), .A2(new_n561_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n861_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n858_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n602_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n493_), .B(new_n935_), .C1(new_n939_), .C2(new_n868_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n870_), .A2(KEYINPUT126), .A3(new_n493_), .A4(new_n935_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n942_), .A2(G169gat), .A3(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n942_), .A2(new_n943_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n870_), .A2(new_n935_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n949_), .A2(new_n258_), .A3(new_n493_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n946_), .A2(new_n947_), .A3(new_n950_), .ZN(G1348gat));
  NOR2_X1   g750(.A1(new_n948_), .A2(new_n661_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(new_n206_), .ZN(G1349gat));
  NOR2_X1   g752(.A1(new_n948_), .A2(new_n663_), .ZN(new_n954_));
  MUX2_X1   g753(.A(G183gat), .B(new_n218_), .S(new_n954_), .Z(G1350gat));
  OAI21_X1  g754(.A(G190gat), .B1(new_n948_), .B2(new_n700_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n662_), .A2(new_n221_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n948_), .B2(new_n957_), .ZN(G1351gat));
  AOI22_X1  g757(.A1(new_n387_), .A2(new_n390_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n308_), .A2(new_n365_), .ZN(new_n960_));
  OAI211_X1 g759(.A(new_n959_), .B(new_n960_), .C1(new_n939_), .C2(new_n868_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n961_), .A2(new_n492_), .ZN(new_n962_));
  XOR2_X1   g761(.A(new_n962_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g762(.A1(new_n961_), .A2(new_n661_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n964_), .A2(G204gat), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n965_), .B1(new_n239_), .B2(new_n964_), .ZN(G1353gat));
  NOR2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  AND2_X1   g766(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n968_));
  NOR4_X1   g767(.A1(new_n961_), .A2(new_n663_), .A3(new_n967_), .A4(new_n968_), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n908_), .A2(new_n602_), .A3(new_n960_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n969_), .B1(new_n970_), .B2(new_n967_), .ZN(G1354gat));
  OAI21_X1  g770(.A(G218gat), .B1(new_n961_), .B2(new_n700_), .ZN(new_n972_));
  INV_X1    g771(.A(G218gat), .ZN(new_n973_));
  NAND4_X1  g772(.A1(new_n908_), .A2(new_n973_), .A3(new_n662_), .A4(new_n960_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n972_), .A2(new_n974_), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n975_), .A2(new_n976_), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n972_), .A2(KEYINPUT127), .A3(new_n974_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n977_), .A2(new_n978_), .ZN(G1355gat));
endmodule


