//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT81), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT24), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  OAI211_X1 g005(.A(new_n203_), .B(KEYINPUT24), .C1(new_n205_), .C2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT23), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n204_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT80), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n209_), .B1(G183gat), .B2(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT82), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(G169gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n210_), .A2(new_n214_), .B1(new_n217_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G227gat), .A2(G233gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT83), .ZN(new_n224_));
  XOR2_X1   g023(.A(new_n224_), .B(KEYINPUT30), .Z(new_n225_));
  XNOR2_X1  g024(.A(new_n222_), .B(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G71gat), .B(G99gat), .Z(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G127gat), .B(G134gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT84), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G113gat), .B(G120gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT31), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G15gat), .B(G43gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n228_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n228_), .A2(new_n235_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G211gat), .B(G218gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G197gat), .B(G204gat), .Z(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(KEYINPUT21), .A3(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT90), .ZN(new_n243_));
  OR3_X1    g042(.A1(new_n241_), .A2(KEYINPUT89), .A3(KEYINPUT21), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT21), .B1(new_n241_), .B2(KEYINPUT89), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n239_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT20), .B1(new_n222_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G226gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT19), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT24), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n211_), .A2(new_n212_), .B1(new_n253_), .B2(new_n202_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n207_), .A2(new_n254_), .A3(new_n209_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT96), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n207_), .A2(new_n254_), .A3(KEYINPUT96), .A4(new_n209_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n215_), .A2(new_n219_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n259_), .A2(KEYINPUT97), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(KEYINPUT97), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n257_), .B(new_n258_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(new_n247_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n263_), .A2(KEYINPUT99), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT99), .ZN(new_n265_));
  NOR3_X1   g064(.A1(new_n262_), .A2(new_n265_), .A3(new_n247_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n252_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n251_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT20), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n269_), .B1(new_n222_), .B2(new_n248_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n262_), .A2(new_n247_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n268_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT98), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  AOI211_X1 g073(.A(KEYINPUT98), .B(new_n268_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n267_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G8gat), .B(G36gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT18), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G64gat), .B(G92gat), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n278_), .B(new_n279_), .Z(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(new_n281_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n267_), .B(new_n280_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT27), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT27), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n248_), .A2(new_n259_), .A3(new_n255_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n251_), .B1(new_n286_), .B2(new_n249_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n270_), .A2(new_n271_), .A3(new_n268_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n285_), .B1(new_n289_), .B2(new_n281_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n283_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n284_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n232_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G141gat), .B(G148gat), .ZN(new_n295_));
  INV_X1    g094(.A(G155gat), .ZN(new_n296_));
  INV_X1    g095(.A(G162gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(KEYINPUT85), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT85), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(G155gat), .B2(G162gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  AOI22_X1  g100(.A1(new_n298_), .A2(new_n300_), .B1(KEYINPUT1), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT86), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n301_), .A2(KEYINPUT1), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n305_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n295_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n301_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n298_), .A2(new_n300_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT87), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NOR3_X1   g112(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  AOI211_X1 g115(.A(new_n308_), .B(new_n309_), .C1(new_n311_), .C2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n294_), .B1(new_n307_), .B2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n307_), .A2(new_n317_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n232_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n318_), .A2(KEYINPUT4), .A3(new_n320_), .ZN(new_n326_));
  OR3_X1    g125(.A1(new_n319_), .A2(new_n232_), .A3(KEYINPUT4), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n322_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G1gat), .B(G29gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(G85gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT0), .B(G57gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n325_), .A2(new_n329_), .A3(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n333_), .B1(new_n324_), .B2(new_n328_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT93), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT29), .B1(new_n307_), .B2(new_n317_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n247_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G228gat), .A2(G233gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n342_), .A3(new_n247_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G78gat), .B(G106gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n347_), .B(KEYINPUT91), .Z(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n339_), .B1(new_n346_), .B2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n344_), .A2(KEYINPUT93), .A3(new_n348_), .A4(new_n345_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n319_), .A2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NOR4_X1   g156(.A1(new_n307_), .A2(new_n317_), .A3(KEYINPUT29), .A4(new_n356_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G22gat), .B(G50gat), .Z(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n360_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n356_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(new_n319_), .B2(new_n354_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n364_), .B2(new_n358_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n350_), .A2(new_n352_), .A3(new_n353_), .A4(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT94), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n351_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n370_), .A2(KEYINPUT94), .A3(new_n353_), .A4(new_n350_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT92), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n346_), .A2(new_n349_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n374_), .A2(new_n351_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n373_), .B1(new_n375_), .B2(new_n366_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n366_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n377_), .B(KEYINPUT92), .C1(new_n374_), .C2(new_n351_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n372_), .A2(new_n379_), .A3(KEYINPUT95), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT95), .B1(new_n372_), .B2(new_n379_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n293_), .B(new_n338_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n280_), .A2(KEYINPUT32), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n289_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n337_), .B(new_n386_), .C1(new_n276_), .C2(new_n385_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT33), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n336_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n321_), .A2(new_n323_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n326_), .A2(new_n322_), .A3(new_n327_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n334_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n282_), .A2(new_n389_), .A3(new_n283_), .A4(new_n392_), .ZN(new_n393_));
  OAI211_X1 g192(.A(KEYINPUT33), .B(new_n333_), .C1(new_n324_), .C2(new_n328_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT100), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n387_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n382_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n380_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n238_), .B1(new_n383_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n380_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n293_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n238_), .A2(new_n338_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n399_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT68), .ZN(new_n405_));
  AND2_X1   g204(.A1(G85gat), .A2(G92gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G85gat), .A2(G92gat), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT8), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT67), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n411_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  OR3_X1    g214(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(KEYINPUT67), .A3(new_n412_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G99gat), .A2(G106gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT6), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(G99gat), .A3(G106gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT66), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n420_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n423_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n410_), .B1(new_n418_), .B2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n413_), .A2(new_n414_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n420_), .A2(new_n422_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n408_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(G85gat), .B2(G92gat), .ZN(new_n432_));
  AND2_X1   g231(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(G85gat), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n436_));
  NOR2_X1   g235(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n432_), .B1(new_n435_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT10), .B(G99gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n429_), .B1(new_n440_), .B2(G106gat), .ZN(new_n441_));
  OAI22_X1  g240(.A1(new_n430_), .A2(KEYINPUT8), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n405_), .B1(new_n427_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n429_), .A2(KEYINPUT66), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n420_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n444_), .A2(new_n415_), .A3(new_n417_), .A4(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT8), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n408_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n429_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n416_), .A2(new_n412_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n409_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n447_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n439_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n441_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n449_), .A2(new_n453_), .A3(new_n456_), .A4(KEYINPUT68), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n443_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT11), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G71gat), .B(G78gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G57gat), .B(G64gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT69), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(G57gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n465_), .A2(G64gat), .ZN(new_n466_));
  INV_X1    g265(.A(G64gat), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n467_), .A2(G57gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT69), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  AOI211_X1 g268(.A(new_n459_), .B(new_n461_), .C1(new_n464_), .C2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n464_), .A2(new_n469_), .A3(new_n459_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n464_), .A2(new_n469_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n460_), .B1(new_n472_), .B2(KEYINPUT11), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n470_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT12), .B1(new_n458_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(KEYINPUT11), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(new_n461_), .A3(new_n471_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n472_), .A2(KEYINPUT11), .A3(new_n460_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n443_), .A2(new_n479_), .A3(new_n457_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n449_), .A2(new_n456_), .A3(new_n453_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n474_), .A2(KEYINPUT12), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n475_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G230gat), .A2(G233gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n458_), .A2(new_n474_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n487_), .A2(new_n480_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n486_), .B1(new_n488_), .B2(new_n485_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G120gat), .B(G148gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT5), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G176gat), .B(G204gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n493_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n486_), .B(new_n495_), .C1(new_n488_), .C2(new_n485_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT13), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n494_), .A2(KEYINPUT13), .A3(new_n496_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT79), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G113gat), .B(G141gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G169gat), .B(G197gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(new_n504_), .Z(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G29gat), .B(G36gat), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n507_), .A2(KEYINPUT70), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(KEYINPUT70), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n508_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518_));
  INV_X1    g317(.A(G1gat), .ZN(new_n519_));
  INV_X1    g318(.A(G8gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT14), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G1gat), .B(G8gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  NOR3_X1   g323(.A1(new_n516_), .A2(new_n517_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n524_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n513_), .A2(new_n514_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n525_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n528_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n526_), .A2(new_n527_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n529_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n506_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n531_), .A2(new_n534_), .A3(new_n506_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n502_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n537_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n539_), .A2(KEYINPUT79), .A3(new_n535_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n501_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n404_), .A2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT72), .B1(new_n458_), .B2(new_n527_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT34), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n547_), .A2(KEYINPUT35), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n516_), .A2(new_n517_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n549_), .B2(new_n481_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n527_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT72), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n443_), .A2(new_n551_), .A3(new_n552_), .A4(new_n457_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n545_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(KEYINPUT35), .A3(new_n547_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT73), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G134gat), .B(G162gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(KEYINPUT36), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n547_), .A2(KEYINPUT35), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n550_), .A2(new_n545_), .A3(new_n562_), .A4(new_n553_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n555_), .A2(new_n561_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT74), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT74), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n555_), .A2(new_n566_), .A3(new_n561_), .A4(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n555_), .A2(new_n563_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n559_), .B(KEYINPUT36), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n568_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(G231gat), .ZN(new_n578_));
  INV_X1    g377(.A(G233gat), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n479_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n477_), .A2(new_n478_), .B1(G231gat), .B2(G233gat), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT76), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n580_), .A2(new_n581_), .A3(KEYINPUT76), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n583_), .A2(new_n526_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n584_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n524_), .B1(new_n586_), .B2(new_n582_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT77), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G127gat), .B(G155gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT16), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G183gat), .B(G211gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n526_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n586_), .A2(new_n524_), .A3(new_n582_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT77), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n588_), .A2(new_n594_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT78), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n595_), .A2(new_n596_), .A3(KEYINPUT78), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n592_), .B(KEYINPUT17), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n577_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n544_), .A2(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n607_), .A2(G1gat), .A3(new_n338_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n608_), .A2(KEYINPUT38), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(KEYINPUT38), .ZN(new_n610_));
  INV_X1    g409(.A(new_n572_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n404_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT101), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n543_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n501_), .A2(KEYINPUT101), .A3(new_n542_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n605_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n612_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n617_), .B2(new_n338_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n609_), .A2(new_n610_), .A3(new_n618_), .ZN(G1324gat));
  OAI21_X1  g418(.A(G8gat), .B1(new_n617_), .B2(new_n293_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT39), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n401_), .A2(new_n520_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n607_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(G1325gat));
  INV_X1    g424(.A(new_n238_), .ZN(new_n626_));
  OR3_X1    g425(.A1(new_n607_), .A2(G15gat), .A3(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n612_), .A2(new_n238_), .A3(new_n616_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT41), .B1(new_n628_), .B2(G15gat), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT102), .Z(G1326gat));
  INV_X1    g432(.A(new_n400_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G22gat), .B1(new_n617_), .B2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT42), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n634_), .A2(G22gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n636_), .B1(new_n607_), .B2(new_n637_), .ZN(G1327gat));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n614_), .A2(new_n615_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n640_), .B2(new_n605_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n605_), .ZN(new_n642_));
  AOI211_X1 g441(.A(KEYINPUT103), .B(new_n642_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n577_), .B1(new_n399_), .B2(new_n403_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n645_), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT43), .B1(new_n645_), .B2(KEYINPUT104), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n644_), .B(KEYINPUT44), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(G29gat), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n338_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n641_), .A2(new_n643_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n645_), .A2(KEYINPUT104), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n645_), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n651_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n657_));
  OAI211_X1 g456(.A(new_n648_), .B(new_n650_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n383_), .A2(new_n398_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n626_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n403_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT106), .ZN(new_n663_));
  INV_X1    g462(.A(new_n543_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n642_), .A2(new_n572_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n662_), .A2(new_n663_), .A3(new_n664_), .A4(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n664_), .B(new_n665_), .C1(new_n399_), .C2(new_n403_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT106), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n649_), .B1(new_n669_), .B2(new_n338_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n658_), .A2(new_n670_), .ZN(G1328gat));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT108), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT109), .Z(new_n674_));
  OAI211_X1 g473(.A(new_n648_), .B(new_n401_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G36gat), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n293_), .A2(KEYINPUT107), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n293_), .A2(KEYINPUT107), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(G36gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n666_), .A2(new_n668_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT45), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n666_), .A2(new_n668_), .A3(KEYINPUT45), .A4(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n676_), .A2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n672_), .A2(KEYINPUT108), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n674_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n686_), .B1(new_n675_), .B2(G36gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n674_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n692_), .A2(new_n689_), .A3(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1329gat));
  INV_X1    g494(.A(G43gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n696_), .B1(new_n669_), .B2(new_n626_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT110), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n626_), .A2(new_n696_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n648_), .B(new_n699_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n698_), .A2(KEYINPUT47), .A3(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT47), .B1(new_n698_), .B2(new_n701_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1330gat));
  OR3_X1    g503(.A1(new_n669_), .A2(G50gat), .A3(new_n634_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n648_), .B(new_n400_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(G50gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n706_), .B2(G50gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1331gat));
  NOR2_X1   g509(.A1(new_n404_), .A2(new_n542_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n577_), .A2(new_n605_), .A3(new_n501_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n465_), .B1(new_n713_), .B2(new_n338_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n501_), .A2(new_n605_), .A3(new_n542_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n612_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n338_), .B2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n717_), .B2(G57gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n714_), .B1(new_n716_), .B2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT113), .ZN(G1332gat));
  NAND3_X1  g520(.A1(new_n612_), .A2(new_n679_), .A3(new_n715_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n723_), .A3(G64gat), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n723_), .B1(new_n722_), .B2(G64gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n679_), .A2(new_n467_), .ZN(new_n727_));
  OAI22_X1  g526(.A1(new_n725_), .A2(new_n726_), .B1(new_n713_), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT114), .ZN(G1333gat));
  OAI21_X1  g528(.A(G71gat), .B1(new_n716_), .B2(new_n626_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT49), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n626_), .A2(G71gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n713_), .B2(new_n732_), .ZN(G1334gat));
  OAI21_X1  g532(.A(G78gat), .B1(new_n716_), .B2(new_n634_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT50), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n634_), .A2(G78gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n713_), .B2(new_n736_), .ZN(G1335gat));
  INV_X1    g536(.A(G85gat), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n501_), .A2(new_n642_), .A3(new_n572_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n711_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n738_), .B1(new_n740_), .B2(new_n338_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT115), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n654_), .A2(new_n655_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n501_), .A2(new_n642_), .A3(new_n542_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n338_), .A2(new_n738_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(G1336gat));
  INV_X1    g546(.A(new_n740_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G92gat), .B1(new_n748_), .B2(new_n401_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n433_), .A2(new_n434_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n680_), .A2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n745_), .B2(new_n751_), .ZN(G1337gat));
  NOR2_X1   g551(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n743_), .A2(new_n238_), .A3(new_n744_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G99gat), .ZN(new_n755_));
  OR3_X1    g554(.A1(new_n740_), .A2(new_n440_), .A3(new_n626_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n753_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n757_), .B(new_n758_), .Z(G1338gat));
  OR3_X1    g558(.A1(new_n740_), .A2(G106gat), .A3(new_n634_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n400_), .B(new_n744_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(new_n762_), .A3(G106gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(G106gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g565(.A(new_n577_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n599_), .A2(new_n604_), .A3(new_n541_), .ZN(new_n769_));
  AND4_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(new_n499_), .A4(new_n500_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n768_), .B1(new_n501_), .B2(new_n769_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT54), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n767_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT121), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n611_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT56), .ZN(new_n780_));
  INV_X1    g579(.A(new_n485_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n475_), .B2(new_n483_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT118), .B(new_n781_), .C1(new_n475_), .C2(new_n483_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n479_), .B1(new_n443_), .B2(new_n457_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n480_), .B(new_n482_), .C1(new_n786_), .C2(KEYINPUT12), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT55), .B1(new_n787_), .B2(new_n781_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT12), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n487_), .A2(new_n789_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n480_), .A2(new_n482_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n790_), .A2(new_n791_), .A3(new_n792_), .A4(new_n485_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n784_), .A2(new_n785_), .B1(new_n788_), .B2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n780_), .B1(new_n794_), .B2(new_n495_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n495_), .A2(new_n780_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT119), .B1(new_n794_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n792_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n787_), .A2(KEYINPUT55), .A3(new_n781_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n785_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT118), .B1(new_n787_), .B2(new_n781_), .ZN(new_n802_));
  OAI22_X1  g601(.A1(new_n799_), .A2(new_n800_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n804_), .A3(new_n796_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n795_), .A2(new_n798_), .A3(new_n805_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n538_), .A2(new_n540_), .A3(new_n496_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OR3_X1    g607(.A1(new_n525_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n532_), .A2(new_n533_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n505_), .B1(new_n810_), .B2(new_n529_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  AOI211_X1 g611(.A(new_n537_), .B(new_n812_), .C1(new_n494_), .C2(new_n496_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n777_), .B(new_n779_), .C1(new_n808_), .C2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n496_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n815_), .A2(new_n537_), .A3(new_n812_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n795_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n794_), .A2(new_n797_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n816_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT58), .B(new_n816_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n577_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n813_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n572_), .A2(KEYINPUT57), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT121), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n778_), .B1(new_n824_), .B2(new_n611_), .ZN(new_n827_));
  AND4_X1   g626(.A1(new_n814_), .A2(new_n823_), .A3(new_n826_), .A4(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n776_), .B1(new_n642_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830_));
  NOR4_X1   g629(.A1(new_n400_), .A2(new_n401_), .A3(new_n338_), .A4(new_n626_), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n827_), .A2(KEYINPUT120), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n778_), .C1(new_n824_), .C2(new_n611_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n814_), .A2(new_n823_), .A3(new_n826_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n605_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n776_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT122), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n838_), .A2(new_n841_), .A3(new_n776_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n831_), .ZN(new_n844_));
  AOI211_X1 g643(.A(new_n541_), .B(new_n832_), .C1(new_n844_), .C2(KEYINPUT59), .ZN(new_n845_));
  INV_X1    g644(.A(G113gat), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n542_), .A2(new_n846_), .ZN(new_n847_));
  OAI22_X1  g646(.A1(new_n845_), .A2(new_n846_), .B1(new_n844_), .B2(new_n847_), .ZN(G1340gat));
  INV_X1    g647(.A(new_n844_), .ZN(new_n849_));
  INV_X1    g648(.A(G120gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n501_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n849_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n850_), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n501_), .B(new_n832_), .C1(new_n844_), .C2(KEYINPUT59), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n850_), .ZN(G1341gat));
  INV_X1    g653(.A(G127gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n849_), .A2(new_n855_), .A3(new_n642_), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n605_), .B(new_n832_), .C1(new_n844_), .C2(KEYINPUT59), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n855_), .ZN(G1342gat));
  INV_X1    g657(.A(G134gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n849_), .A2(new_n859_), .A3(new_n611_), .ZN(new_n860_));
  AOI211_X1 g659(.A(new_n767_), .B(new_n832_), .C1(new_n844_), .C2(KEYINPUT59), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n859_), .ZN(G1343gat));
  NOR4_X1   g661(.A1(new_n679_), .A2(new_n634_), .A3(new_n338_), .A4(new_n238_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n843_), .A2(new_n542_), .A3(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g664(.A(new_n501_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n843_), .A2(new_n866_), .A3(new_n863_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g667(.A1(new_n843_), .A2(new_n642_), .A3(new_n863_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT61), .B(G155gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1346gat));
  NAND4_X1  g670(.A1(new_n843_), .A2(G162gat), .A3(new_n577_), .A4(new_n863_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n840_), .A2(new_n611_), .A3(new_n842_), .A4(new_n863_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n873_), .A2(KEYINPUT123), .A3(new_n297_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT123), .B1(new_n873_), .B2(new_n297_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n872_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  OAI211_X1 g677(.A(KEYINPUT124), .B(new_n872_), .C1(new_n874_), .C2(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1347gat));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n829_), .A2(new_n634_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n402_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n679_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n542_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  AND4_X1   g686(.A1(new_n881_), .A2(new_n886_), .A3(new_n887_), .A4(G169gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n205_), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n886_), .A2(new_n889_), .B1(new_n881_), .B2(new_n887_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT22), .B(G169gat), .Z(new_n891_));
  OAI22_X1  g690(.A1(new_n888_), .A2(new_n890_), .B1(new_n886_), .B2(new_n891_), .ZN(G1348gat));
  INV_X1    g691(.A(new_n882_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n884_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n206_), .B1(new_n895_), .B2(new_n501_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n897_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n843_), .A2(new_n634_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n894_), .A2(G176gat), .A3(new_n866_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  AOI22_X1  g701(.A1(new_n898_), .A2(new_n899_), .B1(new_n900_), .B2(new_n902_), .ZN(G1349gat));
  NOR2_X1   g702(.A1(new_n884_), .A2(new_n605_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n840_), .A2(new_n634_), .A3(new_n842_), .A4(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(G183gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n211_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n893_), .A2(new_n908_), .A3(new_n904_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT127), .Z(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n895_), .B2(new_n767_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n885_), .A2(new_n611_), .A3(new_n212_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1351gat));
  NOR4_X1   g713(.A1(new_n680_), .A2(new_n634_), .A3(new_n337_), .A4(new_n238_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n843_), .A2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n542_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n866_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g719(.A(KEYINPUT63), .B(G211gat), .C1(new_n916_), .C2(new_n642_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT63), .B(G211gat), .Z(new_n922_));
  AND3_X1   g721(.A1(new_n916_), .A2(new_n642_), .A3(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1354gat));
  NAND2_X1  g723(.A1(new_n843_), .A2(new_n915_), .ZN(new_n925_));
  OAI21_X1  g724(.A(G218gat), .B1(new_n925_), .B2(new_n767_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n572_), .A2(G218gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n925_), .B2(new_n927_), .ZN(G1355gat));
endmodule


