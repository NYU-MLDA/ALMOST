//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_;
  INV_X1    g000(.A(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  OR2_X1    g003(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n204_), .B1(new_n207_), .B2(new_n203_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n211_), .B(new_n212_), .C1(G183gat), .C2(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n211_), .A2(new_n212_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n216_), .A2(KEYINPUT78), .ZN(new_n217_));
  INV_X1    g016(.A(new_n204_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(KEYINPUT78), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT24), .A4(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n217_), .A2(new_n219_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n215_), .B(new_n220_), .C1(new_n221_), .C2(KEYINPUT24), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT77), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(G190gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT26), .ZN(new_n225_));
  INV_X1    g024(.A(G183gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT25), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G183gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT76), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n227_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n226_), .A2(KEYINPUT25), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(KEYINPUT76), .ZN(new_n233_));
  NOR3_X1   g032(.A1(new_n225_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n214_), .B1(new_n222_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT30), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n236_), .A2(KEYINPUT80), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G227gat), .A2(G233gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT79), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(G15gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G71gat), .B(G99gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(G43gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n240_), .B(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G113gat), .B(G120gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  NAND2_X1  g048(.A1(new_n236_), .A2(KEYINPUT80), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n237_), .A2(new_n250_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n244_), .B(new_n249_), .C1(new_n251_), .C2(new_n243_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n249_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n244_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n243_), .B1(new_n237_), .B2(new_n250_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT27), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G197gat), .A2(G204gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT85), .B(G197gat), .ZN(new_n260_));
  OAI211_X1 g059(.A(KEYINPUT21), .B(new_n259_), .C1(new_n260_), .C2(G204gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(G211gat), .B(G218gat), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(G204gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(G197gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(new_n260_), .B2(new_n264_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n261_), .B(new_n263_), .C1(new_n266_), .C2(KEYINPUT21), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(KEYINPUT21), .A3(new_n262_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n235_), .A2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(KEYINPUT26), .B(G190gat), .Z(new_n271_));
  NAND2_X1  g070(.A1(new_n229_), .A2(new_n227_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n272_), .A2(KEYINPUT89), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(KEYINPUT89), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n271_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n222_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n207_), .A2(new_n203_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT90), .B1(new_n277_), .B2(new_n218_), .ZN(new_n278_));
  AOI21_X1  g077(.A(G176gat), .B1(new_n205_), .B2(new_n206_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT90), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n204_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n213_), .B(KEYINPUT91), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT92), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n208_), .A2(KEYINPUT90), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n280_), .B1(new_n279_), .B2(new_n204_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT91), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n213_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT92), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n276_), .B1(new_n284_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n269_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n270_), .B(KEYINPUT20), .C1(new_n292_), .C2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G226gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(G64gat), .B(G92gat), .Z(new_n299_));
  XNOR2_X1  g098(.A(G8gat), .B(G36gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  AOI21_X1  g102(.A(new_n297_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT20), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n305_), .B1(new_n235_), .B2(new_n269_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n298_), .A2(new_n303_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n303_), .B1(new_n298_), .B2(new_n307_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n258_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n294_), .A2(new_n297_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n303_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n303_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n294_), .A2(new_n297_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n297_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n276_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n287_), .A2(new_n289_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n269_), .A2(KEYINPUT86), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT86), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n316_), .B(new_n317_), .C1(new_n318_), .C2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n315_), .B1(new_n321_), .B2(new_n306_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n313_), .B1(new_n314_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n312_), .A2(new_n323_), .A3(KEYINPUT27), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n310_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(KEYINPUT83), .A2(G233gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(KEYINPUT83), .A2(G233gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(G228gat), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT84), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n331_));
  INV_X1    g130(.A(G141gat), .ZN(new_n332_));
  INV_X1    g131(.A(G148gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n334_), .A2(new_n336_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340_));
  OR2_X1    g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(KEYINPUT1), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(G155gat), .A3(G162gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n345_), .A3(new_n341_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G141gat), .B(G148gat), .Z(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n342_), .A2(new_n348_), .A3(KEYINPUT82), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT82), .B1(new_n342_), .B2(new_n348_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT29), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n269_), .B(new_n330_), .C1(new_n351_), .C2(new_n352_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n342_), .A2(new_n348_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(new_n352_), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n318_), .A2(new_n355_), .A3(new_n320_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n353_), .B1(new_n356_), .B2(new_n329_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n351_), .A2(new_n352_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT28), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  NOR4_X1   g161(.A1(new_n349_), .A2(new_n350_), .A3(KEYINPUT29), .A4(new_n361_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G78gat), .B(G106gat), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT87), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n362_), .A2(new_n364_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n360_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n366_), .B1(new_n369_), .B2(new_n363_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n357_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n357_), .B1(new_n370_), .B2(new_n368_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(KEYINPUT95), .B(KEYINPUT0), .Z(new_n374_));
  XNOR2_X1  g173(.A(G1gat), .B(G29gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G57gat), .B(G85gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT94), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381_));
  INV_X1    g180(.A(new_n247_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n381_), .B(new_n382_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n382_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n354_), .A2(new_n247_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n380_), .B(new_n383_), .C1(new_n386_), .C2(new_n381_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n384_), .A2(KEYINPUT94), .A3(KEYINPUT4), .A4(new_n385_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n379_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n379_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n386_), .A2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n378_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n384_), .A2(KEYINPUT4), .A3(new_n385_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n383_), .A2(new_n380_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n388_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n391_), .B1(new_n395_), .B2(new_n390_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n378_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n373_), .A2(new_n392_), .A3(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT97), .B1(new_n325_), .B2(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n373_), .A2(new_n392_), .A3(new_n398_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT97), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n401_), .A2(new_n402_), .A3(new_n310_), .A4(new_n324_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n398_), .A2(KEYINPUT33), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n396_), .A2(new_n406_), .A3(new_n397_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n395_), .A2(new_n379_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n409_), .B(new_n378_), .C1(new_n379_), .C2(new_n386_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n298_), .A2(new_n307_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n313_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n410_), .A2(new_n412_), .A3(new_n312_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n408_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n303_), .A2(KEYINPUT32), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT96), .B1(new_n311_), .B2(new_n415_), .ZN(new_n416_));
  AND4_X1   g215(.A1(KEYINPUT96), .A2(new_n298_), .A3(new_n307_), .A4(new_n415_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n282_), .A2(new_n283_), .A3(KEYINPUT92), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n290_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n316_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n305_), .B1(new_n421_), .B2(new_n269_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n315_), .A3(new_n270_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n322_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n415_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n398_), .B2(new_n392_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n418_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n373_), .B1(new_n414_), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n257_), .B1(new_n404_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n398_), .A2(new_n392_), .ZN(new_n430_));
  NOR4_X1   g229(.A1(new_n325_), .A2(new_n257_), .A3(new_n430_), .A4(new_n373_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT73), .B(G15gat), .Z(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(G22gat), .ZN(new_n435_));
  INV_X1    g234(.A(G1gat), .ZN(new_n436_));
  INV_X1    g235(.A(G8gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT14), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT73), .B(G15gat), .ZN(new_n439_));
  INV_X1    g238(.A(G22gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n435_), .A2(new_n438_), .A3(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G1gat), .B(G8gat), .Z(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n435_), .A2(new_n443_), .A3(new_n438_), .A4(new_n441_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G29gat), .B(G36gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G43gat), .B(G50gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G229gat), .A2(G233gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n450_), .B(KEYINPUT15), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n451_), .B(new_n452_), .C1(new_n454_), .C2(new_n447_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n445_), .A2(new_n446_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(new_n450_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n455_), .B1(new_n452_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G113gat), .B(G141gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G169gat), .B(G197gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n461_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n455_), .B(new_n463_), .C1(new_n452_), .C2(new_n457_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n433_), .A2(KEYINPUT98), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT98), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n408_), .A2(new_n413_), .B1(new_n418_), .B2(new_n426_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n400_), .B(new_n403_), .C1(new_n468_), .C2(new_n373_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n431_), .B1(new_n469_), .B2(new_n257_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n465_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n467_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(KEYINPUT5), .B(G176gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT69), .B(G204gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G120gat), .B(G148gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G230gat), .A2(G233gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT7), .ZN(new_n479_));
  INV_X1    g278(.A(G99gat), .ZN(new_n480_));
  INV_X1    g279(.A(G106gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n482_), .A2(new_n485_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(G85gat), .A2(G92gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G85gat), .A2(G92gat), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT8), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT8), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n488_), .A2(new_n494_), .A3(new_n491_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n480_), .A2(KEYINPUT10), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT10), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G99gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT64), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n497_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n500_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n481_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n489_), .A2(KEYINPUT9), .A3(new_n490_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n490_), .A2(KEYINPUT9), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n505_), .A2(new_n485_), .A3(new_n506_), .A4(new_n486_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(G57gat), .A2(G64gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(G57gat), .A2(G64gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT11), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT65), .ZN(new_n513_));
  OR3_X1    g312(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT11), .ZN(new_n514_));
  XOR2_X1   g313(.A(G71gat), .B(G78gat), .Z(new_n515_));
  INV_X1    g314(.A(KEYINPUT65), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n516_), .B(KEYINPUT11), .C1(new_n510_), .C2(new_n511_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .A4(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n515_), .B1(KEYINPUT11), .B2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n516_), .B1(new_n519_), .B2(KEYINPUT11), .ZN(new_n521_));
  INV_X1    g320(.A(new_n517_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n496_), .A2(new_n509_), .A3(new_n518_), .A4(new_n523_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n488_), .A2(new_n494_), .A3(new_n491_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n494_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n498_), .A2(G99gat), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n480_), .A2(KEYINPUT10), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT64), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(G106gat), .B1(new_n529_), .B2(new_n501_), .ZN(new_n530_));
  OAI22_X1  g329(.A1(new_n525_), .A2(new_n526_), .B1(new_n530_), .B2(new_n507_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n523_), .A2(new_n518_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n478_), .B1(new_n524_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT66), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT68), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n531_), .A2(new_n532_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n478_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n536_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  OAI211_X1 g338(.A(KEYINPUT68), .B(new_n478_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n533_), .A2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT67), .B1(new_n525_), .B2(new_n526_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n493_), .A2(new_n545_), .A3(new_n495_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n546_), .A3(new_n509_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(KEYINPUT12), .A3(new_n532_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n541_), .A2(new_n543_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n477_), .B1(new_n535_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT13), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n535_), .A2(new_n549_), .A3(new_n477_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n535_), .A2(new_n549_), .A3(new_n477_), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT13), .B1(new_n555_), .B2(new_n550_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT37), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n547_), .A2(new_n453_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT34), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(KEYINPUT35), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n493_), .A2(new_n495_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n567_), .B2(new_n450_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n563_), .A2(KEYINPUT72), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT71), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n565_), .A2(KEYINPUT35), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n572_), .B(KEYINPUT70), .Z(new_n573_));
  NAND3_X1  g372(.A1(new_n563_), .A2(KEYINPUT71), .A3(new_n568_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n571_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n573_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n569_), .A2(new_n570_), .A3(new_n576_), .ZN(new_n577_));
  AOI211_X1 g376(.A(KEYINPUT36), .B(new_n562_), .C1(new_n575_), .C2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n562_), .A2(KEYINPUT36), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n562_), .A2(KEYINPUT36), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n575_), .A2(new_n580_), .A3(new_n581_), .A4(new_n577_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n558_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(G211gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT16), .B(G183gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT17), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n445_), .A2(new_n590_), .A3(new_n446_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n592_));
  OR3_X1    g391(.A1(new_n591_), .A2(new_n592_), .A3(new_n532_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n532_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n589_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n588_), .A2(KEYINPUT17), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT74), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n593_), .A2(new_n594_), .A3(KEYINPUT74), .A4(new_n596_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n595_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n601_), .A2(KEYINPUT75), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT75), .ZN(new_n603_));
  AOI211_X1 g402(.A(new_n603_), .B(new_n595_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n575_), .A2(new_n581_), .A3(new_n577_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n579_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(KEYINPUT37), .A3(new_n582_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n584_), .A2(new_n605_), .A3(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n466_), .A2(new_n472_), .A3(new_n557_), .A4(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n430_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n612_));
  OR4_X1    g411(.A1(G1gat), .A2(new_n610_), .A3(new_n611_), .A4(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n610_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n436_), .A3(new_n430_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n612_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n607_), .A2(KEYINPUT101), .A3(new_n582_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT101), .B1(new_n607_), .B2(new_n582_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n470_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n557_), .A2(new_n605_), .A3(new_n465_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT100), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G1gat), .B1(new_n624_), .B2(new_n611_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n613_), .A2(new_n616_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT102), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n613_), .A2(new_n616_), .A3(new_n628_), .A4(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(G1324gat));
  XNOR2_X1  g429(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n631_));
  INV_X1    g430(.A(new_n325_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G8gat), .B1(new_n624_), .B2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(KEYINPUT39), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(KEYINPUT39), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n614_), .A2(new_n437_), .A3(new_n325_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n631_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n637_), .B(new_n631_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n640_), .ZN(G1325gat));
  INV_X1    g440(.A(new_n257_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n621_), .A2(new_n642_), .A3(new_n623_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G15gat), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n644_), .A2(KEYINPUT104), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(KEYINPUT104), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n610_), .A2(G15gat), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n651_));
  OR3_X1    g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n257_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n651_), .B1(new_n650_), .B2(new_n257_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n645_), .A2(KEYINPUT41), .A3(new_n646_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n649_), .A2(new_n652_), .A3(new_n653_), .A4(new_n654_), .ZN(G1326gat));
  INV_X1    g454(.A(new_n373_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G22gat), .B1(new_n624_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT42), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n614_), .A2(new_n440_), .A3(new_n373_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1327gat));
  NOR2_X1   g459(.A1(new_n619_), .A2(new_n605_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n466_), .A2(new_n472_), .A3(new_n557_), .A4(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G29gat), .B1(new_n663_), .B2(new_n430_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n584_), .A2(new_n608_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(KEYINPUT106), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n433_), .A2(new_n665_), .A3(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n669_));
  INV_X1    g468(.A(new_n665_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n470_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n557_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n672_), .A2(new_n605_), .A3(new_n471_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n668_), .A2(new_n671_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(G29gat), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n668_), .A2(new_n671_), .A3(KEYINPUT44), .A4(new_n673_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n678_), .A2(new_n430_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n664_), .B1(new_n677_), .B2(new_n679_), .ZN(G1328gat));
  NAND2_X1  g479(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT109), .Z(new_n682_));
  NAND3_X1  g481(.A1(new_n676_), .A2(new_n325_), .A3(new_n678_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n466_), .A2(new_n472_), .A3(new_n557_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n632_), .A2(G36gat), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n684_), .A2(new_n661_), .A3(new_n685_), .A4(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n685_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n686_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n662_), .B2(new_n689_), .ZN(new_n690_));
  AOI22_X1  g489(.A1(new_n683_), .A2(G36gat), .B1(new_n687_), .B2(new_n690_), .ZN(new_n691_));
  OR2_X1    g490(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n682_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n683_), .A2(G36gat), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n687_), .A2(new_n690_), .ZN(new_n695_));
  AND4_X1   g494(.A1(new_n692_), .A2(new_n694_), .A3(new_n695_), .A4(new_n682_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n693_), .A2(new_n696_), .ZN(G1329gat));
  NAND4_X1  g496(.A1(new_n676_), .A2(G43gat), .A3(new_n642_), .A4(new_n678_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n662_), .A2(new_n257_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(G43gat), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g500(.A(G50gat), .B1(new_n663_), .B2(new_n373_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n676_), .A2(G50gat), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n678_), .A2(new_n373_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(G1331gat));
  NOR2_X1   g504(.A1(new_n470_), .A2(new_n465_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n609_), .A2(new_n672_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT110), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G57gat), .B1(new_n710_), .B2(new_n430_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT111), .ZN(new_n712_));
  INV_X1    g511(.A(G57gat), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n557_), .A2(new_n465_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n621_), .A2(new_n605_), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n713_), .B1(new_n430_), .B2(new_n712_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n711_), .B1(new_n714_), .B2(new_n718_), .ZN(G1332gat));
  OAI21_X1  g518(.A(G64gat), .B1(new_n716_), .B2(new_n632_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT48), .Z(new_n721_));
  NOR3_X1   g520(.A1(new_n709_), .A2(G64gat), .A3(new_n632_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n716_), .B2(new_n257_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT49), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n709_), .A2(G71gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n257_), .B2(new_n726_), .ZN(G1334gat));
  OAI21_X1  g526(.A(G78gat), .B1(new_n716_), .B2(new_n656_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT50), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n709_), .A2(G78gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n656_), .B2(new_n730_), .ZN(G1335gat));
  NAND3_X1  g530(.A1(new_n706_), .A2(new_n672_), .A3(new_n661_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n430_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n605_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n668_), .A2(new_n671_), .A3(new_n735_), .A4(new_n715_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n430_), .A2(G85gat), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT112), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n734_), .B1(new_n737_), .B2(new_n739_), .ZN(G1336gat));
  AOI21_X1  g539(.A(G92gat), .B1(new_n733_), .B2(new_n325_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n736_), .A2(new_n632_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n736_), .B2(new_n257_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n733_), .B1(new_n503_), .B2(new_n502_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(new_n257_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g546(.A1(new_n733_), .A2(new_n481_), .A3(new_n373_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G106gat), .B1(new_n736_), .B2(new_n656_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(KEYINPUT52), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(G106gat), .C1(new_n736_), .C2(new_n656_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n748_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT53), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(new_n748_), .C1(new_n750_), .C2(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1339gat));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n609_), .A2(new_n759_), .A3(new_n471_), .A4(new_n557_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n584_), .A2(new_n557_), .A3(new_n605_), .A4(new_n608_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT54), .B1(new_n761_), .B2(new_n465_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT68), .B1(new_n524_), .B2(new_n478_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n540_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n548_), .A2(new_n543_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n538_), .B1(new_n768_), .B2(new_n537_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n541_), .A2(KEYINPUT55), .A3(new_n543_), .A4(new_n548_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n769_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n477_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT56), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n772_), .A2(new_n776_), .A3(new_n773_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n452_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n451_), .B(new_n778_), .C1(new_n454_), .C2(new_n447_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n461_), .C1(new_n778_), .C2(new_n457_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n464_), .A2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n775_), .A2(new_n553_), .A3(new_n777_), .A4(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT58), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n782_), .A2(new_n783_), .A3(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n665_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n772_), .A2(new_n789_), .A3(new_n776_), .A4(new_n773_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n465_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n772_), .A2(new_n773_), .B1(new_n789_), .B2(new_n776_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n791_), .A2(new_n555_), .A3(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n781_), .B1(new_n555_), .B2(new_n550_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n781_), .B(KEYINPUT114), .C1(new_n555_), .C2(new_n550_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n619_), .B1(new_n793_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n789_), .A2(new_n776_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n774_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n553_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n796_), .B(new_n797_), .C1(new_n804_), .C2(new_n791_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(KEYINPUT57), .A3(new_n619_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n788_), .A2(new_n801_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n763_), .B1(new_n807_), .B2(new_n735_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n632_), .A2(new_n430_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n257_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n808_), .A2(new_n373_), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G113gat), .B1(new_n812_), .B2(new_n465_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT116), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n805_), .A2(KEYINPUT57), .A3(new_n619_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT57), .B1(new_n805_), .B2(new_n619_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n605_), .B1(new_n817_), .B2(new_n788_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n656_), .B(new_n810_), .C1(new_n818_), .C2(new_n763_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT59), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n807_), .A2(new_n735_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n763_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n373_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n810_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n820_), .A2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n471_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n814_), .B1(G113gat), .B2(new_n827_), .ZN(G1340gat));
  NAND3_X1  g627(.A1(new_n820_), .A2(new_n825_), .A3(new_n672_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G120gat), .ZN(new_n830_));
  INV_X1    g629(.A(G120gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n557_), .B2(KEYINPUT60), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n831_), .A2(KEYINPUT60), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n823_), .A2(new_n810_), .A3(new_n832_), .A4(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n812_), .A2(KEYINPUT117), .A3(new_n832_), .A4(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n830_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT118), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n830_), .A2(new_n838_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1341gat));
  AOI21_X1  g642(.A(G127gat), .B1(new_n812_), .B2(new_n605_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n826_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n845_), .A2(G127gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n846_), .B2(new_n605_), .ZN(G1342gat));
  AOI21_X1  g646(.A(G134gat), .B1(new_n812_), .B2(new_n620_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n665_), .A2(G134gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n845_), .B2(new_n849_), .ZN(G1343gat));
  NOR2_X1   g649(.A1(new_n808_), .A2(new_n642_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n809_), .A2(new_n656_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n471_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT119), .B(G141gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1344gat));
  NOR2_X1   g655(.A1(new_n853_), .A2(new_n557_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT120), .B(G148gat), .Z(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1345gat));
  OR3_X1    g658(.A1(new_n853_), .A2(KEYINPUT121), .A3(new_n735_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT121), .B1(new_n853_), .B2(new_n735_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT61), .B(G155gat), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1346gat));
  OAI21_X1  g664(.A(G162gat), .B1(new_n853_), .B2(new_n670_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n851_), .A2(new_n620_), .A3(new_n852_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(G162gat), .B2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT122), .ZN(G1347gat));
  NAND3_X1  g668(.A1(new_n325_), .A2(new_n642_), .A3(new_n611_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n871_), .A2(KEYINPUT123), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(KEYINPUT123), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n823_), .A2(new_n465_), .A3(new_n872_), .A4(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(G169gat), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n823_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(new_n207_), .A3(new_n465_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n874_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n877_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n877_), .A2(new_n880_), .A3(KEYINPUT124), .A4(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1348gat));
  NOR2_X1   g685(.A1(new_n878_), .A2(new_n557_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n203_), .ZN(G1349gat));
  AND2_X1   g687(.A1(new_n273_), .A2(new_n274_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(G183gat), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n879_), .B(new_n605_), .C1(new_n889_), .C2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n890_), .B(new_n226_), .C1(new_n878_), .C2(new_n735_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n892_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1350gat));
  OAI21_X1  g696(.A(G190gat), .B1(new_n878_), .B2(new_n670_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n619_), .A2(new_n271_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n878_), .B2(new_n899_), .ZN(G1351gat));
  NOR4_X1   g699(.A1(new_n808_), .A2(new_n642_), .A3(new_n399_), .A4(new_n632_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n465_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n672_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g704(.A(KEYINPUT63), .B(G211gat), .C1(new_n901_), .C2(new_n605_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n901_), .A2(new_n605_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT63), .B(G211gat), .Z(new_n908_));
  AOI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(G1354gat));
  AOI21_X1  g708(.A(G218gat), .B1(new_n901_), .B2(new_n620_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n665_), .A2(G218gat), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n911_), .B(KEYINPUT127), .Z(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n901_), .B2(new_n912_), .ZN(G1355gat));
endmodule


