//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n894_, new_n896_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_;
  XOR2_X1   g000(.A(G1gat), .B(G8gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT75), .ZN(new_n203_));
  OR2_X1    g002(.A1(G15gat), .A2(G22gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G15gat), .A2(G22gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G1gat), .A2(G8gat), .ZN(new_n206_));
  AOI22_X1  g005(.A1(new_n204_), .A2(new_n205_), .B1(KEYINPUT14), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n203_), .B(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G43gat), .A2(G50gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G43gat), .A2(G50gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n210_), .B(new_n211_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G29gat), .ZN(new_n216_));
  INV_X1    g015(.A(G36gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n211_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n218_), .B(new_n212_), .C1(new_n219_), .C2(new_n209_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n215_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n221_), .B1(new_n215_), .B2(new_n220_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n208_), .B(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT79), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G229gat), .A3(G233gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT15), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n215_), .A2(new_n220_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n221_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n215_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(KEYINPUT15), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n229_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n236_), .A2(new_n208_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n208_), .A2(new_n224_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n227_), .A2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G169gat), .B(G197gat), .Z(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT80), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n244_), .B(new_n245_), .Z(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n227_), .A2(new_n241_), .A3(new_n246_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(KEYINPUT10), .B(G99gat), .Z(new_n252_));
  INV_X1    g051(.A(G106gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G85gat), .B(G92gat), .Z(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT9), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G99gat), .A2(G106gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT6), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT6), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(G99gat), .A3(G106gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT9), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(G85gat), .A3(G92gat), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n254_), .A2(new_n256_), .A3(new_n261_), .A4(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT8), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(KEYINPUT65), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT7), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n267_), .B(KEYINPUT64), .C1(G99gat), .C2(G106gat), .ZN(new_n268_));
  INV_X1    g067(.A(G99gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n269_), .B(new_n253_), .C1(new_n270_), .C2(KEYINPUT7), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n267_), .A2(KEYINPUT64), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n268_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n258_), .A2(new_n260_), .A3(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n266_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n265_), .B1(new_n276_), .B2(new_n255_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n255_), .A2(new_n265_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n278_), .B1(new_n261_), .B2(new_n273_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n264_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n235_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n224_), .B(new_n264_), .C1(new_n277_), .C2(new_n279_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(KEYINPUT70), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G232gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT34), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n285_), .A2(KEYINPUT35), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n280_), .A2(new_n235_), .A3(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n283_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n285_), .A2(KEYINPUT35), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n281_), .A2(new_n282_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT71), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n281_), .A2(new_n294_), .A3(new_n282_), .A4(new_n291_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n289_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G190gat), .B(G218gat), .Z(new_n297_));
  XNOR2_X1  g096(.A(G134gat), .B(G162gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT36), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT36), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n299_), .A2(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n296_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT37), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n296_), .A2(KEYINPUT73), .A3(new_n300_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n303_), .A2(new_n306_), .A3(new_n307_), .A4(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n301_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n296_), .A2(new_n305_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT37), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT72), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n312_), .A2(new_n316_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT74), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G57gat), .B(G64gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT11), .ZN(new_n324_));
  XOR2_X1   g123(.A(G71gat), .B(G78gat), .Z(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n324_), .A2(new_n325_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n323_), .A2(KEYINPUT11), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n208_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G231gat), .A2(G233gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT76), .Z(new_n332_));
  XNOR2_X1  g131(.A(new_n330_), .B(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n333_), .A2(KEYINPUT77), .ZN(new_n334_));
  XOR2_X1   g133(.A(G127gat), .B(G155gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G211gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(KEYINPUT16), .B(G183gat), .Z(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT17), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n338_), .A2(KEYINPUT17), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n333_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(new_n334_), .B2(new_n339_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G120gat), .B(G148gat), .ZN(new_n346_));
  INV_X1    g145(.A(G204gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT5), .B(G176gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  INV_X1    g149(.A(KEYINPUT12), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT67), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(new_n280_), .B2(new_n329_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n280_), .A2(new_n329_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n280_), .A2(new_n329_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n354_), .B(new_n355_), .C1(KEYINPUT67), .C2(new_n351_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n353_), .B1(new_n356_), .B2(new_n352_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G230gat), .A2(G233gat), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n358_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT66), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(KEYINPUT66), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n350_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT66), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n357_), .A2(new_n358_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n360_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n350_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n368_), .A2(new_n362_), .A3(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT13), .B1(new_n364_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n361_), .A2(new_n363_), .A3(new_n350_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT13), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n369_), .B1(new_n368_), .B2(new_n362_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n345_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n322_), .A2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n251_), .B1(new_n377_), .B2(KEYINPUT78), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT20), .ZN(new_n379_));
  XOR2_X1   g178(.A(G211gat), .B(G218gat), .Z(new_n380_));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G197gat), .B(G204gat), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT21), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n382_), .A2(new_n381_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n387_), .A2(new_n384_), .A3(new_n380_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n390_));
  INV_X1    g189(.A(G176gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(G169gat), .A2(G176gat), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n392_), .A2(G169gat), .B1(new_n390_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n395_), .A2(KEYINPUT23), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(KEYINPUT83), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT83), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(G183gat), .A3(G190gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n396_), .B1(new_n400_), .B2(KEYINPUT23), .ZN(new_n401_));
  NOR2_X1   g200(.A1(G183gat), .A2(G190gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n394_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT23), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n395_), .A2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(new_n400_), .B2(new_n404_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT25), .B(G183gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT81), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT26), .ZN(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT82), .B(G190gat), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(KEYINPUT82), .A2(G190gat), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(KEYINPUT81), .A3(KEYINPUT26), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n408_), .B1(new_n409_), .B2(G190gat), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n407_), .A2(new_n410_), .A3(new_n412_), .A4(new_n413_), .ZN(new_n414_));
  NOR3_X1   g213(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G169gat), .A2(G176gat), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n415_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n406_), .A2(new_n414_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n403_), .A2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n379_), .B1(new_n389_), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT22), .B(G169gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n391_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n418_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT91), .ZN(new_n427_));
  INV_X1    g226(.A(new_n402_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n406_), .B2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT23), .B1(new_n397_), .B2(new_n399_), .ZN(new_n430_));
  NOR4_X1   g229(.A1(new_n430_), .A2(KEYINPUT91), .A3(new_n402_), .A4(new_n405_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n426_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n383_), .A2(KEYINPUT21), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n433_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n401_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT26), .B(G190gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT90), .ZN(new_n437_));
  INV_X1    g236(.A(new_n407_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n435_), .B(new_n419_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n432_), .A2(new_n434_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n422_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G226gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n441_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n400_), .A2(new_n404_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n405_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n428_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT91), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n406_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n425_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n404_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n419_), .B1(new_n453_), .B2(new_n396_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n437_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n454_), .B1(new_n455_), .B2(new_n407_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n389_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT92), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n434_), .B1(new_n432_), .B2(new_n439_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT92), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n403_), .A2(new_n420_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n379_), .B1(new_n462_), .B2(new_n434_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n458_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n446_), .B1(new_n464_), .B2(new_n445_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G64gat), .B(G92gat), .Z(new_n466_));
  XNOR2_X1  g265(.A(G8gat), .B(G36gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT32), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n465_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G225gat), .A2(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G141gat), .A2(G148gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT87), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT2), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT2), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(KEYINPUT87), .A3(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n481_));
  OR3_X1    g280(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n478_), .A2(new_n480_), .A3(new_n481_), .A4(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G155gat), .B(G162gat), .Z(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(G127gat), .ZN(new_n486_));
  INV_X1    g285(.A(G134gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(G120gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G113gat), .ZN(new_n490_));
  INV_X1    g289(.A(G113gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(G120gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G127gat), .A2(G134gat), .ZN(new_n493_));
  AND4_X1   g292(.A1(new_n488_), .A2(new_n490_), .A3(new_n492_), .A4(new_n493_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n490_), .A2(new_n492_), .B1(new_n488_), .B2(new_n493_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(G141gat), .ZN(new_n497_));
  INV_X1    g296(.A(G148gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(G155gat), .A2(G162gat), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n476_), .B(new_n499_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n485_), .A2(new_n496_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n496_), .B1(new_n485_), .B2(new_n504_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT4), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n507_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n475_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n474_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G1gat), .B(G29gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G57gat), .B(G85gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n485_), .A2(new_n504_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n496_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n485_), .A2(new_n504_), .A3(new_n496_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(KEYINPUT4), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n474_), .B1(new_n524_), .B2(new_n509_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n512_), .ZN(new_n526_));
  OR3_X1    g325(.A1(new_n525_), .A2(new_n518_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n519_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n463_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n529_));
  AOI211_X1 g328(.A(KEYINPUT92), .B(new_n434_), .C1(new_n432_), .C2(new_n439_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n445_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n422_), .A2(new_n440_), .A3(new_n444_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n471_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n473_), .A2(new_n528_), .A3(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n505_), .A2(new_n506_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n518_), .B1(new_n535_), .B2(new_n475_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n524_), .A2(new_n474_), .A3(new_n509_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT33), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n539_), .B1(new_n513_), .B2(new_n518_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n539_), .B(new_n518_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n538_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n470_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT20), .B1(new_n389_), .B2(new_n421_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n457_), .B2(KEYINPUT92), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n444_), .B1(new_n546_), .B2(new_n461_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n532_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n544_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n531_), .A2(new_n470_), .A3(new_n532_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT94), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n543_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(KEYINPUT94), .A3(new_n550_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n534_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n434_), .B1(KEYINPUT29), .B2(new_n520_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G228gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT28), .ZN(new_n558_));
  XOR2_X1   g357(.A(G22gat), .B(G50gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n556_), .B(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n520_), .A2(KEYINPUT29), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G78gat), .B(G106gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT96), .B1(new_n555_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT27), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n551_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n567_), .A2(new_n528_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n465_), .B2(new_n544_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n548_), .B1(new_n464_), .B2(new_n445_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT97), .B1(new_n574_), .B2(new_n470_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n531_), .A2(KEYINPUT97), .A3(new_n470_), .A4(new_n532_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  OAI211_X1 g376(.A(KEYINPUT98), .B(new_n573_), .C1(new_n575_), .C2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT97), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n550_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n576_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT98), .B1(new_n582_), .B2(new_n573_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n571_), .B(new_n572_), .C1(new_n579_), .C2(new_n583_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n547_), .A2(new_n544_), .A3(new_n548_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n470_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n552_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n543_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n554_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n534_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT96), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n592_), .A3(new_n567_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n569_), .A2(new_n584_), .A3(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n421_), .B(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(G71gat), .B(G99gat), .Z(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT30), .B(G43gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n596_), .B(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(KEYINPUT85), .B(G15gat), .Z(new_n601_));
  NAND2_X1  g400(.A1(G227gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n521_), .B(new_n603_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n604_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n594_), .A2(new_n608_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n571_), .B(new_n567_), .C1(new_n579_), .C2(new_n583_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT99), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n573_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n578_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n615_), .A2(new_n616_), .A3(new_n571_), .A4(new_n567_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n528_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n611_), .A2(new_n617_), .A3(new_n607_), .A4(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n609_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n322_), .A2(new_n376_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT78), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n378_), .A2(new_n620_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n378_), .A2(KEYINPUT100), .A3(new_n620_), .A4(new_n623_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(G1gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n528_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n311_), .B1(new_n302_), .B2(new_n301_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n308_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AOI211_X1 g434(.A(new_n635_), .B(new_n345_), .C1(new_n609_), .C2(new_n619_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n371_), .A2(new_n375_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n250_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT101), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G1gat), .B1(new_n640_), .B2(new_n618_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n630_), .A2(new_n631_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n632_), .A2(new_n641_), .A3(new_n642_), .ZN(G1324gat));
  XNOR2_X1  g442(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT40), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n615_), .A2(new_n571_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(G8gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n628_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT102), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n628_), .A2(new_n652_), .A3(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G8gat), .B1(new_n640_), .B2(new_n648_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT39), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n657_), .B(G8gat), .C1(new_n640_), .C2(new_n648_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n646_), .B1(new_n654_), .B2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n652_), .B1(new_n628_), .B2(new_n649_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n649_), .ZN(new_n662_));
  AOI211_X1 g461(.A(KEYINPUT102), .B(new_n662_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n646_), .B(new_n659_), .C1(new_n661_), .C2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n645_), .B1(new_n660_), .B2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n659_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT40), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(new_n664_), .A3(new_n644_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(G1325gat));
  OAI21_X1  g469(.A(G15gat), .B1(new_n640_), .B2(new_n608_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n671_), .A2(KEYINPUT41), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(KEYINPUT41), .ZN(new_n673_));
  OR3_X1    g472(.A1(new_n624_), .A2(G15gat), .A3(new_n608_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(G1326gat));
  OAI21_X1  g474(.A(G22gat), .B1(new_n640_), .B2(new_n567_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT42), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n567_), .A2(G22gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(new_n624_), .B2(new_n678_), .ZN(G1327gat));
  INV_X1    g478(.A(new_n345_), .ZN(new_n680_));
  AOI211_X1 g479(.A(new_n634_), .B(new_n680_), .C1(new_n609_), .C2(new_n619_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n638_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n216_), .A3(new_n528_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n639_), .A2(new_n345_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n687_));
  AOI211_X1 g486(.A(KEYINPUT43), .B(new_n322_), .C1(new_n609_), .C2(new_n619_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n315_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n319_), .A2(new_n320_), .A3(KEYINPUT74), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n318_), .A2(new_n321_), .A3(KEYINPUT105), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n689_), .B1(new_n695_), .B2(new_n620_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n688_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  AOI22_X1  g497(.A1(new_n694_), .A2(new_n693_), .B1(new_n609_), .B2(new_n619_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT106), .B1(new_n699_), .B2(new_n689_), .ZN(new_n700_));
  AOI211_X1 g499(.A(new_n686_), .B(new_n687_), .C1(new_n698_), .C2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n687_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n609_), .A2(new_n619_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n318_), .A2(KEYINPUT105), .A3(new_n321_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT105), .B1(new_n318_), .B2(new_n321_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n697_), .B(KEYINPUT43), .C1(new_n703_), .C2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n688_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n700_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n686_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n702_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n701_), .A2(new_n711_), .A3(new_n618_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n685_), .B1(new_n712_), .B2(new_n216_), .ZN(G1328gat));
  NOR2_X1   g512(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT110), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n683_), .A2(G36gat), .A3(new_n648_), .ZN(new_n717_));
  XOR2_X1   g516(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n709_), .A2(new_n710_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n687_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n709_), .A2(new_n710_), .A3(new_n702_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n647_), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n719_), .B1(new_n723_), .B2(G36gat), .ZN(new_n724_));
  NAND2_X1  g523(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n716_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n701_), .A2(new_n711_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n217_), .B1(new_n728_), .B2(new_n647_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n725_), .B(new_n715_), .C1(new_n729_), .C2(new_n719_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n727_), .A2(new_n730_), .ZN(G1329gat));
  NOR3_X1   g530(.A1(new_n701_), .A2(new_n711_), .A3(new_n608_), .ZN(new_n732_));
  INV_X1    g531(.A(G43gat), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n607_), .A2(new_n733_), .ZN(new_n734_));
  OAI22_X1  g533(.A1(new_n732_), .A2(new_n733_), .B1(new_n683_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(G1330gat));
  NOR3_X1   g536(.A1(new_n701_), .A2(new_n711_), .A3(new_n567_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n738_), .A2(KEYINPUT111), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(KEYINPUT111), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(G50gat), .A3(new_n740_), .ZN(new_n741_));
  OR3_X1    g540(.A1(new_n683_), .A2(G50gat), .A3(new_n567_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1331gat));
  NOR2_X1   g542(.A1(new_n637_), .A2(new_n250_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n636_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(G57gat), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n745_), .A2(new_n746_), .A3(new_n618_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n620_), .A2(new_n322_), .A3(new_n680_), .A4(new_n744_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n618_), .B1(new_n748_), .B2(KEYINPUT112), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(KEYINPUT112), .B2(new_n748_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n747_), .B1(new_n750_), .B2(new_n746_), .ZN(G1332gat));
  OAI21_X1  g550(.A(G64gat), .B1(new_n745_), .B2(new_n648_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT48), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n648_), .A2(G64gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n748_), .B2(new_n754_), .ZN(G1333gat));
  OAI21_X1  g554(.A(G71gat), .B1(new_n745_), .B2(new_n608_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT49), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n608_), .A2(G71gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n748_), .B2(new_n758_), .ZN(G1334gat));
  OAI21_X1  g558(.A(G78gat), .B1(new_n745_), .B2(new_n567_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT50), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n567_), .A2(G78gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n748_), .B2(new_n762_), .ZN(G1335gat));
  NAND2_X1  g562(.A1(new_n681_), .A2(new_n744_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT113), .Z(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(G85gat), .B1(new_n766_), .B2(new_n528_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n709_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n744_), .A2(new_n345_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n528_), .A2(G85gat), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT114), .Z(new_n772_));
  AOI21_X1  g571(.A(new_n767_), .B1(new_n770_), .B2(new_n772_), .ZN(G1336gat));
  NOR3_X1   g572(.A1(new_n765_), .A2(G92gat), .A3(new_n648_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n770_), .A2(new_n647_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(G92gat), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT115), .ZN(G1337gat));
  NAND3_X1  g576(.A1(new_n766_), .A2(new_n607_), .A3(new_n252_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n768_), .A2(new_n608_), .A3(new_n769_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n269_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g580(.A1(new_n766_), .A2(new_n253_), .A3(new_n568_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n709_), .A2(new_n568_), .A3(new_n345_), .A4(new_n744_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n783_), .A2(new_n784_), .A3(G106gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n783_), .B2(G106gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  XOR2_X1   g586(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(G1339gat));
  AND3_X1   g588(.A1(new_n611_), .A2(new_n607_), .A3(new_n617_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT55), .B1(new_n357_), .B2(new_n358_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT117), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n793_), .B(KEYINPUT55), .C1(new_n357_), .C2(new_n358_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n359_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n369_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n359_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT56), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n792_), .A2(new_n794_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n366_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n369_), .A4(new_n795_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n798_), .A2(new_n802_), .A3(new_n372_), .A4(new_n250_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n226_), .A2(new_n240_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n239_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n804_), .B(new_n247_), .C1(new_n240_), .C2(new_n805_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n806_), .A2(new_n249_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n364_), .B2(new_n370_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n803_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT57), .B1(new_n809_), .B2(new_n634_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n811_));
  AOI211_X1 g610(.A(new_n811_), .B(new_n635_), .C1(new_n803_), .C2(new_n808_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n798_), .A2(new_n802_), .A3(new_n372_), .A4(new_n807_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT58), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n322_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n815_), .B2(new_n814_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n680_), .B1(new_n813_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n377_), .A2(new_n251_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n528_), .B(new_n790_), .C1(new_n818_), .C2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT118), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n809_), .A2(new_n634_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n811_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n809_), .A2(KEYINPUT57), .A3(new_n634_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n817_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n345_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n819_), .B(KEYINPUT54), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n528_), .A4(new_n790_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n250_), .B1(new_n824_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n822_), .B1(new_n836_), .B2(KEYINPUT59), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n618_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n790_), .A3(new_n840_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n837_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n251_), .A2(new_n491_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n835_), .A2(new_n491_), .B1(new_n842_), .B2(new_n843_), .ZN(G1340gat));
  OAI21_X1  g643(.A(new_n489_), .B1(new_n637_), .B2(KEYINPUT60), .ZN(new_n845_));
  OAI221_X1 g644(.A(new_n845_), .B1(KEYINPUT60), .B2(new_n489_), .C1(new_n824_), .C2(new_n834_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n637_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n837_), .A2(new_n847_), .A3(new_n841_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(G120gat), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n848_), .A2(new_n849_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n846_), .B1(new_n851_), .B2(new_n852_), .ZN(G1341gat));
  NAND2_X1  g652(.A1(new_n680_), .A2(G127gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT121), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n837_), .A2(new_n841_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n345_), .B1(new_n823_), .B2(new_n833_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(G127gat), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n856_), .B(KEYINPUT122), .C1(new_n857_), .C2(G127gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1342gat));
  OAI21_X1  g661(.A(new_n635_), .B1(new_n824_), .B2(new_n834_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n487_), .A2(KEYINPUT123), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n487_), .A2(KEYINPUT123), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n322_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n863_), .A2(new_n487_), .B1(new_n842_), .B2(new_n866_), .ZN(G1343gat));
  NOR3_X1   g666(.A1(new_n647_), .A2(new_n607_), .A3(new_n567_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n838_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n251_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n497_), .ZN(G1344gat));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n637_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(new_n498_), .ZN(G1345gat));
  NOR2_X1   g672(.A1(new_n869_), .A2(new_n345_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT61), .B(G155gat), .Z(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  INV_X1    g675(.A(new_n869_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n877_), .A2(G162gat), .A3(new_n695_), .ZN(new_n878_));
  AOI21_X1  g677(.A(G162gat), .B1(new_n877_), .B2(new_n635_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1347gat));
  AOI211_X1 g679(.A(new_n648_), .B(new_n528_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n608_), .A2(new_n568_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n250_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n884_), .A3(G169gat), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n883_), .B2(G169gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n881_), .A2(new_n882_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n250_), .A2(new_n423_), .ZN(new_n889_));
  XOR2_X1   g688(.A(new_n889_), .B(KEYINPUT124), .Z(new_n890_));
  OAI22_X1  g689(.A1(new_n886_), .A2(new_n887_), .B1(new_n888_), .B2(new_n890_), .ZN(G1348gat));
  NOR2_X1   g690(.A1(new_n888_), .A2(new_n637_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n391_), .ZN(G1349gat));
  NAND3_X1  g692(.A1(new_n881_), .A2(new_n680_), .A3(new_n882_), .ZN(new_n894_));
  MUX2_X1   g693(.A(new_n407_), .B(G183gat), .S(new_n894_), .Z(G1350gat));
  OAI21_X1  g694(.A(G190gat), .B1(new_n888_), .B2(new_n322_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n634_), .A2(new_n437_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT125), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n888_), .B2(new_n898_), .ZN(G1351gat));
  NOR2_X1   g698(.A1(new_n607_), .A2(new_n567_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n881_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n250_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n847_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n347_), .A2(KEYINPUT126), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n347_), .A2(KEYINPUT126), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n905_), .B2(new_n906_), .ZN(G1353gat));
  AOI21_X1  g708(.A(new_n345_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT127), .Z(new_n911_));
  NOR2_X1   g710(.A1(new_n901_), .A2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1354gat));
  INV_X1    g713(.A(G218gat), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n901_), .A2(new_n915_), .A3(new_n322_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n902_), .A2(new_n635_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n915_), .B2(new_n917_), .ZN(G1355gat));
endmodule


