//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n891_, new_n892_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_;
  XOR2_X1   g000(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(KEYINPUT1), .B2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(KEYINPUT1), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n207_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n206_), .B(KEYINPUT2), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT82), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(G141gat), .B2(G148gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT3), .B1(new_n215_), .B2(KEYINPUT83), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT82), .B1(KEYINPUT83), .B2(KEYINPUT3), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n205_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n213_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n209_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(new_n208_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n212_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT29), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n223_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n202_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n227_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n202_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n225_), .A3(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G22gat), .B(G50gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n228_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n233_), .B1(new_n228_), .B2(new_n231_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G204gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT87), .B1(new_n237_), .B2(G197gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT87), .ZN(new_n239_));
  INV_X1    g038(.A(G197gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(G204gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT21), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(G197gat), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n238_), .A2(new_n241_), .A3(new_n242_), .A4(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n237_), .A2(G197gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n240_), .A2(G204gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT21), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G218gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G211gat), .ZN(new_n249_));
  INV_X1    g048(.A(G211gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G218gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT88), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n249_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n252_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n244_), .B(new_n247_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n249_), .A2(new_n251_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT88), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n238_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n249_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(KEYINPUT21), .A4(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT89), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n255_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n261_), .B1(new_n255_), .B2(new_n260_), .ZN(new_n263_));
  INV_X1    g062(.A(G233gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT86), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n265_), .A2(G228gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(G228gat), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n264_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NOR3_X1   g068(.A1(new_n262_), .A2(new_n263_), .A3(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(new_n224_), .B2(new_n222_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT90), .ZN(new_n272_));
  INV_X1    g071(.A(new_n221_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT83), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n205_), .B2(new_n214_), .ZN(new_n275_));
  OAI22_X1  g074(.A1(new_n275_), .A2(KEYINPUT3), .B1(new_n205_), .B2(new_n217_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n273_), .B1(new_n276_), .B2(new_n213_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n272_), .B(KEYINPUT29), .C1(new_n277_), .C2(new_n212_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT90), .B1(new_n222_), .B2(new_n224_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n255_), .A2(new_n260_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n281_), .A2(KEYINPUT91), .A3(new_n269_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT91), .B1(new_n281_), .B2(new_n269_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n271_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G78gat), .B(G106gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT92), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n286_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n288_), .B(new_n271_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n236_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n287_), .A2(new_n236_), .A3(new_n289_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G226gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT94), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n296_));
  XOR2_X1   g095(.A(new_n295_), .B(new_n296_), .Z(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT20), .ZN(new_n299_));
  NOR3_X1   g098(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n300_));
  INV_X1    g099(.A(G183gat), .ZN(new_n301_));
  INV_X1    g100(.A(G190gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT23), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(G183gat), .A3(G190gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n300_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n307_));
  INV_X1    g106(.A(G169gat), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT76), .B1(G169gat), .B2(G176gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n310_), .A2(KEYINPUT24), .A3(new_n311_), .A4(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n302_), .A2(KEYINPUT26), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT26), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G190gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G183gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n301_), .A2(KEYINPUT25), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n314_), .A2(new_n316_), .A3(new_n318_), .A4(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n306_), .A2(new_n313_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n305_), .A2(KEYINPUT77), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT77), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n323_), .A2(new_n304_), .A3(G183gat), .A4(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n325_), .A2(new_n303_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT22), .B(G169gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n309_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n312_), .B(KEYINPUT95), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n321_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n299_), .B1(new_n331_), .B2(new_n280_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n303_), .A2(new_n305_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n301_), .A2(new_n302_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(G169gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n310_), .A2(new_n311_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT24), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  OR3_X1    g141(.A1(new_n301_), .A2(KEYINPUT75), .A3(KEYINPUT25), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT26), .B(G190gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT25), .B1(new_n301_), .B2(KEYINPUT75), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n342_), .A2(new_n346_), .A3(new_n313_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n303_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n339_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n280_), .A2(KEYINPUT89), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n255_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n298_), .B1(new_n333_), .B2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G8gat), .B(G36gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G64gat), .B(G92gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n306_), .A2(new_n313_), .A3(new_n320_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n325_), .A2(new_n303_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n335_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n330_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n360_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n280_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n299_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n351_), .A2(new_n352_), .A3(new_n350_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n297_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n354_), .A2(new_n359_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT101), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT101), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n354_), .A2(new_n371_), .A3(new_n359_), .A4(new_n368_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n359_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n333_), .A2(new_n353_), .A3(new_n298_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n297_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n373_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n370_), .A2(new_n372_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT27), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n366_), .A2(new_n297_), .A3(new_n367_), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n347_), .A2(new_n349_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n380_), .B(new_n339_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n297_), .B1(new_n381_), .B2(new_n332_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n373_), .B1(new_n379_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT27), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n383_), .A2(new_n384_), .A3(new_n369_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n378_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388_));
  INV_X1    g187(.A(G15gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(G43gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n391_), .B(new_n392_), .Z(new_n393_));
  INV_X1    g192(.A(KEYINPUT78), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n350_), .B(KEYINPUT30), .Z(new_n396_));
  XNOR2_X1  g195(.A(new_n391_), .B(new_n392_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT78), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n395_), .A2(new_n396_), .A3(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n350_), .B(KEYINPUT30), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(KEYINPUT80), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G134gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(G127gat), .ZN(new_n404_));
  INV_X1    g203(.A(G127gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G134gat), .ZN(new_n406_));
  INV_X1    g205(.A(G120gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G113gat), .ZN(new_n408_));
  INV_X1    g207(.A(G113gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(G120gat), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n404_), .A2(new_n406_), .A3(new_n408_), .A4(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT79), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G113gat), .B(G120gat), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n414_), .A2(KEYINPUT79), .A3(new_n404_), .A4(new_n406_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n404_), .A2(new_n406_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n408_), .A2(new_n410_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n413_), .A2(new_n415_), .A3(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n419_), .B(KEYINPUT31), .Z(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n402_), .B(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n219_), .A2(new_n221_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n212_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n419_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n418_), .A2(new_n411_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n222_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n424_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT4), .B1(new_n427_), .B2(new_n428_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n419_), .B2(new_n222_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(KEYINPUT4), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n432_), .B1(new_n435_), .B2(new_n424_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G1gat), .B(G29gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(G85gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT0), .B(G57gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  AOI221_X4 g240(.A(new_n212_), .B1(new_n411_), .B2(new_n418_), .C1(new_n219_), .C2(new_n221_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n419_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT4), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT4), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n429_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n424_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n432_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n440_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n441_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n422_), .A2(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n293_), .A2(new_n387_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT97), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(KEYINPUT33), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n456_), .ZN(new_n458_));
  AOI211_X1 g257(.A(new_n440_), .B(new_n458_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n429_), .A2(new_n431_), .A3(new_n424_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n440_), .B(new_n461_), .C1(new_n435_), .C2(new_n424_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n383_), .A2(new_n462_), .A3(new_n369_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT98), .B1(new_n460_), .B2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n458_), .B1(new_n436_), .B2(new_n440_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n449_), .A2(new_n450_), .A3(new_n456_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n383_), .A2(new_n369_), .A3(new_n462_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT98), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n359_), .A2(KEYINPUT32), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n354_), .A2(new_n368_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT99), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT99), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n354_), .A2(new_n474_), .A3(new_n368_), .A4(new_n471_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n471_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n477_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT100), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT100), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n480_), .B(new_n477_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n476_), .A2(new_n452_), .A3(new_n479_), .A4(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n464_), .A2(new_n470_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n293_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n452_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n387_), .A2(new_n291_), .A3(new_n485_), .A4(new_n292_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n422_), .B(KEYINPUT81), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n454_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT6), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G85gat), .A2(G92gat), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n493_), .A2(KEYINPUT9), .ZN(new_n494_));
  OR2_X1    g293(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n495_));
  INV_X1    g294(.A(G106gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G85gat), .ZN(new_n499_));
  INV_X1    g298(.A(G92gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(KEYINPUT9), .A3(new_n493_), .ZN(new_n502_));
  AND4_X1   g301(.A1(new_n492_), .A2(new_n494_), .A3(new_n498_), .A4(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT7), .ZN(new_n505_));
  INV_X1    g304(.A(G99gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(new_n496_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n492_), .A2(new_n504_), .A3(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n501_), .A2(new_n493_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT64), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT8), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n503_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n508_), .A2(KEYINPUT64), .A3(new_n509_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n491_), .B(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(new_n504_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n509_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT64), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n513_), .A2(new_n519_), .A3(KEYINPUT8), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G57gat), .B(G64gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT11), .ZN(new_n522_));
  XOR2_X1   g321(.A(G71gat), .B(G78gat), .Z(new_n523_));
  OR2_X1    g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n521_), .A2(KEYINPUT11), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n523_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n524_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n512_), .A2(new_n520_), .A3(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(KEYINPUT65), .A2(KEYINPUT12), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G230gat), .A2(G233gat), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n527_), .B1(new_n512_), .B2(new_n520_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(KEYINPUT65), .A2(KEYINPUT12), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT65), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT12), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  AOI211_X1 g336(.A(new_n527_), .B(new_n537_), .C1(new_n512_), .C2(new_n520_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n530_), .B(new_n531_), .C1(new_n534_), .C2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n528_), .ZN(new_n540_));
  OAI211_X1 g339(.A(G230gat), .B(G233gat), .C1(new_n540_), .C2(new_n532_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G120gat), .B(G148gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT5), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G176gat), .B(G204gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n546_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT66), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(KEYINPUT66), .A3(new_n548_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT13), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G1gat), .B(G8gat), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT73), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(G22gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n389_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G15gat), .A2(G22gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G1gat), .A2(G8gat), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n560_), .A2(new_n561_), .B1(KEYINPUT14), .B2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n558_), .B(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G29gat), .B(G36gat), .Z(new_n565_));
  XOR2_X1   g364(.A(G43gat), .B(G50gat), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G29gat), .B(G36gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G43gat), .B(G50gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n564_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT15), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n567_), .A2(KEYINPUT15), .A3(new_n570_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n572_), .B1(new_n564_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G229gat), .A2(G233gat), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n564_), .B(new_n571_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n579_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G113gat), .B(G141gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(G169gat), .B(G197gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n586_), .A2(KEYINPUT74), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n583_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n551_), .A2(KEYINPUT13), .A3(new_n552_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n555_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n490_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT37), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT72), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT36), .Z(new_n598_));
  NAND3_X1  g397(.A1(new_n512_), .A2(new_n520_), .A3(new_n571_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n600_));
  AND2_X1   g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT35), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT69), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT69), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n602_), .A2(new_n606_), .A3(new_n603_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n602_), .A2(new_n603_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n605_), .A2(new_n607_), .B1(KEYINPUT70), .B2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n599_), .A2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n576_), .B1(new_n512_), .B2(new_n520_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT68), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  AOI211_X1 g412(.A(KEYINPUT68), .B(new_n576_), .C1(new_n512_), .C2(new_n520_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n610_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n608_), .A2(KEYINPUT70), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT71), .ZN(new_n618_));
  OAI221_X1 g417(.A(new_n610_), .B1(KEYINPUT70), .B2(new_n608_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n618_), .B1(new_n617_), .B2(new_n619_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n594_), .B(new_n598_), .C1(new_n620_), .C2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n619_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n597_), .A2(KEYINPUT36), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(KEYINPUT71), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n617_), .A2(new_n619_), .A3(new_n618_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n594_), .B1(new_n629_), .B2(new_n598_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n593_), .B1(new_n626_), .B2(new_n630_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n617_), .A2(new_n598_), .A3(new_n619_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(KEYINPUT37), .A3(new_n625_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n527_), .B(new_n636_), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(new_n564_), .ZN(new_n638_));
  XOR2_X1   g437(.A(G127gat), .B(G155gat), .Z(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT16), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G183gat), .B(G211gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT17), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n638_), .A2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n642_), .B(new_n643_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n638_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n635_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n592_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(G1gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(new_n652_), .A3(new_n452_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT38), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n598_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT72), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(new_n622_), .A3(new_n625_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n649_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n592_), .A2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT102), .Z(new_n661_));
  AND2_X1   g460(.A1(new_n661_), .A2(new_n452_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n654_), .B1(new_n662_), .B2(new_n652_), .ZN(G1324gat));
  OAI21_X1  g462(.A(G8gat), .B1(new_n660_), .B2(new_n387_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT39), .ZN(new_n665_));
  INV_X1    g464(.A(G8gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n385_), .B1(new_n377_), .B2(KEYINPUT27), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n651_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(G1325gat));
  NAND3_X1  g470(.A1(new_n651_), .A2(new_n389_), .A3(new_n488_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n389_), .B1(new_n661_), .B2(new_n488_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n673_), .A2(KEYINPUT41), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(KEYINPUT41), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n674_), .B2(new_n675_), .ZN(G1326gat));
  INV_X1    g475(.A(new_n293_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n651_), .A2(new_n559_), .A3(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n559_), .B1(new_n661_), .B2(new_n677_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n679_), .A2(new_n680_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(G1327gat));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n684_), .A2(KEYINPUT43), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(KEYINPUT43), .ZN(new_n686_));
  INV_X1    g485(.A(new_n634_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n657_), .B2(new_n593_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n685_), .B(new_n686_), .C1(new_n490_), .C2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n293_), .A2(new_n453_), .A3(new_n387_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n287_), .A2(new_n236_), .A3(new_n289_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n667_), .A2(new_n691_), .A3(new_n290_), .ZN(new_n692_));
  AOI22_X1  g491(.A1(new_n692_), .A2(new_n485_), .B1(new_n483_), .B2(new_n293_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n690_), .B1(new_n693_), .B2(new_n488_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n694_), .A2(new_n684_), .A3(KEYINPUT43), .A4(new_n635_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n591_), .A2(new_n648_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n689_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n689_), .A2(new_n695_), .A3(KEYINPUT44), .A4(new_n696_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n452_), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G29gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n657_), .A2(new_n648_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n592_), .A2(new_n703_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n485_), .A2(G29gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n702_), .B1(new_n704_), .B2(new_n705_), .ZN(G1328gat));
  NOR2_X1   g505(.A1(new_n387_), .A2(G36gat), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT106), .B1(new_n704_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n592_), .A2(new_n710_), .A3(new_n703_), .A4(new_n707_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n709_), .A2(KEYINPUT45), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT45), .B1(new_n709_), .B2(new_n711_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n699_), .A2(new_n667_), .A3(new_n700_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n699_), .A2(KEYINPUT105), .A3(new_n667_), .A4(new_n700_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G36gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n714_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT46), .B(new_n714_), .C1(new_n717_), .C2(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1329gat));
  INV_X1    g523(.A(G43gat), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n422_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n699_), .A2(new_n700_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT107), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n699_), .A2(new_n729_), .A3(new_n700_), .A4(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n725_), .B1(new_n704_), .B2(new_n489_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT108), .Z(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT47), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n731_), .A2(new_n736_), .A3(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1330gat));
  OR3_X1    g537(.A1(new_n704_), .A2(G50gat), .A3(new_n293_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n699_), .A2(new_n677_), .A3(new_n700_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(new_n741_), .A3(G50gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n740_), .B2(G50gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(G1331gat));
  NAND2_X1  g543(.A1(new_n555_), .A2(new_n590_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n588_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(new_n490_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n659_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G57gat), .B1(new_n748_), .B2(new_n485_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n650_), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n485_), .A2(G57gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(G1332gat));
  OAI21_X1  g551(.A(G64gat), .B1(new_n748_), .B2(new_n387_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT48), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n387_), .A2(G64gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n750_), .B2(new_n755_), .ZN(G1333gat));
  OAI21_X1  g555(.A(G71gat), .B1(new_n748_), .B2(new_n489_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT49), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n489_), .A2(G71gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n750_), .B2(new_n759_), .ZN(G1334gat));
  INV_X1    g559(.A(G78gat), .ZN(new_n761_));
  INV_X1    g560(.A(new_n748_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(new_n677_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n763_), .A2(new_n764_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n293_), .A2(G78gat), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT111), .ZN(new_n769_));
  OAI22_X1  g568(.A1(new_n766_), .A2(new_n767_), .B1(new_n750_), .B2(new_n769_), .ZN(G1335gat));
  AND2_X1   g569(.A1(new_n689_), .A2(new_n695_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n746_), .A2(new_n648_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773_), .B2(new_n485_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n747_), .A2(new_n703_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n499_), .A3(new_n452_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n774_), .A2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT112), .ZN(G1336gat));
  OAI21_X1  g578(.A(G92gat), .B1(new_n773_), .B2(new_n387_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n776_), .A2(new_n500_), .A3(new_n667_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT113), .Z(G1337gat));
  OAI21_X1  g582(.A(G99gat), .B1(new_n773_), .B2(new_n489_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n422_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n775_), .B2(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g587(.A1(new_n776_), .A2(new_n496_), .A3(new_n677_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n771_), .A2(new_n677_), .A3(new_n772_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(new_n791_), .A3(G106gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n790_), .B2(G106gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT53), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n789_), .B(new_n796_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1339gat));
  NOR2_X1   g597(.A1(new_n677_), .A2(new_n667_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n422_), .A2(new_n485_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(KEYINPUT59), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n589_), .A2(new_n547_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n539_), .A2(KEYINPUT116), .A3(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n530_), .B1(new_n534_), .B2(new_n538_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(G230gat), .A3(G233gat), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n804_), .B1(new_n539_), .B2(KEYINPUT116), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n546_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(KEYINPUT118), .A3(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(KEYINPUT56), .B(new_n546_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT118), .B1(new_n810_), .B2(new_n811_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n803_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n581_), .A2(new_n579_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n577_), .A2(new_n579_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n586_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n583_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n586_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n553_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n658_), .B1(new_n816_), .B2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n821_), .A2(new_n547_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n813_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n539_), .A2(KEYINPUT116), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT55), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n805_), .A3(new_n807_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT56), .B1(new_n828_), .B2(new_n546_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n824_), .B1(new_n825_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n631_), .A2(new_n634_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n830_), .A2(new_n831_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n823_), .A2(KEYINPUT57), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n810_), .A2(new_n811_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n840_), .A2(new_n803_), .B1(new_n553_), .B2(new_n821_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n836_), .B1(new_n841_), .B2(new_n658_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n648_), .B1(new_n834_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n588_), .A2(new_n648_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n846_), .A2(new_n555_), .A3(new_n590_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n847_), .A2(new_n688_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n847_), .B2(new_n688_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n802_), .B1(new_n843_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n823_), .B2(new_n835_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT120), .B(new_n836_), .C1(new_n841_), .C2(new_n658_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n834_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n851_), .B1(new_n856_), .B2(new_n649_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n801_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n589_), .B(new_n852_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G113gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n858_), .A2(new_n409_), .A3(new_n589_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1340gat));
  OAI211_X1 g662(.A(new_n745_), .B(new_n852_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G120gat), .ZN(new_n865_));
  INV_X1    g664(.A(new_n745_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n407_), .B1(new_n866_), .B2(KEYINPUT60), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n858_), .B(new_n867_), .C1(KEYINPUT60), .C2(new_n407_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n865_), .A2(new_n868_), .ZN(G1341gat));
  OAI211_X1 g668(.A(new_n648_), .B(new_n852_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G127gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n858_), .A2(new_n405_), .A3(new_n648_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1342gat));
  OAI211_X1 g672(.A(new_n635_), .B(new_n852_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(G134gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n858_), .A2(new_n403_), .A3(new_n658_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1343gat));
  XNOR2_X1  g676(.A(KEYINPUT121), .B(G141gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n856_), .A2(new_n649_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n851_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NOR4_X1   g680(.A1(new_n488_), .A2(new_n485_), .A3(new_n667_), .A4(new_n293_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n878_), .B1(new_n884_), .B2(new_n589_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n878_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n883_), .A2(new_n588_), .A3(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1344gat));
  NAND3_X1  g687(.A1(new_n881_), .A2(new_n745_), .A3(new_n882_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g689(.A1(new_n881_), .A2(new_n648_), .A3(new_n882_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT61), .B(G155gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1346gat));
  OR3_X1    g692(.A1(new_n883_), .A2(G162gat), .A3(new_n657_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G162gat), .B1(new_n883_), .B2(new_n688_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n843_), .A2(new_n851_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n488_), .A2(new_n485_), .A3(new_n667_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n897_), .A2(new_n677_), .A3(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n589_), .A3(new_n327_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n677_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n589_), .B(new_n901_), .C1(new_n843_), .C2(new_n851_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n902_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(G169gat), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n900_), .A2(new_n903_), .A3(new_n906_), .ZN(G1348gat));
  AOI21_X1  g706(.A(G176gat), .B1(new_n899_), .B2(new_n745_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n677_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n866_), .A2(new_n309_), .A3(new_n898_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(G1349gat));
  NOR2_X1   g710(.A1(new_n898_), .A2(new_n649_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G183gat), .B1(new_n909_), .B2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n318_), .A2(new_n319_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n648_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n901_), .B(new_n916_), .C1(new_n843_), .C2(new_n851_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  OAI21_X1  g717(.A(KEYINPUT122), .B1(new_n913_), .B2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920_));
  NOR4_X1   g719(.A1(new_n857_), .A2(new_n677_), .A3(new_n649_), .A4(new_n898_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n920_), .B(new_n917_), .C1(new_n921_), .C2(G183gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n919_), .A2(new_n922_), .ZN(G1350gat));
  NAND3_X1  g722(.A1(new_n899_), .A2(new_n344_), .A3(new_n658_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n635_), .B(new_n901_), .C1(new_n843_), .C2(new_n851_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(G190gat), .ZN(new_n927_));
  AND3_X1   g726(.A1(new_n926_), .A2(new_n925_), .A3(G190gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n924_), .B1(new_n927_), .B2(new_n928_), .ZN(G1351gat));
  NOR4_X1   g728(.A1(new_n488_), .A2(new_n452_), .A3(new_n387_), .A4(new_n293_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n881_), .A2(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(G197gat), .B1(new_n931_), .B2(new_n589_), .ZN(new_n932_));
  AND4_X1   g731(.A1(G197gat), .A2(new_n881_), .A3(new_n589_), .A4(new_n930_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1352gat));
  NAND3_X1  g733(.A1(new_n881_), .A2(new_n745_), .A3(new_n930_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n936_));
  XOR2_X1   g735(.A(new_n935_), .B(new_n936_), .Z(G1353gat));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n938_));
  AND3_X1   g737(.A1(new_n938_), .A2(new_n250_), .A3(KEYINPUT125), .ZN(new_n939_));
  AOI211_X1 g738(.A(new_n939_), .B(new_n649_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n881_), .A2(new_n930_), .A3(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(KEYINPUT125), .B1(new_n938_), .B2(new_n250_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n941_), .B(new_n942_), .ZN(G1354gat));
  NAND2_X1  g742(.A1(new_n931_), .A2(new_n658_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(KEYINPUT126), .B(G218gat), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n688_), .A2(new_n945_), .ZN(new_n946_));
  AOI22_X1  g745(.A1(new_n944_), .A2(new_n945_), .B1(new_n931_), .B2(new_n946_), .ZN(G1355gat));
endmodule


