//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n861_, new_n862_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR3_X1   g004(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  AND3_X1   g006(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT65), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n207_), .A2(new_n210_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(KEYINPUT8), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n217_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(G99gat), .ZN(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n228_), .A2(new_n213_), .A3(new_n215_), .A4(new_n204_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n222_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT8), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n210_), .A2(new_n216_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT9), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT64), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT9), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n220_), .A2(new_n235_), .A3(new_n237_), .A4(new_n221_), .ZN(new_n238_));
  OR2_X1    g037(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n227_), .A3(new_n240_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n234_), .A2(KEYINPUT64), .A3(G85gat), .A4(G92gat), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n238_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n224_), .A2(new_n232_), .B1(new_n233_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G64gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G57gat), .ZN(new_n246_));
  INV_X1    g045(.A(G57gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G64gat), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G71gat), .B(G78gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT11), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n249_), .A2(KEYINPUT11), .ZN(new_n252_));
  INV_X1    g051(.A(new_n250_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT11), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n251_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n244_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT66), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n244_), .A2(new_n256_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n203_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n224_), .A2(new_n232_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n243_), .A2(new_n233_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n256_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n261_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n244_), .A2(KEYINPUT12), .A3(new_n256_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n257_), .B(new_n202_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n260_), .A2(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G120gat), .B(G148gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(G176gat), .B(G204gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n274_), .B(KEYINPUT68), .Z(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n260_), .A2(new_n268_), .A3(new_n274_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT69), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n276_), .A2(new_n280_), .A3(new_n277_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n279_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT13), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n279_), .A2(new_n281_), .A3(new_n282_), .A4(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT80), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G113gat), .B(G141gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G169gat), .B(G197gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G1gat), .ZN(new_n295_));
  INV_X1    g094(.A(G8gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT14), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(G22gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G15gat), .ZN(new_n299_));
  INV_X1    g098(.A(G15gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G22gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n297_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT77), .ZN(new_n303_));
  XOR2_X1   g102(.A(G1gat), .B(G8gat), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n303_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G29gat), .B(G36gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G43gat), .B(G50gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n303_), .B(new_n304_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n309_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G229gat), .A2(G233gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n309_), .B(KEYINPUT15), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n311_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n310_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n294_), .B1(new_n316_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n316_), .A2(new_n320_), .A3(new_n294_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n290_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n323_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(new_n321_), .A3(KEYINPUT80), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT2), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n331_), .A2(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n332_), .B2(new_n331_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT88), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n328_), .B(new_n330_), .C1(new_n336_), .C2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n329_), .B1(KEYINPUT1), .B2(new_n328_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(KEYINPUT1), .B2(new_n328_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n331_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n333_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n344_), .A2(KEYINPUT29), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT28), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G228gat), .ZN(new_n348_));
  INV_X1    g147(.A(G233gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G211gat), .B(G218gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT89), .ZN(new_n353_));
  INV_X1    g152(.A(G197gat), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n354_), .A2(G204gat), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n352_), .B(KEYINPUT21), .C1(new_n353_), .C2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G197gat), .B(G204gat), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n357_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n352_), .A2(KEYINPUT21), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT90), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n344_), .A2(KEYINPUT29), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n351_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G78gat), .B(G106gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n366_), .B(KEYINPUT91), .Z(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n361_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n364_), .A2(new_n369_), .A3(new_n351_), .ZN(new_n370_));
  OR3_X1    g169(.A1(new_n365_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n368_), .B1(new_n365_), .B2(new_n370_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G22gat), .B(G50gat), .Z(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n347_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(new_n346_), .A3(new_n374_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT23), .ZN(new_n383_));
  OR3_X1    g182(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n383_), .B1(new_n386_), .B2(KEYINPUT24), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT23), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n382_), .B(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT24), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n384_), .A2(new_n385_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT82), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT24), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT25), .B(G183gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT26), .B(G190gat), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n386_), .A2(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n389_), .A2(new_n395_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n396_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT22), .B(G169gat), .ZN(new_n404_));
  INV_X1    g203(.A(G176gat), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n406_), .A2(KEYINPUT83), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n383_), .B1(G183gat), .B2(G190gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(KEYINPUT83), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n402_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT84), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n402_), .A2(KEYINPUT84), .A3(new_n410_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n369_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT20), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n400_), .B(KEYINPUT92), .Z(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n399_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n387_), .A2(KEYINPUT94), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT94), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n394_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n397_), .B(KEYINPUT93), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n386_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n419_), .A2(new_n420_), .A3(new_n422_), .A4(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n408_), .A2(new_n406_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n417_), .B1(new_n427_), .B2(new_n361_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n416_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G226gat), .A2(G233gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT19), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n369_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n425_), .A2(new_n369_), .A3(new_n426_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT20), .B(new_n431_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT18), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G64gat), .B(G92gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT20), .B1(new_n434_), .B2(new_n435_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n443_), .A2(new_n431_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n363_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n417_), .B1(new_n445_), .B2(new_n427_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n432_), .B1(new_n446_), .B2(new_n416_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n442_), .B(KEYINPUT27), .C1(new_n441_), .C2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G127gat), .B(G134gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(G113gat), .B(G120gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n344_), .B(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G225gat), .A2(G233gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n344_), .A2(new_n457_), .A3(new_n452_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n455_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n456_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G1gat), .B(G29gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(G57gat), .B(G85gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n464_), .B(new_n465_), .Z(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n456_), .B(new_n468_), .C1(new_n458_), .C2(new_n460_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT27), .ZN(new_n472_));
  INV_X1    g271(.A(new_n441_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n433_), .A2(new_n473_), .A3(new_n436_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n473_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n472_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n449_), .A2(new_n471_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n381_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G71gat), .B(G99gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT85), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n480_), .B(G43gat), .Z(new_n481_));
  NAND2_X1  g280(.A1(G227gat), .A2(G233gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(new_n300_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n481_), .B(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n413_), .A2(KEYINPUT30), .A3(new_n414_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT30), .B1(new_n413_), .B2(new_n414_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n485_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n488_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(new_n486_), .A3(new_n484_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT86), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n489_), .A2(new_n491_), .A3(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n452_), .B(KEYINPUT31), .Z(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n489_), .A2(new_n491_), .A3(new_n494_), .A4(new_n496_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n474_), .A2(new_n475_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT96), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n505_), .A2(KEYINPUT33), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n469_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n469_), .A2(new_n506_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n459_), .A2(new_n454_), .ZN(new_n509_));
  OAI221_X1 g308(.A(new_n466_), .B1(new_n453_), .B2(new_n454_), .C1(new_n458_), .C2(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n504_), .A2(new_n507_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n441_), .A2(KEYINPUT32), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n437_), .A2(new_n513_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n514_), .B(new_n470_), .C1(new_n448_), .C2(new_n513_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n380_), .A2(new_n512_), .A3(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n478_), .A2(new_n503_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n498_), .A2(new_n500_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n518_), .A2(new_n470_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n449_), .A2(KEYINPUT97), .A3(new_n476_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT97), .B1(new_n449_), .B2(new_n476_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n380_), .B(new_n519_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n522_));
  AOI211_X1 g321(.A(new_n289_), .B(new_n327_), .C1(new_n517_), .C2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G232gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(KEYINPUT35), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n527_), .B1(new_n244_), .B2(new_n309_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n528_), .A2(KEYINPUT72), .B1(new_n264_), .B2(new_n318_), .ZN(new_n529_));
  OAI22_X1  g328(.A1(new_n264_), .A2(new_n312_), .B1(KEYINPUT35), .B2(new_n526_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT72), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n526_), .A2(KEYINPUT35), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT75), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n318_), .A2(new_n264_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(new_n528_), .A3(new_n534_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT74), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT74), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n538_), .A2(new_n528_), .A3(new_n541_), .A4(new_n534_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n536_), .A2(new_n537_), .A3(new_n540_), .A4(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n542_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n534_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT75), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G190gat), .B(G218gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT73), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G134gat), .B(G162gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT36), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n543_), .A2(new_n546_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT37), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n550_), .A2(new_n551_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n536_), .A2(new_n556_), .A3(new_n540_), .A4(new_n542_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT76), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n553_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT37), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n558_), .A2(new_n559_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n559_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G127gat), .B(G155gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT16), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G183gat), .B(G211gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n256_), .B(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n311_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n311_), .A2(new_n572_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n570_), .B1(new_n575_), .B2(KEYINPUT78), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n573_), .A2(new_n574_), .A3(new_n569_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT79), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(KEYINPUT17), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n578_), .B1(new_n577_), .B2(KEYINPUT17), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n576_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n581_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n576_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n584_), .A3(new_n579_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n565_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n523_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT98), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n295_), .A3(new_n470_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT38), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n517_), .A2(new_n522_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n554_), .A2(new_n557_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT99), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596_));
  INV_X1    g395(.A(new_n594_), .ZN(new_n597_));
  AOI211_X1 g396(.A(new_n596_), .B(new_n597_), .C1(new_n517_), .C2(new_n522_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n289_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n322_), .A2(new_n323_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(new_n587_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G1gat), .B1(new_n605_), .B2(new_n471_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n592_), .A2(new_n606_), .ZN(G1324gat));
  INV_X1    g406(.A(new_n520_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n521_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n611_), .B(new_n604_), .C1(new_n595_), .C2(new_n598_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT100), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G8gat), .B1(new_n612_), .B2(new_n613_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT39), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n612_), .A2(new_n613_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n618_), .A2(new_n619_), .A3(G8gat), .A4(new_n614_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n590_), .A2(new_n296_), .A3(new_n611_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n621_), .A2(KEYINPUT40), .A3(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1325gat));
  OAI21_X1  g426(.A(G15gat), .B1(new_n605_), .B2(new_n503_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n628_), .A2(KEYINPUT41), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(KEYINPUT41), .ZN(new_n630_));
  INV_X1    g429(.A(new_n503_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n590_), .A2(new_n300_), .A3(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n629_), .A2(new_n630_), .A3(new_n632_), .ZN(G1326gat));
  NAND3_X1  g432(.A1(new_n590_), .A2(new_n298_), .A3(new_n381_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G22gat), .B1(new_n605_), .B2(new_n380_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(KEYINPUT42), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(KEYINPUT42), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n634_), .B1(new_n636_), .B2(new_n637_), .ZN(G1327gat));
  NOR2_X1   g437(.A1(new_n586_), .A2(new_n594_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n523_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(G29gat), .B1(new_n640_), .B2(new_n470_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n603_), .A2(new_n586_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n593_), .B2(new_n565_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n565_), .ZN(new_n645_));
  AOI211_X1 g444(.A(KEYINPUT43), .B(new_n645_), .C1(new_n517_), .C2(new_n522_), .ZN(new_n646_));
  OAI211_X1 g445(.A(KEYINPUT44), .B(new_n642_), .C1(new_n644_), .C2(new_n646_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n647_), .A2(G29gat), .A3(new_n470_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n642_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n641_), .B1(new_n648_), .B2(new_n651_), .ZN(G1328gat));
  INV_X1    g451(.A(G36gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n640_), .A2(new_n653_), .A3(new_n611_), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT46), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n651_), .A2(new_n611_), .A3(new_n647_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(KEYINPUT101), .A3(G36gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT101), .B1(new_n660_), .B2(G36gat), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n656_), .B(new_n659_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n655_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n654_), .B(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n660_), .A2(G36gat), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n660_), .A2(KEYINPUT101), .A3(G36gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT103), .B1(new_n658_), .B2(KEYINPUT46), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n658_), .B2(KEYINPUT46), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n663_), .B1(new_n670_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(G1329gat));
  INV_X1    g473(.A(new_n518_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n651_), .A2(G43gat), .A3(new_n675_), .A4(new_n647_), .ZN(new_n676_));
  XOR2_X1   g475(.A(KEYINPUT105), .B(G43gat), .Z(new_n677_));
  INV_X1    g476(.A(new_n640_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(new_n678_), .B2(new_n503_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g480(.A1(new_n678_), .A2(G50gat), .A3(new_n380_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n651_), .A2(new_n381_), .A3(new_n647_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(new_n684_), .A3(G50gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n683_), .B2(G50gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(G1331gat));
  NAND2_X1  g486(.A1(new_n324_), .A2(new_n326_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n600_), .A2(new_n587_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n599_), .A2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G57gat), .B1(new_n690_), .B2(new_n471_), .ZN(new_n691_));
  AOI211_X1 g490(.A(new_n602_), .B(new_n600_), .C1(new_n517_), .C2(new_n522_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n588_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(new_n247_), .A3(new_n470_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n691_), .A2(new_n695_), .ZN(G1332gat));
  OAI21_X1  g495(.A(G64gat), .B1(new_n690_), .B2(new_n610_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT48), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n694_), .A2(new_n245_), .A3(new_n611_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1333gat));
  OAI21_X1  g499(.A(G71gat), .B1(new_n690_), .B2(new_n503_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT49), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n503_), .A2(G71gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n693_), .B2(new_n703_), .ZN(G1334gat));
  OAI21_X1  g503(.A(G78gat), .B1(new_n690_), .B2(new_n380_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT50), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n380_), .A2(G78gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n693_), .B2(new_n707_), .ZN(G1335gat));
  AND2_X1   g507(.A1(new_n692_), .A2(new_n639_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(new_n218_), .A3(new_n470_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n644_), .A2(new_n646_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n600_), .A2(new_n602_), .A3(new_n586_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n470_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n710_), .B1(new_n715_), .B2(new_n218_), .ZN(G1336gat));
  NAND3_X1  g515(.A1(new_n709_), .A2(new_n219_), .A3(new_n611_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n713_), .A2(new_n611_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n719_), .B2(new_n219_), .ZN(G1337gat));
  AOI21_X1  g519(.A(new_n226_), .B1(new_n713_), .B2(new_n631_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n675_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n709_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(KEYINPUT107), .A2(KEYINPUT51), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(G1338gat));
  NAND3_X1  g524(.A1(new_n709_), .A2(new_n227_), .A3(new_n381_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n711_), .A2(new_n381_), .A3(new_n712_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(G106gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G106gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g531(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT108), .B1(new_n587_), .B2(new_n688_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n327_), .A2(new_n735_), .A3(new_n586_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n733_), .B1(new_n738_), .B2(new_n565_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n733_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n600_), .A2(new_n645_), .A3(new_n737_), .A4(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT57), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n744_));
  INV_X1    g543(.A(new_n275_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n262_), .A2(new_n263_), .A3(new_n256_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT12), .B1(new_n244_), .B2(new_n256_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n263_), .ZN(new_n748_));
  AOI22_X1  g547(.A1(new_n217_), .A2(new_n223_), .B1(new_n231_), .B2(KEYINPUT8), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n261_), .B(new_n265_), .C1(new_n748_), .C2(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n746_), .B1(new_n747_), .B2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT55), .B1(new_n751_), .B2(new_n202_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n202_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(KEYINPUT55), .A3(new_n202_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n745_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n744_), .B1(new_n756_), .B2(KEYINPUT56), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n268_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n257_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n203_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n759_), .A2(new_n755_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n275_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(KEYINPUT110), .A3(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(KEYINPUT56), .A3(new_n275_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n762_), .A2(KEYINPUT111), .A3(KEYINPUT56), .A4(new_n275_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n757_), .A2(new_n765_), .A3(new_n768_), .A4(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n277_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n601_), .A2(new_n771_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n770_), .A2(KEYINPUT112), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT112), .B1(new_n770_), .B2(new_n772_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n310_), .A2(new_n319_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n775_), .B(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(new_n315_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n314_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n293_), .B1(new_n779_), .B2(new_n317_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n321_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n773_), .A2(new_n774_), .A3(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n743_), .B1(new_n783_), .B2(new_n597_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n770_), .A2(new_n772_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n770_), .A2(KEYINPUT112), .A3(new_n772_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(KEYINPUT57), .A3(new_n594_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n756_), .A2(KEYINPUT114), .A3(KEYINPUT56), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n766_), .A2(new_n792_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n791_), .A2(new_n793_), .B1(new_n764_), .B2(new_n763_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n781_), .A2(new_n771_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(KEYINPUT58), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n781_), .A2(new_n771_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n794_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n565_), .A2(new_n797_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n784_), .A2(new_n790_), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n742_), .B1(new_n803_), .B2(new_n587_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n518_), .A2(new_n471_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n610_), .A2(new_n380_), .A3(new_n805_), .ZN(new_n806_));
  OR3_X1    g605(.A1(new_n804_), .A2(KEYINPUT115), .A3(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT115), .B1(new_n804_), .B2(new_n806_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n602_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810_));
  INV_X1    g609(.A(G113gat), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n806_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n597_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n801_), .B1(new_n817_), .B2(KEYINPUT57), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n586_), .B1(new_n818_), .B2(new_n784_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT59), .B(new_n816_), .C1(new_n819_), .C2(new_n742_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n815_), .A2(new_n821_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n822_), .A2(new_n811_), .A3(new_n327_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n810_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n812_), .A2(new_n823_), .A3(new_n824_), .ZN(G1340gat));
  INV_X1    g624(.A(KEYINPUT60), .ZN(new_n826_));
  INV_X1    g625(.A(G120gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n289_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n807_), .A2(new_n808_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n600_), .B1(new_n814_), .B2(new_n820_), .ZN(new_n831_));
  OAI21_X1  g630(.A(G120gat), .B1(new_n831_), .B2(KEYINPUT117), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833_));
  AOI211_X1 g632(.A(new_n833_), .B(new_n600_), .C1(new_n814_), .C2(new_n820_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n830_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT118), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n837_), .B(new_n830_), .C1(new_n832_), .C2(new_n834_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1341gat));
  OAI21_X1  g638(.A(G127gat), .B1(new_n822_), .B2(new_n587_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n587_), .A2(G127gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n807_), .A2(new_n808_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1342gat));
  NAND3_X1  g642(.A1(new_n807_), .A2(new_n597_), .A3(new_n808_), .ZN(new_n844_));
  INV_X1    g643(.A(G134gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT119), .B(G134gat), .Z(new_n847_));
  OAI211_X1 g646(.A(new_n565_), .B(new_n847_), .C1(new_n815_), .C2(new_n821_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT120), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n846_), .A2(new_n851_), .A3(new_n848_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1343gat));
  INV_X1    g652(.A(new_n804_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n631_), .A2(new_n380_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n854_), .A2(new_n470_), .A3(new_n610_), .A4(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n601_), .ZN(new_n857_));
  XOR2_X1   g656(.A(new_n857_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g657(.A1(new_n856_), .A2(new_n600_), .ZN(new_n859_));
  XOR2_X1   g658(.A(new_n859_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g659(.A1(new_n856_), .A2(new_n587_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT61), .B(G155gat), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n861_), .B(new_n862_), .Z(G1346gat));
  OAI21_X1  g662(.A(G162gat), .B1(new_n856_), .B2(new_n645_), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n594_), .A2(G162gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n856_), .B2(new_n865_), .ZN(G1347gat));
  NOR4_X1   g665(.A1(new_n610_), .A2(new_n470_), .A3(new_n381_), .A4(new_n503_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n854_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n602_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n404_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n870_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT62), .B1(new_n870_), .B2(G169gat), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1348gat));
  NAND2_X1  g674(.A1(KEYINPUT121), .A2(G176gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n868_), .B2(new_n600_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT122), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n879_), .B(new_n876_), .C1(new_n868_), .C2(new_n600_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(new_n881_));
  OR2_X1    g680(.A1(KEYINPUT121), .A2(G176gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1349gat));
  NAND2_X1  g682(.A1(new_n869_), .A2(new_n586_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(KEYINPUT123), .B2(G183gat), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n399_), .B1(new_n886_), .B2(G183gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n885_), .B1(new_n884_), .B2(new_n887_), .ZN(G1350gat));
  OAI21_X1  g687(.A(G190gat), .B1(new_n868_), .B2(new_n645_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n597_), .A2(new_n418_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n868_), .B2(new_n890_), .ZN(G1351gat));
  NOR2_X1   g690(.A1(new_n610_), .A2(new_n470_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n855_), .B(new_n892_), .C1(new_n819_), .C2(new_n742_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n894_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  OAI211_X1 g696(.A(KEYINPUT125), .B(new_n354_), .C1(new_n897_), .C2(new_n601_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n601_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(G197gat), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(G197gat), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n898_), .A2(new_n901_), .A3(new_n902_), .ZN(G1352gat));
  NAND2_X1  g702(.A1(new_n895_), .A2(new_n896_), .ZN(new_n904_));
  AND4_X1   g703(.A1(KEYINPUT126), .A2(new_n904_), .A3(G204gat), .A4(new_n289_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT126), .B(G204gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n906_), .B1(new_n904_), .B2(new_n289_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1353gat));
  AOI21_X1  g707(.A(new_n587_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n904_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT127), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n910_), .B(new_n912_), .ZN(G1354gat));
  OR3_X1    g712(.A1(new_n897_), .A2(G218gat), .A3(new_n594_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G218gat), .B1(new_n897_), .B2(new_n645_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1355gat));
endmodule


