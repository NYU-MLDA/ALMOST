//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n878_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT76), .B(G15gat), .ZN(new_n205_));
  INV_X1    g004(.A(G22gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G1gat), .ZN(new_n208_));
  INV_X1    g007(.A(G8gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G1gat), .B(G8gat), .Z(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G29gat), .B(G36gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(KEYINPUT15), .ZN(new_n218_));
  INV_X1    g017(.A(new_n213_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n213_), .B(new_n216_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n221_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n204_), .B1(new_n222_), .B2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n226_), .B(KEYINPUT81), .Z(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(new_n225_), .A3(new_n204_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT82), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n229_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT6), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n235_), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G99gat), .A2(G106gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(KEYINPUT6), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n234_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(KEYINPUT6), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n235_), .A2(G99gat), .A3(G106gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT66), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR3_X1   g043(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(new_n242_), .A3(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(G85gat), .A2(G92gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G85gat), .A2(G92gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(KEYINPUT8), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT67), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n247_), .A2(new_n254_), .A3(new_n251_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n244_), .A2(new_n245_), .A3(new_n256_), .ZN(new_n257_));
  OR3_X1    g056(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT69), .B1(new_n258_), .B2(new_n243_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT68), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT68), .B1(new_n240_), .B2(new_n241_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n250_), .B1(new_n260_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT8), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n253_), .B(new_n255_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT66), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT66), .B1(new_n240_), .B2(new_n241_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT10), .B(G99gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G106gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT9), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n248_), .B1(new_n276_), .B2(new_n249_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT64), .B(G92gat), .ZN(new_n278_));
  INV_X1    g077(.A(G85gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n276_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n277_), .B1(new_n281_), .B2(KEYINPUT65), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n275_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n267_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n218_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n247_), .A2(new_n254_), .A3(new_n251_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n254_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n258_), .A2(new_n243_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n256_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n263_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n258_), .A2(KEYINPUT69), .A3(new_n243_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n261_), .A4(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n250_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT8), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n285_), .B1(new_n291_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n216_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G232gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT34), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n288_), .B(new_n301_), .C1(KEYINPUT35), .C2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(KEYINPUT35), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G190gat), .B(G218gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G134gat), .B(G162gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n309_), .B(KEYINPUT36), .Z(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT75), .B1(new_n306_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT37), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n309_), .A2(KEYINPUT36), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n306_), .A2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(new_n306_), .B2(new_n311_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n313_), .B(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G231gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n213_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G57gat), .B(G64gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT11), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n322_));
  INV_X1    g121(.A(G64gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G57gat), .ZN(new_n324_));
  INV_X1    g123(.A(G57gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(G64gat), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT11), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G71gat), .B(G78gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n322_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n330_));
  AND2_X1   g129(.A1(G71gat), .A2(G78gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G71gat), .A2(G78gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n333_), .B(KEYINPUT70), .C1(new_n320_), .C2(KEYINPUT11), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n329_), .A2(new_n330_), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n330_), .B1(new_n329_), .B2(new_n334_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n321_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n324_), .A2(new_n326_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT11), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT70), .B1(new_n340_), .B2(new_n333_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n327_), .A2(new_n322_), .A3(new_n328_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT71), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n321_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n329_), .A2(new_n330_), .A3(new_n334_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n337_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n319_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT17), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G183gat), .B(G211gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT78), .ZN(new_n352_));
  XOR2_X1   g151(.A(G127gat), .B(G155gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n349_), .A2(new_n350_), .A3(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT79), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n356_), .B(KEYINPUT17), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n349_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n317_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G230gat), .A2(G233gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI211_X1 g163(.A(KEYINPUT73), .B(new_n364_), .C1(new_n300_), .C2(new_n347_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT73), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n347_), .A2(new_n267_), .A3(new_n286_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n367_), .B2(new_n363_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT72), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT12), .ZN(new_n371_));
  OAI22_X1  g170(.A1(new_n300_), .A2(new_n347_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n337_), .A2(new_n346_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n287_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT74), .B1(new_n369_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n367_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n300_), .A2(new_n347_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n364_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n372_), .A2(new_n375_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT74), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n381_), .B(new_n382_), .C1(new_n368_), .C2(new_n365_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n377_), .A2(new_n380_), .A3(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G120gat), .B(G148gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT5), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G176gat), .B(G204gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  OR2_X1    g187(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n384_), .A2(new_n388_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n389_), .A2(KEYINPUT13), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT13), .B1(new_n389_), .B2(new_n390_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n362_), .A2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n233_), .B1(new_n394_), .B2(KEYINPUT80), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT24), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G169gat), .A2(G176gat), .ZN(new_n398_));
  MUX2_X1   g197(.A(new_n397_), .B(KEYINPUT24), .S(new_n398_), .Z(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT26), .B(G190gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401_));
  INV_X1    g200(.A(G183gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT25), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n402_), .A2(KEYINPUT25), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n400_), .B(new_n403_), .C1(new_n404_), .C2(new_n401_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G183gat), .A2(G190gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT84), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT23), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n406_), .ZN(new_n410_));
  OAI22_X1  g209(.A1(new_n409_), .A2(KEYINPUT85), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n409_), .A2(KEYINPUT85), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n399_), .B(new_n405_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT22), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(KEYINPUT86), .A3(G169gat), .ZN(new_n415_));
  INV_X1    g214(.A(G176gat), .ZN(new_n416_));
  AND2_X1   g215(.A1(KEYINPUT86), .A2(G169gat), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n415_), .B(new_n416_), .C1(new_n414_), .C2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n407_), .A2(KEYINPUT23), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n419_), .B1(KEYINPUT23), .B2(new_n410_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G183gat), .A2(G190gat), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n396_), .B(new_n418_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n413_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G15gat), .B(G43gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT89), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n423_), .B(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(KEYINPUT87), .B(KEYINPUT30), .Z(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G227gat), .A2(G233gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT88), .ZN(new_n430_));
  INV_X1    g229(.A(G71gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n428_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G127gat), .B(G134gat), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n434_), .A2(KEYINPUT90), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(KEYINPUT90), .ZN(new_n436_));
  XOR2_X1   g235(.A(G113gat), .B(G120gat), .Z(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT91), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n435_), .A2(new_n436_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n437_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n440_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT31), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(G99gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n433_), .B(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(G1gat), .B(G29gat), .Z(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT104), .B(KEYINPUT0), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G57gat), .B(G85gat), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n451_), .B(new_n452_), .Z(new_n453_));
  NAND2_X1  g252(.A1(G225gat), .A2(G233gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G155gat), .A2(G162gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT92), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT1), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT93), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n457_), .A2(KEYINPUT93), .A3(new_n458_), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n456_), .B(KEYINPUT92), .Z(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT1), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G155gat), .A2(G162gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n461_), .A2(new_n462_), .A3(new_n464_), .A4(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G141gat), .A2(G148gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(G141gat), .A2(G148gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n467_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n470_), .B(KEYINPUT3), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n468_), .B(KEYINPUT2), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n457_), .A2(new_n465_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n472_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n444_), .A2(new_n478_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n467_), .A2(new_n471_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n443_), .A2(new_n438_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n455_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT4), .B1(new_n444_), .B2(new_n478_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n482_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n485_), .B2(KEYINPUT4), .ZN(new_n486_));
  AOI211_X1 g285(.A(new_n453_), .B(new_n483_), .C1(new_n486_), .C2(new_n455_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n453_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(KEYINPUT4), .ZN(new_n489_));
  INV_X1    g288(.A(new_n484_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n455_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n483_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n488_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n487_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n448_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT25), .B(G183gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n400_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n399_), .A2(new_n498_), .ZN(new_n499_));
  OR3_X1    g298(.A1(new_n420_), .A2(new_n499_), .A3(KEYINPUT101), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT101), .B1(new_n420_), .B2(new_n499_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT103), .ZN(new_n503_));
  INV_X1    g302(.A(G204gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(G197gat), .ZN(new_n505_));
  INV_X1    g304(.A(G197gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n506_), .A2(G204gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT21), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G211gat), .B(G218gat), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n507_), .B1(KEYINPUT96), .B2(new_n505_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(KEYINPUT96), .B2(new_n505_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n508_), .B(new_n509_), .C1(new_n511_), .C2(KEYINPUT21), .ZN(new_n512_));
  INV_X1    g311(.A(new_n509_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(KEYINPUT21), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n421_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT22), .B(G169gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n416_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n396_), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n521_), .B(KEYINPUT102), .Z(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n502_), .A2(new_n503_), .A3(new_n516_), .A4(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G226gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT20), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AND4_X1   g328(.A1(new_n516_), .A2(new_n523_), .A3(new_n501_), .A4(new_n500_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT103), .B1(new_n423_), .B2(new_n515_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n524_), .B(new_n529_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n527_), .B(KEYINPUT100), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n516_), .B1(new_n502_), .B2(new_n523_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT20), .B1(new_n423_), .B2(new_n515_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n534_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G8gat), .B(G36gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT18), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G64gat), .B(G92gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  NAND3_X1  g340(.A1(new_n532_), .A2(new_n537_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT106), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n541_), .B(KEYINPUT105), .Z(new_n544_));
  NOR3_X1   g343(.A1(new_n535_), .A2(new_n536_), .A3(new_n534_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n527_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n528_), .B1(new_n423_), .B2(new_n515_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n523_), .B(new_n516_), .C1(new_n420_), .C2(new_n499_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n544_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT106), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n532_), .A2(new_n537_), .A3(new_n551_), .A4(new_n541_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n543_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT27), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n532_), .A2(new_n537_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n541_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT27), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(new_n542_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G22gat), .B(G50gat), .Z(new_n561_));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT29), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n480_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n562_), .B1(new_n480_), .B2(new_n563_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n564_), .A2(new_n565_), .A3(KEYINPUT94), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT28), .B1(new_n478_), .B2(KEYINPUT29), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n480_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n561_), .B1(new_n566_), .B2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT94), .B1(new_n564_), .B2(new_n565_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n568_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n561_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G78gat), .B(G106gat), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n577_), .A2(KEYINPUT97), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n571_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n576_), .B1(new_n571_), .B2(new_n575_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n516_), .B1(new_n478_), .B2(KEYINPUT29), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT95), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n579_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n574_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n577_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n571_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n584_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G228gat), .A2(G233gat), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT98), .Z(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n583_), .A2(new_n589_), .A3(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n582_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n587_), .A2(new_n588_), .A3(new_n584_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n591_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n496_), .A2(new_n560_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT107), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n493_), .A2(KEYINPUT33), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT33), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n483_), .B1(new_n486_), .B2(new_n455_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n602_), .B1(new_n603_), .B2(new_n488_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n486_), .A2(new_n455_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n488_), .B1(new_n485_), .B2(new_n454_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n557_), .B(new_n542_), .C1(new_n606_), .C2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n541_), .A2(KEYINPUT32), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n609_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n610_), .B1(new_n555_), .B2(new_n609_), .ZN(new_n611_));
  OAI22_X1  g410(.A1(new_n605_), .A2(new_n608_), .B1(new_n494_), .B2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n593_), .B2(new_n596_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n592_), .B1(new_n583_), .B2(new_n589_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n594_), .A2(new_n591_), .A3(new_n595_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n614_), .A2(new_n560_), .A3(new_n615_), .A4(new_n494_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n600_), .B1(new_n617_), .B2(new_n448_), .ZN(new_n618_));
  AOI211_X1 g417(.A(KEYINPUT107), .B(new_n447_), .C1(new_n613_), .C2(new_n616_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n599_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI211_X1 g420(.A(new_n395_), .B(new_n621_), .C1(KEYINPUT80), .C2(new_n394_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n208_), .A3(new_n495_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT38), .ZN(new_n624_));
  INV_X1    g423(.A(new_n393_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n233_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n620_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n316_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n361_), .A2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n631_), .A2(new_n495_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n624_), .B1(new_n208_), .B2(new_n632_), .ZN(G1324gat));
  INV_X1    g432(.A(new_n560_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n209_), .B1(new_n631_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n622_), .A2(new_n209_), .A3(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(G1325gat));
  INV_X1    g440(.A(G15gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n631_), .B2(new_n447_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT41), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n622_), .A2(new_n642_), .A3(new_n447_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1326gat));
  AOI21_X1  g445(.A(new_n206_), .B1(new_n631_), .B2(new_n597_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT42), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n622_), .A2(new_n597_), .A3(new_n206_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1327gat));
  INV_X1    g449(.A(new_n361_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n316_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n628_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n495_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n625_), .A2(new_n651_), .A3(new_n626_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n620_), .A2(new_n656_), .A3(new_n317_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n620_), .B2(new_n317_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n655_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(KEYINPUT44), .B(new_n655_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n495_), .A2(G29gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n654_), .B1(new_n663_), .B2(new_n664_), .ZN(G1328gat));
  XNOR2_X1  g464(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(new_n634_), .A3(new_n662_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G36gat), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT108), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT108), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n667_), .A2(new_n670_), .A3(G36gat), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT109), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n560_), .A2(G36gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n653_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n628_), .A2(new_n652_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n674_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT109), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n675_), .A2(KEYINPUT45), .A3(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT45), .B1(new_n675_), .B2(new_n678_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n666_), .B1(new_n672_), .B2(new_n681_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n667_), .A2(new_n670_), .A3(G36gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n670_), .B1(new_n667_), .B2(G36gat), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n681_), .B(new_n666_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n682_), .A2(new_n686_), .ZN(G1329gat));
  NAND3_X1  g486(.A1(new_n663_), .A2(G43gat), .A3(new_n447_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n676_), .A2(new_n448_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(G43gat), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g490(.A1(new_n663_), .A2(new_n597_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G50gat), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n598_), .A2(G50gat), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT111), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n676_), .B2(new_n695_), .ZN(G1331gat));
  NOR2_X1   g495(.A1(new_n393_), .A2(new_n233_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n620_), .A2(new_n697_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(new_n630_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G57gat), .B1(new_n700_), .B2(new_n494_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n698_), .A2(new_n362_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n325_), .A3(new_n495_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1332gat));
  AOI21_X1  g503(.A(new_n323_), .B1(new_n699_), .B2(new_n634_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT48), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n702_), .A2(new_n323_), .A3(new_n634_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1333gat));
  AOI21_X1  g507(.A(new_n431_), .B1(new_n699_), .B2(new_n447_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n702_), .A2(new_n431_), .A3(new_n447_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1334gat));
  INV_X1    g512(.A(G78gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n699_), .B2(new_n597_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT50), .Z(new_n716_));
  NAND3_X1  g515(.A1(new_n702_), .A2(new_n714_), .A3(new_n597_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1335gat));
  NOR2_X1   g517(.A1(new_n657_), .A2(new_n658_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n697_), .A2(new_n361_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n279_), .B1(new_n721_), .B2(new_n495_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n698_), .A2(new_n652_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n723_), .A2(new_n279_), .A3(new_n495_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1336gat));
  AOI21_X1  g524(.A(G92gat), .B1(new_n723_), .B2(new_n634_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n560_), .A2(new_n278_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n721_), .B2(new_n727_), .ZN(G1337gat));
  INV_X1    g527(.A(new_n720_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n447_), .B(new_n729_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G99gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n723_), .A2(new_n272_), .A3(new_n447_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(KEYINPUT114), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n731_), .A2(new_n732_), .A3(KEYINPUT113), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(KEYINPUT51), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT115), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT51), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n733_), .A2(new_n734_), .A3(new_n739_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n737_), .A2(new_n738_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n738_), .B1(new_n737_), .B2(new_n740_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1338gat));
  NAND2_X1  g542(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G106gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n721_), .B2(new_n597_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n746_), .A2(new_n748_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n723_), .A2(new_n273_), .A3(new_n597_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n749_), .A2(new_n750_), .A3(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g554(.A1(new_n394_), .A2(new_n233_), .ZN(new_n756_));
  XOR2_X1   g555(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n757_));
  XNOR2_X1  g556(.A(new_n756_), .B(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n233_), .A2(new_n389_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n377_), .A2(new_n761_), .A3(new_n383_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n368_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n367_), .A2(new_n366_), .A3(new_n363_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n376_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n372_), .A2(new_n367_), .A3(new_n375_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n765_), .A2(KEYINPUT55), .B1(new_n364_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n762_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT119), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT119), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n762_), .A2(new_n767_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT56), .B1(new_n772_), .B2(new_n388_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n762_), .A2(new_n770_), .A3(new_n767_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n770_), .B1(new_n762_), .B2(new_n767_), .ZN(new_n775_));
  OAI211_X1 g574(.A(KEYINPUT56), .B(new_n388_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n760_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n389_), .A2(new_n390_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n220_), .A2(new_n224_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n204_), .B1(new_n223_), .B2(new_n221_), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n230_), .A2(new_n231_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n629_), .B1(new_n778_), .B2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT57), .B1(new_n784_), .B2(KEYINPUT120), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n388_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n759_), .B1(new_n788_), .B2(new_n776_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n783_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n316_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT57), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n389_), .A2(new_n782_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT121), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n389_), .A2(new_n782_), .A3(KEYINPUT121), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT122), .B1(new_n802_), .B2(new_n317_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n788_), .A2(new_n776_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT122), .B(new_n317_), .C1(new_n804_), .C2(KEYINPUT58), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(KEYINPUT58), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n785_), .B(new_n794_), .C1(new_n803_), .C2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n758_), .B1(new_n808_), .B2(new_n361_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NOR4_X1   g609(.A1(new_n448_), .A2(new_n597_), .A3(new_n494_), .A4(new_n634_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(G113gat), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n233_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(KEYINPUT123), .A3(KEYINPUT59), .ZN(new_n816_));
  OR2_X1    g615(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n817_));
  NAND2_X1  g616(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n812_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n626_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n815_), .B1(new_n820_), .B2(new_n814_), .ZN(G1340gat));
  INV_X1    g620(.A(G120gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n393_), .B2(KEYINPUT60), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n813_), .B(new_n823_), .C1(KEYINPUT60), .C2(new_n822_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n393_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n822_), .ZN(G1341gat));
  AOI21_X1  g625(.A(G127gat), .B1(new_n813_), .B2(new_n651_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n816_), .A2(new_n819_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n651_), .A2(G127gat), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT124), .Z(new_n830_));
  AOI21_X1  g629(.A(new_n827_), .B1(new_n828_), .B2(new_n830_), .ZN(G1342gat));
  INV_X1    g630(.A(G134gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n813_), .A2(new_n832_), .A3(new_n629_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n317_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n835_), .B2(new_n832_), .ZN(G1343gat));
  NOR4_X1   g635(.A1(new_n598_), .A2(new_n494_), .A3(new_n634_), .A4(new_n447_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n810_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n233_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n625_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g642(.A1(new_n838_), .A2(KEYINPUT125), .A3(new_n361_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT125), .B1(new_n838_), .B2(new_n361_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1346gat));
  OR3_X1    g647(.A1(new_n838_), .A2(G162gat), .A3(new_n316_), .ZN(new_n849_));
  OAI21_X1  g648(.A(G162gat), .B1(new_n838_), .B2(new_n834_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1347gat));
  INV_X1    g650(.A(new_n496_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n597_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NOR4_X1   g653(.A1(new_n809_), .A2(new_n626_), .A3(new_n560_), .A4(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT126), .ZN(new_n856_));
  OAI21_X1  g655(.A(G169gat), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n785_), .A2(new_n794_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n802_), .A2(new_n317_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n651_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n853_), .B(new_n634_), .C1(new_n863_), .C2(new_n758_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n864_), .A2(KEYINPUT126), .A3(new_n626_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT127), .B1(new_n857_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT126), .B1(new_n864_), .B2(new_n626_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n855_), .A2(new_n856_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT127), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .A4(G169gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n866_), .A2(KEYINPUT62), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT62), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT127), .B(new_n872_), .C1(new_n857_), .C2(new_n865_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n855_), .A2(new_n519_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n871_), .A2(new_n873_), .A3(new_n874_), .ZN(G1348gat));
  NOR2_X1   g674(.A1(new_n864_), .A2(new_n393_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n416_), .ZN(G1349gat));
  NOR2_X1   g676(.A1(new_n864_), .A2(new_n361_), .ZN(new_n878_));
  MUX2_X1   g677(.A(G183gat), .B(new_n497_), .S(new_n878_), .Z(G1350gat));
  OAI21_X1  g678(.A(G190gat), .B1(new_n864_), .B2(new_n834_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n629_), .A2(new_n400_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n864_), .B2(new_n881_), .ZN(G1351gat));
  NOR2_X1   g681(.A1(new_n809_), .A2(new_n560_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n883_), .A2(new_n494_), .A3(new_n597_), .A4(new_n448_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n626_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n506_), .ZN(G1352gat));
  NOR2_X1   g685(.A1(new_n884_), .A2(new_n393_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n504_), .ZN(G1353gat));
  NOR2_X1   g687(.A1(new_n884_), .A2(new_n361_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n889_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT63), .B(G211gat), .Z(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n889_), .B2(new_n891_), .ZN(G1354gat));
  OAI21_X1  g691(.A(G218gat), .B1(new_n884_), .B2(new_n834_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n316_), .A2(G218gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n884_), .B2(new_n894_), .ZN(G1355gat));
endmodule


