//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_;
  XNOR2_X1  g000(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G127gat), .B(G155gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G183gat), .B(G211gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT77), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G15gat), .ZN(new_n211_));
  INV_X1    g010(.A(G22gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G15gat), .A2(G22gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G1gat), .A2(G8gat), .ZN(new_n215_));
  AOI22_X1  g014(.A1(new_n213_), .A2(new_n214_), .B1(KEYINPUT14), .B2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n210_), .B(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G57gat), .B(G64gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT69), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n218_), .A2(KEYINPUT69), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT11), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G71gat), .B(G78gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n218_), .A2(KEYINPUT69), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n219_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(new_n224_), .A3(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(KEYINPUT11), .B(new_n223_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n229_));
  INV_X1    g028(.A(G231gat), .ZN(new_n230_));
  INV_X1    g029(.A(G233gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n228_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n217_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n228_), .A2(new_n229_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n232_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n217_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n234_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n207_), .B1(new_n242_), .B2(KEYINPUT79), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT79), .ZN(new_n244_));
  AOI211_X1 g043(.A(new_n244_), .B(new_n206_), .C1(new_n237_), .C2(new_n241_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n203_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  NOR3_X1   g045(.A1(new_n235_), .A2(new_n217_), .A3(new_n236_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n240_), .B1(new_n239_), .B2(new_n234_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT79), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n206_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n242_), .A2(KEYINPUT79), .A3(new_n207_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n202_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n242_), .A2(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n246_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT17), .B1(new_n246_), .B2(new_n252_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT37), .ZN(new_n258_));
  INV_X1    g057(.A(G99gat), .ZN(new_n259_));
  INV_X1    g058(.A(G106gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(new_n260_), .A3(KEYINPUT64), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT7), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G99gat), .A2(G106gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT6), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT6), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(G99gat), .A3(G106gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT7), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n268_), .A2(new_n259_), .A3(new_n260_), .A4(KEYINPUT64), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n262_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n271_));
  AND2_X1   g070(.A1(G85gat), .A2(G92gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G85gat), .A2(G92gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(G85gat), .ZN(new_n275_));
  INV_X1    g074(.A(G92gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G85gat), .A2(G92gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(KEYINPUT66), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT68), .B1(new_n270_), .B2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n262_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(new_n274_), .A4(new_n279_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(KEYINPUT8), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(KEYINPUT65), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n262_), .A2(new_n267_), .A3(new_n287_), .A4(new_n269_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT8), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n274_), .A2(new_n279_), .A3(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT67), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n286_), .A2(new_n293_), .A3(new_n288_), .A4(new_n290_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n285_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G29gat), .B(G36gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G43gat), .B(G50gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(KEYINPUT10), .B(G99gat), .Z(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n260_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n277_), .A2(KEYINPUT9), .A3(new_n278_), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n278_), .A2(KEYINPUT9), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .A4(new_n267_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n295_), .A2(new_n298_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n295_), .A2(KEYINPUT73), .A3(new_n298_), .A4(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n295_), .A2(new_n303_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n298_), .B(KEYINPUT15), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT35), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G232gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n309_), .A2(new_n310_), .B1(new_n311_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n308_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n315_), .A2(new_n311_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n318_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n308_), .A2(new_n320_), .A3(new_n316_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G190gat), .B(G218gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT74), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G134gat), .B(G162gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT36), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT75), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n319_), .A2(new_n321_), .A3(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n258_), .B1(new_n329_), .B2(KEYINPUT76), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n325_), .B(KEYINPUT36), .ZN(new_n331_));
  INV_X1    g130(.A(new_n321_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n320_), .B1(new_n308_), .B2(new_n316_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n329_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n334_), .B(new_n329_), .C1(KEYINPUT76), .C2(new_n258_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n257_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n295_), .A2(new_n238_), .A3(new_n303_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G230gat), .A2(G233gat), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT12), .ZN(new_n342_));
  INV_X1    g141(.A(new_n238_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(new_n309_), .B2(new_n343_), .ZN(new_n344_));
  AOI211_X1 g143(.A(KEYINPUT12), .B(new_n238_), .C1(new_n295_), .C2(new_n303_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n341_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n309_), .A2(new_n343_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n339_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n340_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G120gat), .B(G148gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G176gat), .B(G204gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n346_), .A2(new_n350_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n346_), .A2(new_n350_), .A3(KEYINPUT71), .A4(new_n356_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n340_), .B1(new_n347_), .B2(new_n339_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n303_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n264_), .A2(new_n266_), .B1(new_n261_), .B2(KEYINPUT7), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n280_), .B1(new_n269_), .B2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n289_), .B1(new_n365_), .B2(new_n283_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n366_), .A2(new_n281_), .B1(KEYINPUT67), .B2(new_n291_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n363_), .B1(new_n367_), .B2(new_n294_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT12), .B1(new_n368_), .B2(new_n238_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n309_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n362_), .B1(new_n371_), .B2(new_n341_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n372_), .A2(new_n356_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n361_), .A2(KEYINPUT13), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT13), .B1(new_n361_), .B2(new_n373_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n338_), .A2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT80), .Z(new_n378_));
  NAND2_X1  g177(.A1(G229gat), .A2(G233gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n240_), .A2(new_n310_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n217_), .A2(new_n381_), .A3(new_n298_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n217_), .B2(new_n298_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n379_), .B(new_n380_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G113gat), .B(G141gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G169gat), .B(G197gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  NOR2_X1   g187(.A1(new_n217_), .A2(new_n298_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n384_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n390_), .B2(new_n382_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n385_), .B(new_n388_), .C1(new_n391_), .C2(new_n379_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  OAI22_X1  g192(.A1(new_n383_), .A2(new_n384_), .B1(new_n217_), .B2(new_n298_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n379_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n388_), .B1(new_n396_), .B2(new_n385_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n393_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(G71gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G99gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(G15gat), .B(G43gat), .Z(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT84), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n402_), .B(new_n404_), .Z(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G169gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G183gat), .A2(G190gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT23), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT23), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(G183gat), .A3(G190gat), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT83), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n409_), .B2(KEYINPUT23), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT82), .B(G190gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n417_), .A2(G183gat), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n408_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n410_), .A2(new_n412_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G169gat), .A2(G176gat), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n417_), .B2(KEYINPUT26), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT25), .B(G183gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n420_), .B(new_n425_), .C1(new_n427_), .C2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n419_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT30), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT85), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n432_), .A2(KEYINPUT85), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n406_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n405_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G127gat), .B(G134gat), .Z(new_n438_));
  XOR2_X1   g237(.A(G113gat), .B(G120gat), .Z(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n440_), .B(KEYINPUT31), .Z(new_n441_));
  AND3_X1   g240(.A1(new_n436_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n441_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(G155gat), .A2(G162gat), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G155gat), .A2(G162gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G141gat), .A2(G148gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT3), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G141gat), .A2(G148gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT87), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT2), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n453_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n447_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(KEYINPUT1), .A2(new_n445_), .B1(new_n448_), .B2(KEYINPUT86), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n451_), .A2(KEYINPUT86), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(G141gat), .B2(G148gat), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT1), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n447_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(KEYINPUT88), .B(new_n447_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n460_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT29), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n471_));
  INV_X1    g270(.A(G204gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(G197gat), .ZN(new_n473_));
  INV_X1    g272(.A(G197gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G204gat), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n473_), .A2(new_n475_), .A3(KEYINPUT90), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT21), .B1(new_n473_), .B2(KEYINPUT90), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n471_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G211gat), .B(G218gat), .Z(new_n479_));
  INV_X1    g278(.A(KEYINPUT21), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n473_), .A2(new_n475_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n479_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n473_), .A2(new_n475_), .A3(KEYINPUT90), .ZN(new_n483_));
  OR3_X1    g282(.A1(new_n474_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n483_), .A2(new_n484_), .A3(KEYINPUT91), .A4(KEYINPUT21), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n478_), .A2(new_n482_), .A3(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n481_), .A2(new_n480_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n479_), .A2(KEYINPUT92), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G211gat), .B(G218gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT92), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n487_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n486_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n470_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G228gat), .A2(G233gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n495_), .B(KEYINPUT89), .Z(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n470_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT28), .B1(new_n469_), .B2(KEYINPUT29), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n458_), .A2(new_n459_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT28), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT29), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .A4(new_n468_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G22gat), .B(G50gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n501_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n501_), .A2(new_n505_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n506_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G78gat), .B(G106gat), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n500_), .A2(new_n507_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n511_), .B(KEYINPUT93), .Z(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n500_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n500_), .A2(new_n514_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT94), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n510_), .B2(new_n507_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n515_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n515_), .B1(new_n518_), .B2(new_n516_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n512_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n486_), .A2(new_n419_), .A3(new_n492_), .A4(new_n430_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n486_), .A2(new_n492_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n423_), .A2(new_n424_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n421_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT26), .B(G190gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT95), .ZN(new_n529_));
  INV_X1    g328(.A(new_n426_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT95), .ZN(new_n531_));
  NAND2_X1  g330(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n529_), .A2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n527_), .B1(new_n534_), .B2(new_n428_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n413_), .A2(new_n415_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n420_), .B1(G183gat), .B2(G190gat), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n535_), .A2(new_n536_), .B1(new_n408_), .B2(new_n537_), .ZN(new_n538_));
  OAI211_X1 g337(.A(KEYINPUT20), .B(new_n523_), .C1(new_n524_), .C2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G226gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT19), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT20), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n524_), .B2(new_n538_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n541_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n493_), .A2(new_n431_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G8gat), .B(G36gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G64gat), .B(G92gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT32), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n542_), .A2(new_n547_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n544_), .A2(new_n546_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n541_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n528_), .A2(KEYINPUT95), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n531_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n428_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n536_), .A3(new_n425_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n537_), .A2(new_n408_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n543_), .B1(new_n562_), .B2(new_n493_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(new_n545_), .A3(new_n523_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n556_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n554_), .B1(new_n566_), .B2(new_n553_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n440_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n469_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n502_), .A2(new_n440_), .A3(new_n468_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G225gat), .A2(G233gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n440_), .B1(new_n502_), .B2(new_n468_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT4), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n572_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n569_), .A2(new_n570_), .A3(KEYINPUT4), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G1gat), .B(G29gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(G85gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT0), .B(G57gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n583_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n573_), .A2(new_n578_), .A3(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n567_), .A2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n577_), .B(new_n572_), .C1(KEYINPUT4), .C2(new_n569_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n571_), .A2(G225gat), .A3(G233gat), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n583_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n586_), .A2(new_n593_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n571_), .A2(new_n572_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(new_n585_), .A3(new_n592_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n591_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n552_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n545_), .B1(new_n563_), .B2(new_n523_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n560_), .A2(new_n486_), .A3(new_n492_), .A4(new_n561_), .ZN(new_n600_));
  AND4_X1   g399(.A1(KEYINPUT20), .A2(new_n546_), .A3(new_n545_), .A4(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n598_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n542_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT97), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n602_), .A2(new_n603_), .A3(KEYINPUT97), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n597_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n588_), .B1(new_n606_), .B2(KEYINPUT99), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT99), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n597_), .B(new_n608_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n522_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n565_), .A2(new_n598_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT100), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(KEYINPUT27), .A4(new_n603_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n603_), .A2(KEYINPUT27), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n552_), .B1(new_n556_), .B2(new_n564_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT100), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n602_), .A2(new_n603_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n613_), .B(new_n616_), .C1(KEYINPUT27), .C2(new_n617_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n587_), .B(new_n512_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n444_), .B1(new_n610_), .B2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n522_), .A2(new_n618_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n587_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n444_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n398_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n378_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n587_), .A2(G1gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(KEYINPUT38), .A3(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n605_), .A2(new_n604_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n589_), .A2(new_n590_), .A3(new_n583_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n592_), .B1(new_n595_), .B2(new_n585_), .ZN(new_n632_));
  AND4_X1   g431(.A1(new_n573_), .A2(new_n578_), .A3(new_n585_), .A4(new_n592_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n631_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT99), .B1(new_n630_), .B2(new_n634_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n567_), .A2(new_n587_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n609_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n620_), .B1(new_n637_), .B2(new_n521_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n444_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n625_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n335_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n398_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n376_), .A2(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n641_), .A2(new_n257_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n623_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G1gat), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT38), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n378_), .A2(new_n626_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n628_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n647_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n629_), .A2(new_n646_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(G1324gat));
  INV_X1    g452(.A(new_n618_), .ZN(new_n654_));
  OR3_X1    g453(.A1(new_n648_), .A2(G8gat), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n644_), .A2(new_n618_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n656_), .A2(new_n657_), .A3(G8gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n656_), .B2(G8gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n655_), .B(KEYINPUT40), .C1(new_n658_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  AOI21_X1  g463(.A(new_n211_), .B1(new_n644_), .B2(new_n639_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT41), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n627_), .A2(new_n211_), .A3(new_n639_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1326gat));
  AOI21_X1  g467(.A(new_n212_), .B1(new_n644_), .B2(new_n522_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT42), .Z(new_n670_));
  NOR2_X1   g469(.A1(new_n521_), .A2(G22gat), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT102), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n648_), .B2(new_n672_), .ZN(G1327gat));
  OR2_X1    g472(.A1(new_n374_), .A2(new_n375_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n335_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n257_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n257_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT105), .B1(new_n678_), .B2(new_n335_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n674_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n626_), .A2(new_n680_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n681_), .A2(G29gat), .A3(new_n587_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n643_), .A2(new_n678_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n336_), .A2(KEYINPUT104), .A3(new_n337_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT104), .B1(new_n336_), .B2(new_n337_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n684_), .B1(new_n640_), .B2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n336_), .A2(new_n337_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n689_), .A2(KEYINPUT43), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n683_), .B1(new_n688_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  OAI211_X1 g493(.A(KEYINPUT44), .B(new_n683_), .C1(new_n688_), .C2(new_n691_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n623_), .A3(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n682_), .B1(new_n696_), .B2(G29gat), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  AOI211_X1 g498(.A(KEYINPUT106), .B(new_n682_), .C1(new_n696_), .C2(G29gat), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1328gat));
  NAND3_X1  g500(.A1(new_n694_), .A2(new_n618_), .A3(new_n695_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G36gat), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n654_), .A2(G36gat), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n680_), .A2(new_n640_), .A3(new_n642_), .A4(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT107), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n626_), .A2(new_n707_), .A3(new_n680_), .A4(new_n704_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n706_), .A2(KEYINPUT45), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT45), .B1(new_n706_), .B2(new_n708_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n703_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n703_), .B2(new_n711_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1329gat));
  NAND4_X1  g514(.A1(new_n694_), .A2(G43gat), .A3(new_n639_), .A4(new_n695_), .ZN(new_n716_));
  INV_X1    g515(.A(G43gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n717_), .B1(new_n681_), .B2(new_n444_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(G1330gat));
  NAND3_X1  g520(.A1(new_n694_), .A2(new_n522_), .A3(new_n695_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G50gat), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n521_), .A2(G50gat), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT110), .Z(new_n725_));
  OAI21_X1  g524(.A(new_n723_), .B1(new_n681_), .B2(new_n725_), .ZN(G1331gat));
  NOR2_X1   g525(.A1(new_n376_), .A2(new_n642_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n640_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n338_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(G57gat), .B1(new_n730_), .B2(new_n623_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n678_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n675_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n733_), .A2(G57gat), .A3(new_n623_), .A4(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(KEYINPUT111), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(KEYINPUT111), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n731_), .A2(new_n736_), .A3(new_n737_), .ZN(G1332gat));
  NAND2_X1  g537(.A1(new_n733_), .A2(new_n734_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G64gat), .B1(new_n739_), .B2(new_n654_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT48), .ZN(new_n741_));
  OR3_X1    g540(.A1(new_n729_), .A2(G64gat), .A3(new_n654_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT112), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n741_), .A2(new_n745_), .A3(new_n742_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n739_), .B2(new_n444_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT49), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n730_), .A2(new_n400_), .A3(new_n639_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1334gat));
  OAI21_X1  g550(.A(G78gat), .B1(new_n739_), .B2(new_n521_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n752_), .B(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n521_), .A2(G78gat), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT114), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n729_), .B2(new_n756_), .ZN(G1335gat));
  NAND2_X1  g556(.A1(new_n640_), .A2(new_n727_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n759_));
  AOI21_X1  g558(.A(G85gat), .B1(new_n759_), .B2(new_n623_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n688_), .A2(new_n691_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n727_), .A2(new_n257_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n623_), .A2(G85gat), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT115), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n760_), .B1(new_n763_), .B2(new_n765_), .ZN(G1336gat));
  NAND3_X1  g565(.A1(new_n759_), .A2(new_n276_), .A3(new_n618_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n763_), .A2(new_n618_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n769_), .B2(new_n276_), .ZN(G1337gat));
  AND3_X1   g569(.A1(new_n759_), .A2(new_n639_), .A3(new_n299_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n763_), .A2(new_n639_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(G99gat), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n773_), .B(new_n774_), .ZN(G1338gat));
  NAND3_X1  g574(.A1(new_n759_), .A2(new_n260_), .A3(new_n522_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n762_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n522_), .B(new_n777_), .C1(new_n688_), .C2(new_n691_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(new_n779_), .A3(G106gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G106gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n776_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g582(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n388_), .B1(new_n394_), .B2(new_n379_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n390_), .A2(new_n382_), .B1(new_n240_), .B2(new_n310_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n395_), .B1(new_n787_), .B2(KEYINPUT117), .ZN(new_n788_));
  OAI211_X1 g587(.A(KEYINPUT117), .B(new_n380_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n392_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n361_), .B2(new_n373_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT71), .B1(new_n372_), .B2(new_n356_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n360_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n642_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n346_), .A2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n339_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n349_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n341_), .B(KEYINPUT55), .C1(new_n344_), .C2(new_n345_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n802_), .A2(new_n355_), .B1(KEYINPUT116), .B2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n796_), .A2(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n802_), .A2(KEYINPUT116), .A3(new_n803_), .A4(new_n355_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n793_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n785_), .B1(new_n807_), .B2(new_n675_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n804_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n398_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n806_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n793_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(KEYINPUT57), .A3(new_n335_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n802_), .A2(new_n355_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT56), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n792_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n802_), .A2(new_n803_), .A3(new_n355_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n816_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n816_), .A2(new_n817_), .A3(KEYINPUT58), .A4(new_n818_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n821_), .A2(new_n337_), .A3(new_n336_), .A4(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n808_), .A2(new_n814_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n257_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT54), .B1(new_n377_), .B2(new_n642_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n338_), .A2(new_n376_), .A3(new_n827_), .A4(new_n398_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n825_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n622_), .A2(new_n623_), .A3(new_n639_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT118), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n784_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n824_), .A2(new_n257_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n832_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(KEYINPUT120), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n834_), .A2(new_n835_), .A3(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT121), .B1(new_n833_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n784_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n830_), .A2(new_n832_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n841_), .B(new_n842_), .C1(new_n843_), .C2(new_n837_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n839_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(G113gat), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n398_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n830_), .A2(KEYINPUT119), .A3(new_n832_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n850_), .A3(new_n642_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n845_), .A2(new_n847_), .B1(new_n846_), .B2(new_n851_), .ZN(G1340gat));
  OAI21_X1  g651(.A(new_n841_), .B1(new_n843_), .B2(new_n837_), .ZN(new_n853_));
  OAI21_X1  g652(.A(G120gat), .B1(new_n853_), .B2(new_n376_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n376_), .A2(KEYINPUT60), .ZN(new_n855_));
  MUX2_X1   g654(.A(new_n855_), .B(KEYINPUT60), .S(G120gat), .Z(new_n856_));
  NAND3_X1  g655(.A1(new_n848_), .A2(new_n850_), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n858_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n854_), .B1(new_n859_), .B2(new_n860_), .ZN(G1341gat));
  INV_X1    g660(.A(G127gat), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n257_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n848_), .A2(new_n850_), .A3(new_n678_), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n845_), .A2(new_n863_), .B1(new_n862_), .B2(new_n864_), .ZN(G1342gat));
  XOR2_X1   g664(.A(KEYINPUT123), .B(G134gat), .Z(new_n866_));
  NOR2_X1   g665(.A1(new_n689_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(G134gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n848_), .A2(new_n850_), .A3(new_n675_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n845_), .A2(new_n867_), .B1(new_n868_), .B2(new_n869_), .ZN(G1343gat));
  NAND3_X1  g669(.A1(new_n522_), .A2(new_n623_), .A3(new_n444_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n834_), .A2(new_n618_), .A3(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n642_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT124), .B(G141gat), .Z(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n674_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g676(.A1(new_n872_), .A2(new_n678_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT61), .B(G155gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  AOI21_X1  g679(.A(G162gat), .B1(new_n872_), .B2(new_n675_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n687_), .A2(G162gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n872_), .B2(new_n882_), .ZN(G1347gat));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n624_), .A2(new_n618_), .ZN(new_n885_));
  NOR4_X1   g684(.A1(new_n834_), .A2(new_n522_), .A3(new_n398_), .A4(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT22), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G169gat), .ZN(new_n889_));
  INV_X1    g688(.A(G169gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n886_), .B2(new_n884_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n888_), .B2(new_n891_), .ZN(G1348gat));
  NAND2_X1  g691(.A1(new_n830_), .A2(new_n521_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n885_), .ZN(new_n894_));
  AOI21_X1  g693(.A(G176gat), .B1(new_n894_), .B2(new_n674_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(KEYINPUT125), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n834_), .A2(new_n522_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT125), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n896_), .A2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n885_), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n674_), .A2(G176gat), .A3(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n895_), .B1(new_n900_), .B2(new_n902_), .ZN(G1349gat));
  NAND4_X1  g702(.A1(new_n896_), .A2(new_n899_), .A3(new_n678_), .A4(new_n901_), .ZN(new_n904_));
  INV_X1    g703(.A(G183gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n257_), .A2(new_n428_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n904_), .A2(new_n905_), .B1(new_n894_), .B2(new_n906_), .ZN(G1350gat));
  AOI21_X1  g706(.A(new_n335_), .B1(new_n529_), .B2(new_n533_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n897_), .A2(new_n901_), .A3(new_n908_), .ZN(new_n909_));
  NOR4_X1   g708(.A1(new_n834_), .A2(new_n522_), .A3(new_n689_), .A4(new_n885_), .ZN(new_n910_));
  INV_X1    g709(.A(G190gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n909_), .B(KEYINPUT126), .C1(new_n911_), .C2(new_n910_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1351gat));
  NOR2_X1   g715(.A1(new_n654_), .A2(new_n639_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n619_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n834_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n642_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n674_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g723(.A(new_n919_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n830_), .A2(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n257_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT127), .B1(new_n926_), .B2(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n920_), .A2(new_n931_), .A3(new_n927_), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n929_), .A2(new_n930_), .A3(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n930_), .B1(new_n929_), .B2(new_n932_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1354gat));
  OR3_X1    g734(.A1(new_n926_), .A2(G218gat), .A3(new_n335_), .ZN(new_n936_));
  OAI21_X1  g735(.A(G218gat), .B1(new_n926_), .B2(new_n689_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1355gat));
endmodule


