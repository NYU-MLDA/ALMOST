//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT78), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(KEYINPUT24), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT23), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT26), .B(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(G183gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT25), .B1(new_n210_), .B2(KEYINPUT77), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n210_), .A2(KEYINPUT25), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n209_), .B(new_n211_), .C1(new_n212_), .C2(KEYINPUT77), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n208_), .B(new_n213_), .C1(KEYINPUT24), .C2(new_n203_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n207_), .B1(G183gat), .B2(G190gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n215_), .A2(new_n204_), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(G169gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT22), .B1(new_n218_), .B2(KEYINPUT79), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n218_), .A2(KEYINPUT22), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n217_), .B(new_n219_), .C1(new_n220_), .C2(KEYINPUT79), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n216_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n214_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G227gat), .A2(G233gat), .ZN(new_n224_));
  INV_X1    g023(.A(G15gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT30), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n223_), .B(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G71gat), .B(G99gat), .Z(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G43gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n228_), .B(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G127gat), .B(G134gat), .Z(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G120gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n236_), .B(KEYINPUT31), .Z(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT82), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n231_), .A2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n237_), .A2(KEYINPUT82), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n231_), .B1(new_n241_), .B2(new_n239_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G211gat), .B(G218gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G197gat), .B(G204gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT91), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n245_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n249_), .A2(KEYINPUT21), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n249_), .B(KEYINPUT21), .C1(new_n247_), .C2(new_n245_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G155gat), .B(G162gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G141gat), .A2(G148gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT83), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT84), .B(KEYINPUT2), .Z(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT85), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT85), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n261_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n262_));
  INV_X1    g061(.A(G141gat), .ZN(new_n263_));
  INV_X1    g062(.A(G148gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT3), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(G141gat), .B2(G148gat), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n260_), .A2(new_n262_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n258_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n254_), .B1(new_n269_), .B2(KEYINPUT86), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(KEYINPUT86), .B2(new_n269_), .ZN(new_n271_));
  AND2_X1   g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n272_), .A2(KEYINPUT1), .B1(new_n263_), .B2(new_n264_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n256_), .B(new_n273_), .C1(KEYINPUT1), .C2(new_n254_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n253_), .B1(new_n275_), .B2(KEYINPUT29), .ZN(new_n276_));
  INV_X1    g075(.A(G228gat), .ZN(new_n277_));
  INV_X1    g076(.A(G233gat), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(KEYINPUT89), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(KEYINPUT89), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n277_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT90), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n276_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G78gat), .B(G106gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n287_), .B(KEYINPUT92), .Z(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT93), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n286_), .A2(KEYINPUT93), .A3(new_n288_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n291_), .B(new_n292_), .C1(new_n288_), .C2(new_n286_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n275_), .A2(KEYINPUT29), .ZN(new_n294_));
  XOR2_X1   g093(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G22gat), .B(G50gat), .Z(new_n297_));
  OR2_X1    g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n297_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT88), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n298_), .A2(new_n302_), .A3(new_n299_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n293_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n285_), .A2(new_n287_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n300_), .A2(new_n289_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n275_), .B(new_n236_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT4), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n271_), .A2(new_n274_), .ZN(new_n313_));
  OR3_X1    g112(.A1(new_n313_), .A2(KEYINPUT4), .A3(new_n236_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT96), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n314_), .A2(new_n315_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n310_), .B(new_n312_), .C1(new_n316_), .C2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G1gat), .B(G29gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT97), .B(G85gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT0), .B(G57gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  NAND2_X1  g122(.A1(new_n311_), .A2(new_n309_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n318_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT33), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n202_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n209_), .ZN(new_n329_));
  XOR2_X1   g128(.A(KEYINPUT25), .B(G183gat), .Z(new_n330_));
  OAI221_X1 g129(.A(new_n208_), .B1(KEYINPUT24), .B2(new_n328_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT22), .B(G169gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n216_), .B1(G176gat), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n331_), .A2(new_n253_), .A3(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n335_), .A2(KEYINPUT20), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT19), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n223_), .A2(new_n252_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT20), .B1(new_n223_), .B2(new_n252_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n253_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n338_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT95), .ZN(new_n346_));
  XOR2_X1   g145(.A(G8gat), .B(G36gat), .Z(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G64gat), .B(G92gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n345_), .A2(new_n346_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n351_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n341_), .A2(new_n353_), .A3(new_n344_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n346_), .B1(new_n345_), .B2(new_n351_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n325_), .A2(new_n326_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n323_), .B1(new_n311_), .B2(new_n310_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n312_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n359_), .B1(new_n360_), .B2(new_n310_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n327_), .A2(new_n357_), .A3(new_n358_), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n318_), .A2(new_n324_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n323_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n325_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n353_), .A2(KEYINPUT32), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n341_), .A2(new_n367_), .A3(new_n344_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n342_), .A2(new_n343_), .A3(new_n338_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n336_), .A2(new_n340_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n338_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n366_), .B(new_n368_), .C1(new_n367_), .C2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n308_), .B1(new_n362_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n307_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(new_n304_), .B2(new_n293_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n377_));
  OAI211_X1 g176(.A(KEYINPUT27), .B(new_n354_), .C1(new_n371_), .C2(new_n353_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n375_), .A2(new_n379_), .A3(new_n366_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n244_), .B1(new_n373_), .B2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n308_), .A2(new_n379_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n366_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n243_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G29gat), .B(G36gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G43gat), .B(G50gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n388_), .B(KEYINPUT15), .Z(new_n389_));
  XOR2_X1   g188(.A(G15gat), .B(G22gat), .Z(new_n390_));
  XOR2_X1   g189(.A(KEYINPUT70), .B(G1gat), .Z(new_n391_));
  XOR2_X1   g190(.A(KEYINPUT71), .B(G8gat), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n390_), .B1(new_n393_), .B2(KEYINPUT14), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G1gat), .B(G8gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n389_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n388_), .B2(new_n396_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G229gat), .A2(G233gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n396_), .B(new_n388_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(G229gat), .A3(G233gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G113gat), .B(G141gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G169gat), .B(G197gat), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n404_), .B(new_n405_), .Z(new_n406_));
  XNOR2_X1  g205(.A(new_n403_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT75), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n408_), .A2(KEYINPUT76), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(KEYINPUT76), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n385_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G99gat), .A2(G106gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT6), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(G99gat), .A3(G106gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n418_));
  INV_X1    g217(.A(G106gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G85gat), .ZN(new_n422_));
  INV_X1    g221(.A(G92gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G85gat), .A2(G92gat), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(KEYINPUT9), .A3(new_n425_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n425_), .A2(KEYINPUT9), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n417_), .A2(new_n421_), .A3(new_n426_), .A4(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n424_), .A2(new_n425_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n414_), .A2(new_n416_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT7), .ZN(new_n433_));
  INV_X1    g232(.A(G99gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n434_), .A3(new_n419_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n431_), .B1(new_n432_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT8), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n415_), .B1(G99gat), .B2(G106gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n413_), .A2(KEYINPUT6), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n436_), .B(new_n435_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT8), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(new_n431_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n429_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n388_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G232gat), .A2(G233gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT34), .ZN(new_n448_));
  INV_X1    g247(.A(new_n436_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AOI211_X1 g250(.A(KEYINPUT8), .B(new_n430_), .C1(new_n451_), .C2(new_n417_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n443_), .B1(new_n442_), .B2(new_n431_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT66), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT66), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n439_), .A2(new_n455_), .A3(new_n444_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n429_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  OAI221_X1 g256(.A(new_n446_), .B1(KEYINPUT35), .B2(new_n448_), .C1(new_n457_), .C2(new_n389_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n448_), .A2(KEYINPUT35), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n459_), .B(KEYINPUT68), .Z(new_n460_));
  XNOR2_X1  g259(.A(new_n458_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G190gat), .B(G218gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G134gat), .B(G162gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n464_), .A2(KEYINPUT36), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n464_), .B(KEYINPUT36), .Z(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n461_), .A2(new_n468_), .ZN(new_n469_));
  OR3_X1    g268(.A1(new_n466_), .A2(new_n469_), .A3(KEYINPUT37), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n467_), .B(KEYINPUT69), .Z(new_n471_));
  NOR2_X1   g270(.A1(new_n461_), .A2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT37), .B1(new_n466_), .B2(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT17), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G127gat), .B(G155gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT16), .ZN(new_n477_));
  XOR2_X1   g276(.A(G183gat), .B(G211gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G57gat), .B(G64gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G71gat), .B(G78gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(KEYINPUT11), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(KEYINPUT11), .ZN(new_n483_));
  INV_X1    g282(.A(new_n481_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n480_), .A2(KEYINPUT11), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n482_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G231gat), .A2(G233gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(new_n396_), .ZN(new_n490_));
  AOI211_X1 g289(.A(new_n475_), .B(new_n479_), .C1(new_n490_), .C2(KEYINPUT72), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n491_), .B1(KEYINPUT72), .B2(new_n490_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n479_), .B(new_n475_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT73), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n490_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n474_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(G230gat), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n487_), .B(new_n428_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT64), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT64), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n445_), .A2(new_n501_), .A3(new_n487_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n428_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n487_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n503_), .A2(KEYINPUT65), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n500_), .A2(new_n502_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT65), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AOI211_X1 g308(.A(new_n498_), .B(new_n278_), .C1(new_n506_), .C2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT67), .B(KEYINPUT12), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n452_), .A2(new_n453_), .A3(KEYINPUT66), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n455_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n428_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n505_), .A2(KEYINPUT12), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n513_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n498_), .A2(new_n278_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(new_n445_), .B2(new_n487_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n510_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G120gat), .B(G148gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT5), .ZN(new_n526_));
  XOR2_X1   g325(.A(G176gat), .B(G204gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  OR3_X1    g328(.A1(new_n510_), .A2(new_n523_), .A3(new_n528_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT13), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(KEYINPUT13), .A3(new_n530_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n497_), .A2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n536_), .B(KEYINPUT74), .Z(new_n537_));
  AND2_X1   g336(.A1(new_n412_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n391_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n366_), .A3(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n466_), .A2(new_n469_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(new_n496_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n385_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n408_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n535_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT100), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT100), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n535_), .A2(new_n550_), .A3(new_n547_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n546_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(G1gat), .B1(new_n554_), .B2(new_n383_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n542_), .A2(new_n555_), .ZN(G1324gat));
  INV_X1    g355(.A(new_n392_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n538_), .A2(new_n557_), .A3(new_n379_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT39), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n553_), .A2(new_n379_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n559_), .B1(new_n560_), .B2(G8gat), .ZN(new_n561_));
  INV_X1    g360(.A(G8gat), .ZN(new_n562_));
  AOI211_X1 g361(.A(KEYINPUT39), .B(new_n562_), .C1(new_n553_), .C2(new_n379_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n558_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT40), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OAI211_X1 g365(.A(KEYINPUT40), .B(new_n558_), .C1(new_n561_), .C2(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(G1325gat));
  NAND3_X1  g367(.A1(new_n538_), .A2(new_n225_), .A3(new_n243_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT101), .Z(new_n570_));
  AOI21_X1  g369(.A(new_n225_), .B1(new_n553_), .B2(new_n243_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT41), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(G1326gat));
  INV_X1    g372(.A(G22gat), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n574_), .B1(new_n553_), .B2(new_n308_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n538_), .A2(new_n574_), .A3(new_n308_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(G1327gat));
  NAND4_X1  g378(.A1(new_n412_), .A2(new_n535_), .A3(new_n496_), .A4(new_n543_), .ZN(new_n580_));
  OR3_X1    g379(.A1(new_n580_), .A2(G29gat), .A3(new_n383_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n549_), .A2(new_n551_), .A3(new_n496_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT103), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT43), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n385_), .B2(new_n474_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n474_), .ZN(new_n587_));
  AOI211_X1 g386(.A(KEYINPUT43), .B(new_n587_), .C1(new_n381_), .C2(new_n384_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n584_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT44), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n584_), .B(KEYINPUT44), .C1(new_n586_), .C2(new_n588_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n366_), .A3(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(KEYINPUT104), .ZN(new_n594_));
  OAI21_X1  g393(.A(G29gat), .B1(new_n593_), .B2(KEYINPUT104), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n581_), .B1(new_n594_), .B2(new_n595_), .ZN(G1328gat));
  NAND3_X1  g395(.A1(new_n591_), .A2(new_n379_), .A3(new_n592_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(G36gat), .ZN(new_n598_));
  INV_X1    g397(.A(new_n379_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n599_), .A2(G36gat), .ZN(new_n600_));
  OR3_X1    g399(.A1(new_n580_), .A2(KEYINPUT45), .A3(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT45), .B1(new_n580_), .B2(new_n600_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT46), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n598_), .A2(new_n603_), .A3(KEYINPUT46), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(G1329gat));
  NOR3_X1   g407(.A1(new_n580_), .A2(G43gat), .A3(new_n244_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n591_), .A2(new_n243_), .A3(new_n592_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n610_), .B2(G43gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n612_), .ZN(new_n614_));
  AOI211_X1 g413(.A(new_n609_), .B(new_n614_), .C1(new_n610_), .C2(G43gat), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n613_), .A2(new_n615_), .ZN(G1330gat));
  NAND3_X1  g415(.A1(new_n591_), .A2(new_n308_), .A3(new_n592_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(G50gat), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n375_), .A2(G50gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT106), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n618_), .B1(new_n580_), .B2(new_n620_), .ZN(G1331gat));
  INV_X1    g420(.A(new_n535_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n385_), .A2(new_n408_), .A3(new_n622_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n623_), .A2(new_n496_), .A3(new_n474_), .ZN(new_n624_));
  AOI21_X1  g423(.A(G57gat), .B1(new_n624_), .B2(new_n366_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT107), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n545_), .A2(new_n535_), .A3(new_n411_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n366_), .A2(G57gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n626_), .B1(new_n627_), .B2(new_n628_), .ZN(G1332gat));
  INV_X1    g428(.A(G64gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n627_), .B2(new_n379_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT48), .Z(new_n632_));
  NAND3_X1  g431(.A1(new_n624_), .A2(new_n630_), .A3(new_n379_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1333gat));
  INV_X1    g433(.A(G71gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n627_), .B2(new_n243_), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n624_), .A2(new_n635_), .A3(new_n243_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1334gat));
  INV_X1    g439(.A(G78gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n624_), .A2(new_n641_), .A3(new_n308_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT50), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n627_), .A2(new_n308_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n644_), .B2(G78gat), .ZN(new_n645_));
  AOI211_X1 g444(.A(KEYINPUT50), .B(new_n641_), .C1(new_n627_), .C2(new_n308_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT109), .ZN(G1335gat));
  INV_X1    g447(.A(new_n496_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n535_), .A2(new_n547_), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n650_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G85gat), .B1(new_n651_), .B2(new_n383_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n543_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n623_), .A2(new_n649_), .A3(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(new_n422_), .A3(new_n366_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(G1336gat));
  OAI21_X1  g455(.A(G92gat), .B1(new_n651_), .B2(new_n599_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n654_), .A2(new_n423_), .A3(new_n379_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1337gat));
  OAI21_X1  g458(.A(G99gat), .B1(new_n651_), .B2(new_n244_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n243_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT110), .B1(new_n654_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g463(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n308_), .B(new_n650_), .C1(new_n586_), .C2(new_n588_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT111), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(G106gat), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT52), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n668_), .B1(new_n667_), .B2(G106gat), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n667_), .A2(G106gat), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT52), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(KEYINPUT111), .A3(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n654_), .A2(new_n419_), .A3(new_n308_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n666_), .B1(new_n672_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n671_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(KEYINPUT52), .A3(new_n669_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n680_), .A2(new_n675_), .A3(new_n676_), .A4(new_n665_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(G1339gat));
  INV_X1    g481(.A(KEYINPUT113), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n411_), .A2(new_n536_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n684_), .B2(KEYINPUT54), .ZN(new_n685_));
  OR4_X1    g484(.A1(new_n683_), .A2(new_n411_), .A3(new_n536_), .A4(KEYINPUT54), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(KEYINPUT54), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n685_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT114), .B1(new_n519_), .B2(new_n507_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n511_), .B1(new_n445_), .B2(new_n487_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n690_), .B1(new_n457_), .B2(new_n517_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT114), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n691_), .A2(new_n692_), .A3(new_n503_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n520_), .B1(new_n689_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT115), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT115), .B(new_n520_), .C1(new_n689_), .C2(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT55), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n522_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n519_), .A2(KEYINPUT55), .A3(new_n521_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT116), .B1(new_n698_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT116), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n705_), .B(new_n702_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n528_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT56), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT56), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n709_), .B(new_n528_), .C1(new_n704_), .C2(new_n706_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n708_), .A2(new_n547_), .A3(new_n530_), .A4(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT117), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n530_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n707_), .B2(KEYINPUT56), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n715_), .A2(KEYINPUT117), .A3(new_n547_), .A4(new_n710_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n403_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n398_), .A2(G229gat), .A3(G233gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n406_), .B1(new_n401_), .B2(new_n399_), .ZN(new_n719_));
  AOI22_X1  g518(.A1(new_n717_), .A2(new_n406_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n531_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n713_), .A2(new_n716_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n653_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n721_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n543_), .B1(new_n728_), .B2(new_n716_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT57), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n708_), .A2(new_n530_), .A3(new_n710_), .A4(new_n720_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT58), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n715_), .A2(KEYINPUT58), .A3(new_n710_), .A4(new_n720_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n474_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT119), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n733_), .A2(KEYINPUT119), .A3(new_n474_), .A4(new_n734_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n726_), .A2(new_n730_), .A3(new_n737_), .A4(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n688_), .B1(new_n739_), .B2(new_n496_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n382_), .A2(new_n366_), .A3(new_n243_), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT59), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n726_), .A2(new_n730_), .A3(new_n735_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n688_), .B1(new_n743_), .B2(new_n496_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n741_), .A2(KEYINPUT59), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT120), .B1(new_n744_), .B2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n735_), .B1(new_n729_), .B2(new_n724_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n722_), .A2(KEYINPUT57), .A3(new_n653_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n496_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n685_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT120), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n745_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n742_), .A2(new_n747_), .A3(new_n411_), .A4(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(G113gat), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n737_), .B(new_n738_), .C1(new_n729_), .C2(new_n724_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n496_), .B1(new_n757_), .B2(new_n749_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n751_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n741_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n761_), .A2(G113gat), .A3(new_n408_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n756_), .A2(new_n762_), .ZN(G1340gat));
  NAND4_X1  g562(.A1(new_n742_), .A2(new_n747_), .A3(new_n622_), .A4(new_n754_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(G120gat), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT122), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT60), .ZN(new_n767_));
  AOI21_X1  g566(.A(G120gat), .B1(new_n622_), .B2(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT121), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n767_), .B2(G120gat), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n766_), .B1(new_n761_), .B2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n759_), .A2(KEYINPUT122), .A3(new_n760_), .A4(new_n770_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n765_), .A2(new_n774_), .ZN(G1341gat));
  NAND4_X1  g574(.A1(new_n742_), .A2(new_n747_), .A3(new_n649_), .A4(new_n754_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(G127gat), .ZN(new_n777_));
  OR3_X1    g576(.A1(new_n761_), .A2(G127gat), .A3(new_n496_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1342gat));
  NOR3_X1   g578(.A1(new_n740_), .A2(new_n653_), .A3(new_n741_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT123), .B1(new_n780_), .B2(G134gat), .ZN(new_n781_));
  INV_X1    g580(.A(G134gat), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n587_), .A2(new_n782_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n742_), .A2(new_n747_), .A3(new_n754_), .A4(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT123), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n782_), .C1(new_n761_), .C2(new_n653_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n781_), .A2(new_n784_), .A3(new_n786_), .ZN(G1343gat));
  NOR4_X1   g586(.A1(new_n375_), .A2(new_n383_), .A3(new_n379_), .A4(new_n243_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n759_), .A2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(new_n408_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(new_n263_), .ZN(G1344gat));
  NOR2_X1   g590(.A1(new_n789_), .A2(new_n535_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(new_n264_), .ZN(G1345gat));
  NOR2_X1   g592(.A1(new_n789_), .A2(new_n496_), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT61), .B(G155gat), .Z(new_n795_));
  XNOR2_X1  g594(.A(new_n794_), .B(new_n795_), .ZN(G1346gat));
  OAI21_X1  g595(.A(G162gat), .B1(new_n789_), .B2(new_n587_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n653_), .A2(G162gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n789_), .B2(new_n798_), .ZN(G1347gat));
  NOR3_X1   g598(.A1(new_n599_), .A2(new_n366_), .A3(new_n244_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT124), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(new_n308_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n408_), .B(new_n803_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT125), .B1(new_n804_), .B2(new_n218_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n752_), .A2(new_n547_), .A3(new_n802_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT125), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(G169gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(KEYINPUT62), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT62), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT125), .B(new_n810_), .C1(new_n804_), .C2(new_n218_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n804_), .A2(new_n332_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(new_n811_), .A3(new_n812_), .ZN(G1348gat));
  NOR2_X1   g612(.A1(new_n744_), .A2(new_n803_), .ZN(new_n814_));
  AOI21_X1  g613(.A(G176gat), .B1(new_n814_), .B2(new_n622_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n740_), .A2(new_n308_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n801_), .A2(new_n217_), .A3(new_n535_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(G1349gat));
  INV_X1    g617(.A(new_n801_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n816_), .A2(new_n649_), .A3(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n649_), .A2(new_n330_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n820_), .A2(new_n210_), .B1(new_n814_), .B2(new_n821_), .ZN(G1350gat));
  NAND3_X1  g621(.A1(new_n814_), .A2(new_n209_), .A3(new_n543_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n744_), .A2(new_n587_), .A3(new_n803_), .ZN(new_n824_));
  INV_X1    g623(.A(G190gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(G1351gat));
  NAND4_X1  g625(.A1(new_n308_), .A2(new_n383_), .A3(new_n379_), .A4(new_n244_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n740_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n547_), .ZN(new_n829_));
  INV_X1    g628(.A(G197gat), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n830_), .A2(KEYINPUT126), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(KEYINPUT126), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n828_), .A2(KEYINPUT126), .A3(new_n830_), .A4(new_n547_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(G1352gat));
  NAND2_X1  g634(.A1(new_n828_), .A2(new_n622_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g636(.A(new_n496_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT127), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n828_), .A2(new_n839_), .ZN(new_n840_));
  OR2_X1    g639(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(G1354gat));
  INV_X1    g641(.A(G218gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n828_), .A2(new_n843_), .A3(new_n543_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n740_), .A2(new_n587_), .A3(new_n827_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n843_), .ZN(G1355gat));
endmodule


