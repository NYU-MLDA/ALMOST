//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_;
  INV_X1    g000(.A(KEYINPUT101), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(G169gat), .ZN(new_n208_));
  INV_X1    g007(.A(G183gat), .ZN(new_n209_));
  INV_X1    g008(.A(G190gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT23), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(KEYINPUT81), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT81), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n215_), .B(KEYINPUT23), .C1(new_n209_), .C2(new_n210_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n208_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  INV_X1    g022(.A(G176gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT26), .B(G190gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT77), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n227_), .B1(new_n228_), .B2(G183gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n209_), .A2(KEYINPUT77), .A3(KEYINPUT25), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT78), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n228_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n209_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n226_), .B(new_n231_), .C1(new_n235_), .C2(KEYINPUT79), .ZN(new_n236_));
  INV_X1    g035(.A(new_n234_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n238_));
  OAI211_X1 g037(.A(KEYINPUT79), .B(G183gat), .C1(new_n237_), .C2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n220_), .B(new_n225_), .C1(new_n236_), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n211_), .A2(new_n213_), .ZN(new_n242_));
  OR3_X1    g041(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(G183gat), .B1(new_n237_), .B2(new_n238_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT79), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n248_), .A2(new_n239_), .A3(new_n226_), .A4(new_n231_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n220_), .B1(new_n249_), .B2(new_n225_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n219_), .B1(new_n245_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G204gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT90), .B1(new_n252_), .B2(G197gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT90), .ZN(new_n254_));
  INV_X1    g053(.A(G197gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(G204gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(G197gat), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G211gat), .B(G218gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT21), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n261_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT92), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n257_), .A2(new_n260_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT91), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT92), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(new_n262_), .A4(new_n265_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n263_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n269_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n274_), .B1(new_n275_), .B2(new_n264_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n264_), .B1(G197gat), .B2(G204gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n258_), .A2(new_n259_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n277_), .B1(new_n278_), .B2(G197gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT89), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  OAI211_X1 g080(.A(KEYINPUT89), .B(new_n277_), .C1(new_n278_), .C2(G197gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n273_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n251_), .A2(new_n285_), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n268_), .A2(new_n272_), .B1(new_n276_), .B2(new_n283_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n242_), .B1(G183gat), .B2(G190gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n208_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT25), .B(G183gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n226_), .A2(new_n291_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n292_), .A2(new_n225_), .A3(new_n243_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n217_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT96), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT96), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n225_), .A3(new_n243_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n296_), .B1(new_n297_), .B2(new_n217_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n290_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT20), .B1(new_n287_), .B2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n206_), .B1(new_n286_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G8gat), .B(G36gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT18), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G64gat), .B(G92gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n303_), .B(new_n304_), .Z(new_n305_));
  NAND2_X1  g104(.A1(new_n251_), .A2(new_n285_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n205_), .A2(KEYINPUT20), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(new_n287_), .B2(new_n299_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n301_), .A2(new_n305_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT97), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT97), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n301_), .A2(new_n312_), .A3(new_n305_), .A4(new_n309_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n301_), .A2(new_n309_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n305_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n311_), .A2(new_n313_), .A3(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT100), .B(KEYINPUT27), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n225_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT80), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(new_n287_), .A3(new_n219_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT96), .B1(new_n293_), .B2(new_n294_), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n297_), .A2(new_n296_), .A3(new_n217_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n289_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n285_), .A2(new_n325_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n322_), .A2(new_n326_), .A3(KEYINPUT20), .A4(new_n205_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT20), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n290_), .B1(new_n294_), .B2(new_n293_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n328_), .B1(new_n287_), .B2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n205_), .B1(new_n306_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n327_), .B1(new_n331_), .B2(KEYINPUT99), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT99), .ZN(new_n333_));
  AOI211_X1 g132(.A(new_n333_), .B(new_n205_), .C1(new_n306_), .C2(new_n330_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n315_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n310_), .A2(KEYINPUT27), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n317_), .A2(new_n318_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT87), .ZN(new_n338_));
  INV_X1    g137(.A(G141gat), .ZN(new_n339_));
  INV_X1    g138(.A(G148gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n344_), .B1(KEYINPUT1), .B2(new_n345_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n345_), .A2(KEYINPUT1), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n343_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT2), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n342_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT86), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT86), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n342_), .A2(new_n352_), .A3(new_n349_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NOR3_X1   g156(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n354_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G155gat), .B(G162gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n348_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n338_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n361_), .B1(new_n354_), .B2(new_n359_), .ZN(new_n366_));
  NOR4_X1   g165(.A1(new_n366_), .A2(KEYINPUT87), .A3(new_n348_), .A4(KEYINPUT29), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT28), .B(G22gat), .ZN(new_n368_));
  INV_X1    g167(.A(G50gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n365_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n353_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n352_), .B1(new_n342_), .B2(new_n349_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  OR3_X1    g174(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n362_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n348_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n364_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT87), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n363_), .A2(new_n338_), .A3(new_n364_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n370_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT93), .B1(new_n372_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G228gat), .A2(G233gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n363_), .A2(new_n364_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n285_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n385_), .B1(new_n287_), .B2(new_n387_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT94), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n371_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n381_), .A2(new_n382_), .A3(new_n370_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT93), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G78gat), .B(G106gat), .Z(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n397_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT94), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n384_), .A2(new_n391_), .A3(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n393_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n397_), .B(new_n398_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n384_), .A2(new_n391_), .A3(new_n401_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n401_), .B1(new_n384_), .B2(new_n391_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(G85gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT0), .B(G57gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n409_), .B(new_n410_), .Z(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G134gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G127gat), .ZN(new_n414_));
  INV_X1    g213(.A(G127gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G134gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(G120gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(G113gat), .ZN(new_n419_));
  INV_X1    g218(.A(G113gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G120gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G127gat), .B(G134gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G113gat), .B(G120gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n423_), .A2(new_n426_), .A3(KEYINPUT83), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  OAI22_X1  g229(.A1(new_n427_), .A2(new_n430_), .B1(new_n366_), .B2(new_n348_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G225gat), .A2(G233gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n423_), .A2(new_n426_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n378_), .A2(new_n379_), .A3(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT98), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT98), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n431_), .A2(new_n437_), .A3(new_n432_), .A4(new_n434_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n378_), .A2(new_n379_), .A3(new_n433_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n423_), .A2(new_n426_), .A3(KEYINPUT83), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n378_), .A2(new_n379_), .B1(new_n441_), .B2(new_n429_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT4), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT4), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n431_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n432_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n412_), .B1(new_n439_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n432_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n444_), .B1(new_n431_), .B2(new_n434_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n442_), .A2(KEYINPUT4), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n451_), .A2(new_n411_), .A3(new_n436_), .A4(new_n438_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n447_), .A2(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n403_), .A2(new_n407_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n448_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n440_), .A2(new_n442_), .A3(new_n432_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n455_), .A2(new_n411_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n452_), .A2(KEYINPUT33), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n436_), .A2(new_n438_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n411_), .A4(new_n451_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n457_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n462_), .A2(new_n311_), .A3(new_n313_), .A4(new_n316_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n305_), .A2(KEYINPUT32), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n322_), .A2(new_n326_), .A3(KEYINPUT20), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n467_), .A2(new_n206_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n468_), .A2(new_n464_), .B1(new_n452_), .B2(new_n447_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n463_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n403_), .A2(new_n407_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n337_), .A2(new_n454_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n441_), .A2(new_n429_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT31), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT82), .B(G15gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G227gat), .A2(G233gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n251_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n479_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n321_), .A2(new_n219_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G71gat), .B(G99gat), .ZN(new_n484_));
  INV_X1    g283(.A(G43gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT30), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n480_), .A2(new_n487_), .A3(new_n482_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n476_), .B1(new_n491_), .B2(KEYINPUT84), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT84), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n489_), .A2(new_n493_), .A3(new_n490_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT85), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n489_), .A2(new_n493_), .A3(new_n496_), .A4(new_n490_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n492_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n491_), .A2(KEYINPUT84), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n495_), .A2(new_n497_), .B1(new_n499_), .B2(new_n475_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n202_), .B1(new_n473_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n495_), .A2(new_n497_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n492_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n492_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(new_n453_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n317_), .A2(new_n318_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n336_), .A2(new_n335_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n472_), .A3(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n505_), .A2(new_n506_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n454_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n463_), .A2(new_n470_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n515_));
  OAI211_X1 g314(.A(KEYINPUT101), .B(new_n513_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n502_), .A2(new_n512_), .A3(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G29gat), .B(G36gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT67), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n518_), .A2(KEYINPUT67), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(KEYINPUT67), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n520_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT74), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT71), .B(G15gat), .ZN(new_n529_));
  INV_X1    g328(.A(G22gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G1gat), .ZN(new_n532_));
  INV_X1    g331(.A(G8gat), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT14), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G1gat), .B(G8gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n528_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n526_), .B(KEYINPUT15), .ZN(new_n539_));
  INV_X1    g338(.A(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n526_), .B(KEYINPUT74), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n540_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n538_), .A2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n543_), .B1(new_n546_), .B2(new_n542_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT76), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G169gat), .B(G197gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT75), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n548_), .B(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n517_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT102), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT6), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT6), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(G99gat), .A3(G106gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT65), .ZN(new_n562_));
  XOR2_X1   g361(.A(KEYINPUT10), .B(G99gat), .Z(new_n563_));
  INV_X1    g362(.A(G106gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(G85gat), .ZN(new_n566_));
  INV_X1    g365(.A(G92gat), .ZN(new_n567_));
  OR3_X1    g366(.A1(new_n566_), .A2(new_n567_), .A3(KEYINPUT9), .ZN(new_n568_));
  XOR2_X1   g367(.A(G85gat), .B(G92gat), .Z(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT9), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n562_), .A2(new_n565_), .A3(new_n568_), .A4(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT66), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT8), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT7), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(new_n562_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n561_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n573_), .B1(new_n578_), .B2(new_n569_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n572_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G57gat), .B(G64gat), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n582_), .A2(KEYINPUT11), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G71gat), .B(G78gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n583_), .A2(new_n584_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n582_), .A2(KEYINPUT11), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT12), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n581_), .A2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n577_), .A2(new_n579_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(new_n571_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n589_), .B1(new_n594_), .B2(new_n588_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT64), .Z(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n588_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n592_), .A2(new_n595_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n597_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n598_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n594_), .A2(new_n588_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n600_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G120gat), .B(G148gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT5), .ZN(new_n606_));
  XOR2_X1   g405(.A(G176gat), .B(G204gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n604_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT13), .ZN(new_n610_));
  XOR2_X1   g409(.A(G190gat), .B(G218gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT68), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G134gat), .B(G162gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT36), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT34), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n572_), .A2(new_n580_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n539_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n594_), .A2(new_n526_), .ZN(new_n622_));
  OAI211_X1 g421(.A(KEYINPUT35), .B(new_n618_), .C1(new_n621_), .C2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n581_), .A2(new_n539_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT35), .ZN(new_n625_));
  INV_X1    g424(.A(new_n618_), .ZN(new_n626_));
  AOI22_X1  g425(.A1(new_n594_), .A2(new_n526_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n625_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n624_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n616_), .B1(new_n623_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT36), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n614_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT69), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n623_), .A2(new_n630_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT70), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n623_), .A2(KEYINPUT70), .A3(new_n630_), .A4(new_n634_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n631_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT37), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n537_), .B(new_n641_), .Z(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(new_n588_), .ZN(new_n643_));
  XOR2_X1   g442(.A(G127gat), .B(G155gat), .Z(new_n644_));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT17), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(KEYINPUT17), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n643_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(KEYINPUT73), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT73), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n653_), .B1(new_n643_), .B2(new_n649_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n651_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n640_), .A2(new_n656_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n556_), .A2(new_n610_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n453_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n532_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT38), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n454_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n471_), .A2(new_n472_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n501_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n511_), .B1(new_n665_), .B2(KEYINPUT101), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n639_), .B1(new_n666_), .B2(new_n502_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n610_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n554_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n656_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G1gat), .B1(new_n671_), .B2(new_n453_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n660_), .A2(new_n661_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n662_), .A2(new_n672_), .A3(new_n673_), .ZN(G1324gat));
  OAI21_X1  g473(.A(G8gat), .B1(new_n671_), .B2(new_n337_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT39), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n337_), .A2(G8gat), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n658_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n677_), .B1(new_n658_), .B2(new_n678_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n681_), .B(new_n683_), .ZN(G1325gat));
  INV_X1    g483(.A(G15gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n658_), .A2(new_n685_), .A3(new_n501_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G15gat), .B1(new_n671_), .B2(new_n513_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT41), .Z(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1326gat));
  INV_X1    g488(.A(new_n472_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n658_), .A2(new_n530_), .A3(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G22gat), .B1(new_n671_), .B2(new_n472_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT42), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n656_), .A2(new_n639_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n668_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n556_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n659_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n668_), .A2(new_n669_), .A3(new_n655_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n517_), .A2(new_n640_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(KEYINPUT105), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n517_), .A2(new_n640_), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n702_), .B1(new_n706_), .B2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n700_), .B1(new_n711_), .B2(KEYINPUT44), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT37), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n639_), .B(new_n713_), .ZN(new_n714_));
  AOI211_X1 g513(.A(new_n714_), .B(new_n708_), .C1(new_n666_), .C2(new_n502_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n704_), .B1(new_n517_), .B2(new_n640_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n701_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(KEYINPUT106), .A3(new_n718_), .ZN(new_n719_));
  AOI22_X1  g518(.A1(new_n712_), .A2(new_n719_), .B1(KEYINPUT44), .B2(new_n711_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n659_), .A2(G29gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n699_), .B1(new_n720_), .B2(new_n721_), .ZN(G1328gat));
  NOR2_X1   g521(.A1(new_n337_), .A2(G36gat), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OR3_X1    g523(.A1(new_n697_), .A2(KEYINPUT45), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT45), .B1(new_n697_), .B2(new_n724_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n337_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n728_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n712_), .B2(new_n719_), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n730_), .A2(KEYINPUT107), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n337_), .B1(new_n711_), .B2(KEYINPUT44), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n714_), .B1(new_n666_), .B2(new_n502_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n710_), .B1(new_n735_), .B2(new_n704_), .ZN(new_n736_));
  AOI211_X1 g535(.A(new_n700_), .B(KEYINPUT44), .C1(new_n736_), .C2(new_n701_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT106), .B1(new_n717_), .B2(new_n718_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n733_), .B1(new_n739_), .B2(G36gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n727_), .B1(new_n732_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(KEYINPUT46), .B(new_n727_), .C1(new_n732_), .C2(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1329gat));
  NAND3_X1  g544(.A1(new_n720_), .A2(G43gat), .A3(new_n501_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n485_), .B1(new_n697_), .B2(new_n513_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g548(.A1(new_n698_), .A2(new_n369_), .A3(new_n690_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n720_), .A2(new_n690_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n751_), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT108), .B1(new_n751_), .B2(G50gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(G1331gat));
  INV_X1    g553(.A(G57gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n554_), .B1(new_n666_), .B2(new_n502_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n640_), .A2(new_n610_), .A3(new_n656_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n755_), .B1(new_n758_), .B2(new_n453_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT109), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n668_), .A2(new_n669_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n761_), .A2(new_n656_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n667_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n763_), .A2(new_n755_), .A3(new_n453_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n760_), .A2(new_n764_), .ZN(G1332gat));
  OAI21_X1  g564(.A(G64gat), .B1(new_n763_), .B2(new_n337_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT48), .Z(new_n767_));
  NOR3_X1   g566(.A1(new_n758_), .A2(G64gat), .A3(new_n337_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT110), .ZN(G1333gat));
  OAI21_X1  g569(.A(G71gat), .B1(new_n763_), .B2(new_n513_), .ZN(new_n771_));
  XOR2_X1   g570(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n513_), .A2(G71gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n758_), .B2(new_n774_), .ZN(G1334gat));
  OAI21_X1  g574(.A(G78gat), .B1(new_n763_), .B2(new_n472_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT50), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n472_), .A2(G78gat), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT112), .Z(new_n779_));
  OAI21_X1  g578(.A(new_n777_), .B1(new_n758_), .B2(new_n779_), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n695_), .A2(new_n610_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n756_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n566_), .A3(new_n659_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n761_), .A2(new_n655_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n736_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n659_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n787_), .B2(new_n566_), .ZN(G1336gat));
  NAND3_X1  g587(.A1(new_n782_), .A2(new_n567_), .A3(new_n728_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n728_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n789_), .B1(new_n791_), .B2(new_n567_), .ZN(G1337gat));
  NAND3_X1  g591(.A1(new_n736_), .A2(new_n501_), .A3(new_n784_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(G99gat), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n782_), .A2(new_n501_), .A3(new_n563_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT113), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n797_), .A2(KEYINPUT51), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n796_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n800_), .A2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n797_), .A2(new_n801_), .A3(KEYINPUT51), .A4(new_n799_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1338gat));
  NAND2_X1  g605(.A1(new_n785_), .A2(new_n690_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n782_), .A2(new_n564_), .A3(new_n690_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT115), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT52), .B1(new_n807_), .B2(G106gat), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(G1339gat));
  INV_X1    g614(.A(new_n639_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n604_), .A2(new_n608_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n554_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n592_), .A2(new_n595_), .A3(KEYINPUT55), .A4(new_n598_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n600_), .A2(KEYINPUT118), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n599_), .B(new_n819_), .C1(new_n822_), .C2(new_n820_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n821_), .A2(new_n823_), .A3(KEYINPUT119), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT119), .B1(new_n821_), .B2(new_n823_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n608_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT56), .B(new_n608_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n818_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n542_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n546_), .A2(new_n831_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n538_), .A2(new_n541_), .A3(new_n831_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n552_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n547_), .A2(new_n551_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n609_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n816_), .B1(new_n830_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT57), .B(new_n816_), .C1(new_n830_), .C2(new_n837_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n826_), .A2(KEYINPUT120), .A3(new_n827_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n817_), .A2(new_n836_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n828_), .A2(new_n846_), .A3(new_n829_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(KEYINPUT58), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n640_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT58), .B1(new_n845_), .B2(new_n847_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n840_), .B(new_n841_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n656_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n714_), .A2(new_n610_), .A3(new_n655_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n554_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n657_), .A2(KEYINPUT117), .A3(new_n669_), .A4(new_n610_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n856_), .A3(KEYINPUT54), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n853_), .B(new_n858_), .C1(new_n854_), .C2(new_n554_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n852_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n510_), .A2(new_n513_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n659_), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n420_), .A3(new_n554_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n860_), .B1(new_n851_), .B2(new_n656_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n453_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(KEYINPUT59), .A3(new_n863_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n669_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n866_), .B1(new_n872_), .B2(new_n420_), .ZN(G1340gat));
  OAI21_X1  g672(.A(new_n418_), .B1(new_n610_), .B2(KEYINPUT60), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n418_), .A2(KEYINPUT60), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(KEYINPUT121), .B2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n865_), .B(new_n876_), .C1(KEYINPUT121), .C2(new_n874_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n610_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n418_), .ZN(G1341gat));
  AOI21_X1  g678(.A(G127gat), .B1(new_n865_), .B2(new_n655_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n868_), .A2(new_n871_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT122), .B(G127gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n655_), .A2(new_n882_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT123), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n880_), .B1(new_n881_), .B2(new_n884_), .ZN(G1342gat));
  NAND3_X1  g684(.A1(new_n865_), .A2(new_n413_), .A3(new_n639_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n714_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n413_), .ZN(G1343gat));
  NOR3_X1   g687(.A1(new_n728_), .A2(new_n501_), .A3(new_n472_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n870_), .A2(new_n554_), .A3(new_n889_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g690(.A1(new_n870_), .A2(new_n668_), .A3(new_n889_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g692(.A1(new_n870_), .A2(new_n655_), .A3(new_n889_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1346gat));
  AND4_X1   g695(.A1(G162gat), .A2(new_n870_), .A3(new_n640_), .A4(new_n889_), .ZN(new_n897_));
  AND4_X1   g696(.A1(new_n659_), .A2(new_n862_), .A3(new_n639_), .A4(new_n889_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT124), .B1(new_n898_), .B2(G162gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n870_), .A2(new_n639_), .A3(new_n889_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n901_));
  INV_X1    g700(.A(G162gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n897_), .B1(new_n899_), .B2(new_n903_), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n507_), .A2(new_n690_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NOR4_X1   g705(.A1(new_n869_), .A2(new_n337_), .A3(new_n669_), .A4(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT22), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n223_), .B1(new_n907_), .B2(new_n911_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n910_), .B1(new_n912_), .B2(new_n913_), .ZN(G1348gat));
  NOR2_X1   g713(.A1(new_n869_), .A2(new_n337_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n915_), .A2(new_n668_), .A3(new_n905_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g716(.A1(new_n915_), .A2(new_n655_), .A3(new_n905_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n291_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n919_), .B1(new_n209_), .B2(new_n918_), .ZN(G1350gat));
  NAND2_X1  g719(.A1(new_n639_), .A2(new_n226_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(KEYINPUT125), .Z(new_n922_));
  NAND3_X1  g721(.A1(new_n915_), .A2(new_n905_), .A3(new_n922_), .ZN(new_n923_));
  NOR4_X1   g722(.A1(new_n869_), .A2(new_n337_), .A3(new_n714_), .A4(new_n906_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n924_), .B2(new_n210_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(KEYINPUT126), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n923_), .B(new_n927_), .C1(new_n210_), .C2(new_n924_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1351gat));
  AND2_X1   g728(.A1(new_n513_), .A2(new_n454_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n915_), .A2(new_n554_), .A3(new_n930_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G197gat), .ZN(G1352gat));
  AND4_X1   g731(.A1(new_n278_), .A2(new_n915_), .A3(new_n668_), .A4(new_n930_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n915_), .A2(new_n668_), .A3(new_n930_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n252_), .B2(new_n934_), .ZN(G1353gat));
  AND2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  AOI211_X1 g736(.A(new_n936_), .B(new_n656_), .C1(KEYINPUT127), .C2(new_n937_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n915_), .A2(new_n930_), .A3(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n937_), .A2(KEYINPUT127), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n939_), .B(new_n940_), .ZN(G1354gat));
  NAND2_X1  g740(.A1(new_n915_), .A2(new_n930_), .ZN(new_n942_));
  OAI21_X1  g741(.A(G218gat), .B1(new_n942_), .B2(new_n714_), .ZN(new_n943_));
  OR2_X1    g742(.A1(new_n816_), .A2(G218gat), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n942_), .B2(new_n944_), .ZN(G1355gat));
endmodule


