//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n580_, new_n581_, new_n582_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  AOI22_X1  g004(.A1(new_n205_), .A2(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n206_));
  INV_X1    g005(.A(G183gat), .ZN(new_n207_));
  INV_X1    g006(.A(G190gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT23), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT82), .Z(new_n210_));
  NOR3_X1   g009(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT23), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  OAI221_X1 g012(.A(new_n206_), .B1(KEYINPUT81), .B2(new_n205_), .C1(new_n212_), .C2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(KEYINPUT24), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT79), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT25), .B(G183gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n215_), .A2(KEYINPUT79), .A3(KEYINPUT24), .A4(new_n216_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n219_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT80), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n225_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n209_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(new_n211_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n215_), .A2(KEYINPUT24), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n226_), .A2(new_n227_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n214_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G204gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G197gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT85), .B(G197gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n235_), .B1(new_n236_), .B2(new_n234_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G211gat), .B(G218gat), .Z(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(KEYINPUT21), .A3(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n237_), .A2(KEYINPUT21), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT21), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n241_), .B1(G197gat), .B2(G204gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n236_), .B2(G204gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n238_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n239_), .B1(new_n240_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n233_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G226gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT19), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n222_), .A2(new_n217_), .A3(new_n231_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n203_), .B(KEYINPUT89), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(G176gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n216_), .B(KEYINPUT88), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n229_), .B2(new_n213_), .ZN(new_n255_));
  OAI22_X1  g054(.A1(new_n212_), .A2(new_n251_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT20), .B1(new_n256_), .B2(new_n246_), .ZN(new_n257_));
  OR3_X1    g056(.A1(new_n248_), .A2(new_n250_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n233_), .A2(new_n247_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n246_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT20), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(new_n250_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n202_), .B1(new_n258_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G8gat), .B(G36gat), .ZN(new_n265_));
  INV_X1    g064(.A(G92gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT18), .B(G64gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n262_), .A2(new_n202_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n264_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n271_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n269_), .B1(new_n273_), .B2(new_n263_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT27), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n250_), .B1(new_n248_), .B2(new_n257_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n250_), .B2(new_n261_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n276_), .B1(new_n278_), .B2(new_n269_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n275_), .A2(new_n276_), .B1(new_n272_), .B2(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(G141gat), .A2(G148gat), .ZN(new_n284_));
  OR2_X1    g083(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT2), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n284_), .A2(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n288_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n290_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n283_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT84), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n281_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n282_), .B1(new_n295_), .B2(KEYINPUT1), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n296_), .B1(KEYINPUT1), .B2(new_n295_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n297_), .A2(new_n284_), .A3(new_n287_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n294_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G113gat), .B(G120gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(G127gat), .B(G134gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n299_), .B(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT4), .ZN(new_n304_));
  INV_X1    g103(.A(new_n299_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(new_n306_), .A3(new_n302_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n308_), .B(KEYINPUT91), .Z(new_n309_));
  NAND3_X1  g108(.A1(new_n304_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n303_), .A2(new_n308_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G57gat), .B(G85gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(G1gat), .B(G29gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(KEYINPUT92), .B(KEYINPUT0), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n310_), .A2(new_n311_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n316_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n246_), .B1(new_n299_), .B2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G78gat), .B(G106gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(G228gat), .B(G233gat), .C1(new_n247_), .C2(KEYINPUT86), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT87), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n299_), .A2(new_n320_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT28), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G22gat), .B(G50gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n327_), .B(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n333_), .A2(new_n329_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n326_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n329_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n328_), .A2(new_n330_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(KEYINPUT87), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n325_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT87), .B1(new_n336_), .B2(new_n337_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n323_), .A2(new_n324_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n323_), .A2(new_n324_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G71gat), .B(G99gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(G43gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n233_), .B(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G227gat), .A2(G233gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n302_), .B(new_n348_), .Z(new_n349_));
  XOR2_X1   g148(.A(KEYINPUT30), .B(G15gat), .Z(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT31), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n349_), .B(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n347_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n347_), .A2(new_n352_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n280_), .A2(new_n319_), .A3(new_n344_), .A4(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n270_), .A2(KEYINPUT32), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n264_), .A2(new_n358_), .A3(new_n271_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n278_), .A2(KEYINPUT32), .A3(new_n270_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n359_), .B(new_n360_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n310_), .A2(new_n311_), .A3(new_n316_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n310_), .A2(KEYINPUT33), .A3(new_n311_), .A4(new_n316_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n304_), .A2(new_n308_), .A3(new_n307_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n316_), .B1(new_n303_), .B2(new_n309_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n364_), .A2(new_n365_), .A3(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n361_), .B1(new_n369_), .B2(new_n275_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n339_), .A2(new_n319_), .A3(new_n343_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n370_), .A2(new_n344_), .B1(new_n371_), .B2(new_n280_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n357_), .B1(new_n372_), .B2(new_n356_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G57gat), .B(G64gat), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n374_), .A2(KEYINPUT11), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(KEYINPUT11), .ZN(new_n376_));
  XOR2_X1   g175(.A(G71gat), .B(G78gat), .Z(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n376_), .A2(new_n377_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G85gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n266_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G85gat), .A2(G92gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(KEYINPUT8), .ZN(new_n385_));
  AND2_X1   g184(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n386_));
  NOR2_X1   g185(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n387_));
  OAI22_X1  g186(.A1(new_n386_), .A2(new_n387_), .B1(G99gat), .B2(G106gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(G99gat), .A2(G106gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  AND3_X1   g191(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n385_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT67), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT67), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n399_), .B(new_n385_), .C1(new_n392_), .C2(new_n396_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n396_), .B1(new_n392_), .B2(KEYINPUT68), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT68), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n388_), .A2(new_n402_), .A3(new_n391_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n384_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT8), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n398_), .B(new_n400_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT65), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT9), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n408_), .A2(KEYINPUT64), .ZN(new_n409_));
  AND2_X1   g208(.A1(G85gat), .A2(G92gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT10), .B(G99gat), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n395_), .B(new_n411_), .C1(G106gat), .C2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n408_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT64), .B1(new_n410_), .B2(KEYINPUT9), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n407_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(G99gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT10), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT10), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G99gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(G106gat), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n422_), .A2(new_n423_), .B1(new_n410_), .B2(new_n409_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G85gat), .A2(G92gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT9), .B1(new_n410_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n383_), .A2(new_n408_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(KEYINPUT64), .A3(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n424_), .A2(new_n428_), .A3(KEYINPUT65), .A4(new_n395_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n417_), .A2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT69), .B1(new_n406_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n398_), .A2(new_n400_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT66), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT7), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n389_), .B1(new_n435_), .B2(new_n390_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n389_), .A2(new_n390_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT68), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(new_n403_), .A3(new_n395_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n384_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n405_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n430_), .B(KEYINPUT69), .C1(new_n432_), .C2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n380_), .B1(new_n431_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n430_), .B1(new_n432_), .B2(new_n441_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT69), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n380_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n442_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G230gat), .A2(G233gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT12), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n380_), .A2(new_n454_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n445_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n455_), .A2(new_n451_), .A3(new_n444_), .A4(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n453_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G120gat), .B(G148gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(new_n234_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT5), .B(G176gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n462_), .B(new_n463_), .Z(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n453_), .A2(new_n459_), .A3(new_n464_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n469_), .A2(KEYINPUT13), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(KEYINPUT13), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G15gat), .B(G22gat), .ZN(new_n474_));
  INV_X1    g273(.A(G1gat), .ZN(new_n475_));
  INV_X1    g274(.A(G8gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT14), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G1gat), .B(G8gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G43gat), .B(G50gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(G29gat), .B(G36gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n480_), .B(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(G229gat), .A3(G233gat), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n485_), .A2(KEYINPUT75), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(KEYINPUT75), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n480_), .A2(new_n483_), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n483_), .B(KEYINPUT15), .Z(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n489_), .B2(new_n480_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G229gat), .A2(G233gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT76), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n486_), .A2(new_n487_), .A3(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G113gat), .B(G141gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G169gat), .B(G197gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n495_), .B(new_n500_), .Z(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n473_), .A2(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n373_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G190gat), .B(G218gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G134gat), .B(G162gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n505_), .B(new_n506_), .Z(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT36), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n447_), .A2(new_n442_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n510_), .A2(new_n483_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT35), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT34), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n445_), .A2(new_n489_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n515_), .A2(new_n512_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n517_), .A2(new_n518_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n508_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n517_), .A2(new_n518_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n507_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT36), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n525_), .A3(new_n519_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT37), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n527_), .A2(KEYINPUT70), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n522_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(KEYINPUT70), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT71), .Z(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n380_), .B(new_n480_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G231gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n536_), .A2(KEYINPUT72), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G127gat), .B(G155gat), .ZN(new_n538_));
  INV_X1    g337(.A(G211gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT16), .B(G183gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT17), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n537_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n537_), .A2(new_n544_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n542_), .A2(KEYINPUT17), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n536_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n545_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT73), .Z(new_n550_));
  NAND4_X1  g349(.A1(new_n522_), .A2(new_n526_), .A3(new_n528_), .A4(new_n531_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n533_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n552_), .B(KEYINPUT74), .Z(new_n553_));
  NAND2_X1  g352(.A1(new_n504_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n319_), .B(KEYINPUT93), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n475_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT38), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n550_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n522_), .A2(new_n526_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n504_), .A2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(G1gat), .B1(new_n563_), .B2(new_n319_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n557_), .A2(new_n558_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n559_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT94), .Z(G1324gat));
  INV_X1    g366(.A(new_n280_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n555_), .A2(new_n476_), .A3(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(G8gat), .B1(new_n563_), .B2(new_n280_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n570_), .A2(KEYINPUT39), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(KEYINPUT39), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n569_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g373(.A(G15gat), .B1(new_n563_), .B2(new_n355_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT41), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(KEYINPUT41), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n554_), .A2(G15gat), .A3(new_n355_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(G1326gat));
  OAI21_X1  g378(.A(G22gat), .B1(new_n563_), .B2(new_n344_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT42), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n344_), .A2(G22gat), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n581_), .B1(new_n554_), .B2(new_n582_), .ZN(G1327gat));
  AND2_X1   g382(.A1(new_n560_), .A2(new_n561_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n504_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT97), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n504_), .A2(KEYINPUT97), .A3(new_n584_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n319_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(G29gat), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n533_), .A2(new_n551_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n370_), .A2(new_n344_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n371_), .A2(new_n280_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n356_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n357_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n594_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT43), .B1(new_n593_), .B2(KEYINPUT95), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n373_), .A2(KEYINPUT95), .A3(KEYINPUT43), .A4(new_n594_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n601_), .A2(new_n602_), .A3(new_n503_), .A4(new_n560_), .ZN(new_n603_));
  XOR2_X1   g402(.A(KEYINPUT96), .B(KEYINPUT44), .Z(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n550_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(KEYINPUT96), .A2(KEYINPUT44), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n606_), .A2(new_n503_), .A3(new_n602_), .A4(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n556_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n592_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n591_), .A2(new_n592_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT98), .ZN(G1328gat));
  NOR2_X1   g412(.A1(new_n280_), .A2(G36gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n587_), .A2(new_n588_), .A3(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT45), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n280_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT99), .ZN(new_n618_));
  OAI21_X1  g417(.A(G36gat), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  AOI211_X1 g418(.A(KEYINPUT99), .B(new_n280_), .C1(new_n605_), .C2(new_n608_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n616_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT46), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n616_), .B(KEYINPUT46), .C1(new_n619_), .C2(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1329gat));
  INV_X1    g424(.A(G43gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n589_), .A2(new_n626_), .A3(new_n356_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n355_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n627_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT47), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(G1330gat));
  INV_X1    g430(.A(G50gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n344_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n589_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n344_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n632_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1331gat));
  NOR2_X1   g437(.A1(new_n472_), .A2(new_n501_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n373_), .A2(new_n639_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n640_), .A2(new_n553_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G57gat), .B1(new_n641_), .B2(new_n556_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n562_), .ZN(new_n643_));
  INV_X1    g442(.A(G57gat), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n319_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n642_), .A2(new_n645_), .ZN(G1332gat));
  INV_X1    g445(.A(G64gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n641_), .A2(new_n647_), .A3(new_n568_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G64gat), .B1(new_n643_), .B2(new_n280_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(KEYINPUT48), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(KEYINPUT48), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n648_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT101), .ZN(G1333gat));
  OAI21_X1  g452(.A(G71gat), .B1(new_n643_), .B2(new_n355_), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT102), .B(KEYINPUT49), .Z(new_n655_));
  OR2_X1    g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n655_), .ZN(new_n657_));
  INV_X1    g456(.A(G71gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n641_), .A2(new_n658_), .A3(new_n356_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n656_), .A2(new_n657_), .A3(new_n659_), .ZN(G1334gat));
  OAI21_X1  g459(.A(G78gat), .B1(new_n643_), .B2(new_n344_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT50), .ZN(new_n662_));
  INV_X1    g461(.A(G78gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n641_), .A2(new_n663_), .A3(new_n633_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1335gat));
  NAND3_X1  g464(.A1(new_n606_), .A2(new_n602_), .A3(new_n639_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n666_), .A2(KEYINPUT103), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(KEYINPUT103), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n590_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G85gat), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n640_), .A2(new_n584_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n381_), .A3(new_n556_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n670_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT104), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n670_), .A2(new_n676_), .A3(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1336gat));
  AOI21_X1  g477(.A(G92gat), .B1(new_n672_), .B2(new_n568_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n667_), .A2(new_n668_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n280_), .A2(new_n266_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n680_), .B2(new_n681_), .ZN(G1337gat));
  NAND3_X1  g481(.A1(new_n667_), .A2(new_n356_), .A3(new_n668_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G99gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n672_), .A2(new_n422_), .A3(new_n356_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT51), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT51), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n684_), .A2(new_n688_), .A3(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1338gat));
  NAND3_X1  g489(.A1(new_n672_), .A2(new_n423_), .A3(new_n633_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n666_), .A2(new_n344_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT52), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(G106gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n692_), .B2(G106gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT105), .B(KEYINPUT53), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n691_), .B(new_n697_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1339gat));
  NAND2_X1  g500(.A1(new_n472_), .A2(new_n502_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(new_n552_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT54), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT54), .B1(new_n702_), .B2(new_n552_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n704_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n501_), .A2(new_n467_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n452_), .A2(KEYINPUT55), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n457_), .B1(new_n509_), .B2(new_n380_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n455_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n452_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n712_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n713_), .A2(new_n455_), .A3(new_n715_), .A4(new_n452_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT55), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n459_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n459_), .A2(new_n721_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT107), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(new_n722_), .A3(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(KEYINPUT56), .A3(new_n465_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT56), .B1(new_n725_), .B2(new_n465_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(KEYINPUT109), .ZN(new_n728_));
  AOI22_X1  g527(.A1(new_n718_), .A2(new_n717_), .B1(new_n723_), .B2(KEYINPUT107), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n464_), .B1(new_n729_), .B2(new_n722_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n730_), .A2(new_n731_), .A3(KEYINPUT56), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n711_), .B1(new_n728_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n495_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n493_), .B1(new_n490_), .B2(KEYINPUT110), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n735_), .B1(KEYINPUT110), .B2(new_n490_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n500_), .B1(new_n484_), .B2(new_n493_), .ZN(new_n737_));
  AOI22_X1  g536(.A1(new_n734_), .A2(new_n500_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n468_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n561_), .B1(new_n733_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT57), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT57), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n731_), .B1(new_n730_), .B2(KEYINPUT56), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n725_), .A2(new_n465_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(KEYINPUT109), .A3(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(new_n748_), .A3(new_n726_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n739_), .B1(new_n749_), .B2(new_n711_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT111), .B(new_n744_), .C1(new_n750_), .C2(new_n561_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n727_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n726_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n738_), .A2(new_n467_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n727_), .B2(KEYINPUT112), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT58), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n593_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n754_), .A2(KEYINPUT58), .A3(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n743_), .A2(new_n751_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n560_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n710_), .A2(new_n763_), .ZN(new_n764_));
  NOR4_X1   g563(.A1(new_n610_), .A2(new_n633_), .A3(new_n568_), .A4(new_n355_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT113), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G113gat), .B1(new_n768_), .B2(new_n501_), .ZN(new_n769_));
  XOR2_X1   g568(.A(KEYINPUT114), .B(KEYINPUT59), .Z(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n767_), .B1(new_n772_), .B2(KEYINPUT59), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n502_), .A2(KEYINPUT115), .ZN(new_n776_));
  MUX2_X1   g575(.A(KEYINPUT115), .B(new_n776_), .S(G113gat), .Z(new_n777_));
  AOI21_X1  g576(.A(new_n769_), .B1(new_n775_), .B2(new_n777_), .ZN(G1340gat));
  XOR2_X1   g577(.A(KEYINPUT116), .B(G120gat), .Z(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n774_), .B2(new_n472_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT60), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n472_), .B2(new_n779_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n768_), .B(new_n782_), .C1(new_n781_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n783_), .ZN(G1341gat));
  INV_X1    g583(.A(G127gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n767_), .B2(new_n560_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n771_), .A2(new_n773_), .A3(G127gat), .A4(new_n550_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n787_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n788_), .A2(new_n789_), .A3(new_n790_), .ZN(G1342gat));
  AOI21_X1  g590(.A(G134gat), .B1(new_n768_), .B2(new_n561_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n594_), .A2(G134gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n775_), .B2(new_n793_), .ZN(G1343gat));
  OAI21_X1  g593(.A(KEYINPUT111), .B1(new_n750_), .B2(new_n561_), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n795_), .A2(KEYINPUT57), .B1(new_n760_), .B2(new_n759_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n550_), .B1(new_n796_), .B2(new_n751_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n708_), .A2(new_n709_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n556_), .A2(new_n633_), .A3(new_n280_), .A4(new_n355_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n501_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n473_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g604(.A(KEYINPUT61), .B(G155gat), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n801_), .A2(new_n808_), .A3(new_n550_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n801_), .B2(new_n550_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n807_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n811_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(new_n809_), .A3(new_n806_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1346gat));
  INV_X1    g614(.A(G162gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n801_), .A2(new_n816_), .A3(new_n561_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n799_), .A2(new_n593_), .A3(new_n800_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n816_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT119), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n817_), .B(new_n821_), .C1(new_n816_), .C2(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(G1347gat));
  NOR3_X1   g622(.A1(new_n556_), .A2(new_n280_), .A3(new_n355_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n344_), .B(new_n824_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT120), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n764_), .A2(new_n827_), .A3(new_n344_), .A4(new_n824_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n252_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n501_), .A3(new_n830_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n825_), .A2(new_n502_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT62), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n832_), .A2(new_n833_), .A3(G169gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(G169gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(G1348gat));
  NAND2_X1  g635(.A1(new_n764_), .A2(new_n344_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT121), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n764_), .A2(new_n839_), .A3(new_n344_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n472_), .A2(new_n204_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n838_), .A2(new_n840_), .A3(new_n824_), .A4(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT122), .ZN(new_n843_));
  INV_X1    g642(.A(new_n824_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n837_), .B2(KEYINPUT121), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n840_), .A4(new_n841_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n826_), .A2(new_n473_), .A3(new_n828_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n204_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n843_), .A2(new_n847_), .A3(new_n849_), .ZN(G1349gat));
  NAND3_X1  g649(.A1(new_n845_), .A2(new_n550_), .A3(new_n840_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n560_), .A2(new_n220_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n851_), .A2(new_n207_), .B1(new_n829_), .B2(new_n852_), .ZN(G1350gat));
  NAND3_X1  g652(.A1(new_n829_), .A2(new_n221_), .A3(new_n561_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n826_), .A2(new_n594_), .A3(new_n828_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n855_), .A2(new_n856_), .A3(G190gat), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n855_), .B2(G190gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n854_), .B1(new_n857_), .B2(new_n858_), .ZN(G1351gat));
  NOR4_X1   g658(.A1(new_n280_), .A2(new_n344_), .A3(new_n590_), .A4(new_n356_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n764_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n501_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g663(.A1(new_n861_), .A2(new_n472_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  XOR2_X1   g666(.A(KEYINPUT124), .B(G204gat), .Z(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n865_), .B2(new_n868_), .ZN(G1353gat));
  INV_X1    g668(.A(KEYINPUT63), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT126), .B1(new_n870_), .B2(new_n539_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n550_), .B1(new_n870_), .B2(new_n539_), .ZN(new_n872_));
  XOR2_X1   g671(.A(new_n872_), .B(KEYINPUT125), .Z(new_n873_));
  AOI21_X1  g672(.A(new_n871_), .B1(new_n862_), .B2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n870_), .A2(new_n539_), .A3(KEYINPUT126), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1354gat));
  INV_X1    g675(.A(G218gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n862_), .A2(new_n877_), .A3(new_n561_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT127), .ZN(new_n879_));
  OAI21_X1  g678(.A(G218gat), .B1(new_n861_), .B2(new_n593_), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n878_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1355gat));
endmodule


