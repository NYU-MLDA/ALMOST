//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT13), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G120gat), .B(G148gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(G204gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT5), .B(G176gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT69), .Z(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n211_), .B(KEYINPUT6), .Z(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT10), .B(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n212_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G92gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(G85gat), .B1(new_n217_), .B2(KEYINPUT9), .ZN(new_n218_));
  NAND2_X1  g017(.A1(KEYINPUT9), .A2(G92gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n221_));
  XOR2_X1   g020(.A(new_n221_), .B(KEYINPUT65), .Z(new_n222_));
  OAI21_X1  g021(.A(new_n216_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G85gat), .B(G92gat), .Z(new_n224_));
  INV_X1    g023(.A(G99gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n213_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT7), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n224_), .B1(new_n227_), .B2(new_n212_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT8), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n223_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(KEYINPUT8), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n227_), .A2(KEYINPUT66), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n212_), .B1(new_n227_), .B2(KEYINPUT66), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G57gat), .B(G64gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT11), .ZN(new_n241_));
  XOR2_X1   g040(.A(G71gat), .B(G78gat), .Z(new_n242_));
  OR2_X1    g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n238_), .B(KEYINPUT67), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n241_), .A2(new_n246_), .A3(new_n242_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n243_), .A2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n237_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT12), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n237_), .A2(new_n248_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G230gat), .A2(G233gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n231_), .A2(new_n254_), .A3(new_n236_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n223_), .A2(new_n230_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT68), .B1(new_n256_), .B2(new_n235_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(KEYINPUT12), .A3(new_n248_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n252_), .A2(new_n253_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n249_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n253_), .B1(new_n262_), .B2(new_n251_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n210_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n265_));
  INV_X1    g064(.A(new_n263_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n260_), .A2(new_n266_), .A3(new_n209_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n265_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n204_), .B(new_n205_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n264_), .A2(new_n267_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT70), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n272_), .A2(new_n202_), .A3(new_n273_), .A4(new_n203_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G15gat), .B(G22gat), .ZN(new_n277_));
  INV_X1    g076(.A(G1gat), .ZN(new_n278_));
  INV_X1    g077(.A(G8gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT14), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G1gat), .B(G8gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G43gat), .B(G50gat), .Z(new_n284_));
  XNOR2_X1  g083(.A(G29gat), .B(G36gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(KEYINPUT15), .Z(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(new_n283_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G229gat), .A2(G233gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n283_), .B(new_n286_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n290_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G113gat), .B(G141gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G169gat), .B(G197gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(KEYINPUT79), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n295_), .B(new_n300_), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n276_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G228gat), .A2(G233gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n303_), .B(KEYINPUT88), .Z(new_n304_));
  INV_X1    g103(.A(KEYINPUT90), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308_));
  INV_X1    g107(.A(G141gat), .ZN(new_n309_));
  INV_X1    g108(.A(G148gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(KEYINPUT3), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  AND2_X1   g114(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n316_));
  NOR2_X1   g115(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(G141gat), .B(G148gat), .C1(KEYINPUT85), .C2(KEYINPUT2), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n314_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT86), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT86), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n314_), .A2(new_n318_), .A3(new_n322_), .A4(new_n319_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT87), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT87), .B1(new_n329_), .B2(new_n324_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n321_), .A2(new_n323_), .A3(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT84), .B1(new_n327_), .B2(KEYINPUT1), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT84), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT1), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(G155gat), .A4(G162gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n327_), .A2(KEYINPUT1), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n334_), .A2(new_n337_), .A3(new_n338_), .A4(new_n325_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n309_), .A2(new_n310_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n339_), .A2(new_n340_), .A3(new_n315_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n308_), .B1(new_n333_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT21), .ZN(new_n344_));
  INV_X1    g143(.A(G197gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT89), .ZN(new_n347_));
  INV_X1    g146(.A(G204gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n347_), .B1(G197gat), .B2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(G197gat), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n344_), .B(new_n346_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G211gat), .B(G218gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n345_), .A2(G204gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(G197gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT21), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n351_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n352_), .A2(new_n344_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n346_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(new_n305_), .B2(new_n304_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n307_), .B1(new_n343_), .B2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G78gat), .B(G106gat), .Z(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G211gat), .B(G218gat), .Z(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(KEYINPUT21), .B2(new_n355_), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n367_), .A2(new_n351_), .B1(new_n359_), .B2(new_n358_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n304_), .A2(new_n305_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n331_), .B1(new_n320_), .B2(KEYINPUT86), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n341_), .B1(new_n371_), .B2(new_n323_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n370_), .B(new_n306_), .C1(new_n372_), .C2(new_n308_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n363_), .A2(new_n365_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n365_), .B1(new_n363_), .B2(new_n373_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G22gat), .B(G50gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT28), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n372_), .A2(new_n379_), .A3(new_n308_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n372_), .B2(new_n308_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n378_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n382_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(new_n380_), .A3(new_n377_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n376_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT92), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n363_), .A2(new_n373_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n364_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n363_), .A2(new_n365_), .A3(new_n373_), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT91), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT91), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n385_), .B(new_n383_), .C1(new_n375_), .C2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n388_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(KEYINPUT91), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n396_), .A2(new_n386_), .A3(new_n397_), .A4(KEYINPUT92), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n387_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT98), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT19), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G183gat), .A2(G190gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n406_), .A2(KEYINPUT23), .ZN(new_n407_));
  AND2_X1   g206(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n408_));
  NOR2_X1   g207(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n407_), .B1(new_n410_), .B2(new_n406_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(G169gat), .A2(G176gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(KEYINPUT24), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n405_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n413_), .A2(KEYINPUT24), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(G183gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT80), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT80), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G183gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n421_), .A3(KEYINPUT25), .ZN(new_n422_));
  NOR2_X1   g221(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G190gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT26), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT26), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(G190gat), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n417_), .B1(new_n425_), .B2(new_n430_), .ZN(new_n431_));
  OR2_X1    g230(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n432_));
  NAND2_X1  g231(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n406_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n407_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n414_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(KEYINPUT82), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n415_), .A2(new_n431_), .A3(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(KEYINPUT83), .A2(G176gat), .ZN(new_n440_));
  AND2_X1   g239(.A1(KEYINPUT83), .A2(G176gat), .ZN(new_n441_));
  AND2_X1   g240(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n443_));
  OAI22_X1  g242(.A1(new_n440_), .A2(new_n441_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n419_), .A2(new_n421_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(G190gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n406_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT23), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n432_), .A2(new_n433_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n450_), .B2(new_n447_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n416_), .B(new_n444_), .C1(new_n446_), .C2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n439_), .A2(new_n368_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT24), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT93), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT93), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT24), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n412_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n413_), .A2(new_n456_), .A3(new_n458_), .A4(new_n416_), .ZN(new_n461_));
  AND2_X1   g260(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n427_), .B(new_n429_), .C1(new_n462_), .C2(new_n423_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n460_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n434_), .A2(new_n435_), .B1(new_n418_), .B2(new_n426_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n444_), .A2(new_n416_), .ZN(new_n466_));
  OAI22_X1  g265(.A1(new_n464_), .A2(new_n451_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n454_), .B1(new_n467_), .B2(new_n361_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n404_), .B1(new_n453_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n439_), .A2(new_n452_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n361_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT20), .B1(new_n467_), .B2(new_n361_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n474_), .A3(new_n404_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G8gat), .B(G36gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(G92gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT18), .B(G64gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n470_), .A2(new_n475_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT27), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n368_), .B1(new_n439_), .B2(new_n452_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n403_), .B1(new_n483_), .B2(new_n473_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n453_), .A2(new_n468_), .A3(new_n404_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n480_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n401_), .B1(new_n482_), .B2(new_n486_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n483_), .A2(new_n473_), .A3(new_n403_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n479_), .B1(new_n488_), .B2(new_n469_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n481_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT27), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n486_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n493_), .A2(KEYINPUT98), .A3(new_n481_), .A4(KEYINPUT27), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n487_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n400_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G1gat), .B(G29gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(G85gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT0), .B(G57gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G225gat), .A2(G233gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n333_), .A2(new_n342_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT94), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G127gat), .B(G134gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G113gat), .B(G120gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n333_), .A2(new_n342_), .A3(new_n507_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(KEYINPUT4), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT4), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n503_), .A2(new_n504_), .A3(new_n512_), .A4(new_n508_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n502_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n502_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n503_), .A2(new_n508_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n516_), .B2(new_n510_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n501_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n372_), .A2(KEYINPUT94), .A3(new_n507_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n510_), .A2(KEYINPUT4), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n513_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n515_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n517_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n500_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n518_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G71gat), .B(G99gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G43gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n471_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G227gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n507_), .B(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT30), .B(G15gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT31), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n530_), .B(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n528_), .A2(new_n533_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n525_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n496_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT99), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n500_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n541_));
  AOI211_X1 g340(.A(new_n501_), .B(new_n517_), .C1(new_n521_), .C2(new_n515_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n543_), .A2(new_n487_), .A3(new_n492_), .A4(new_n494_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n399_), .A2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT95), .B1(new_n541_), .B2(KEYINPUT33), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n516_), .A2(new_n515_), .A3(new_n510_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n500_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT96), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT96), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n547_), .A2(new_n550_), .A3(new_n500_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n502_), .B(new_n513_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n490_), .B1(new_n549_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT33), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n518_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n541_), .A2(KEYINPUT33), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n546_), .A2(new_n554_), .A3(new_n557_), .A4(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n480_), .A2(KEYINPUT32), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n488_), .A2(new_n469_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n562_), .B2(new_n560_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n563_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT97), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n525_), .A2(KEYINPUT97), .A3(new_n563_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n559_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n545_), .B1(new_n399_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n536_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n540_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n564_), .A2(new_n565_), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT97), .B1(new_n525_), .B2(new_n563_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n400_), .B1(new_n574_), .B2(new_n559_), .ZN(new_n575_));
  OAI211_X1 g374(.A(KEYINPUT99), .B(new_n536_), .C1(new_n575_), .C2(new_n545_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n539_), .B1(new_n571_), .B2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n302_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT37), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n579_), .A2(KEYINPUT76), .ZN(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n581_));
  NAND2_X1  g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT35), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n288_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT73), .ZN(new_n588_));
  OAI22_X1  g387(.A1(new_n587_), .A2(new_n588_), .B1(new_n286_), .B2(new_n237_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n587_), .A2(new_n588_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n585_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT74), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT74), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n593_), .B(new_n585_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n589_), .A2(new_n590_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n583_), .B(KEYINPUT35), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n592_), .A2(new_n594_), .A3(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599_));
  INV_X1    g398(.A(G162gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT75), .B(G134gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n603_), .A2(new_n604_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n598_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n591_), .A2(KEYINPUT74), .B1(new_n595_), .B2(new_n596_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n608_), .A2(new_n604_), .A3(new_n603_), .A4(new_n594_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n580_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n609_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT76), .B(KEYINPUT37), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n610_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT77), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n283_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n248_), .B(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(G127gat), .B(G155gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(G211gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(KEYINPUT16), .B(G183gat), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n623_), .A2(KEYINPUT17), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(KEYINPUT17), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n619_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT78), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n619_), .A2(new_n624_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n629_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n615_), .A2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n578_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n278_), .A3(new_n525_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT100), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n637_), .A2(KEYINPUT38), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(KEYINPUT38), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n612_), .A2(new_n632_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n578_), .A2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT101), .Z(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n543_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n638_), .A2(new_n639_), .A3(new_n644_), .ZN(G1324gat));
  INV_X1    g444(.A(new_n495_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G8gat), .B1(new_n641_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT39), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n634_), .A2(new_n279_), .A3(new_n495_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(G1325gat));
  INV_X1    g451(.A(G15gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n642_), .B2(new_n570_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n655_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n634_), .A2(new_n653_), .A3(new_n570_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(G1326gat));
  INV_X1    g458(.A(G22gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n642_), .B2(new_n400_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT42), .Z(new_n662_));
  NAND3_X1  g461(.A1(new_n634_), .A2(new_n660_), .A3(new_n400_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1327gat));
  NOR2_X1   g463(.A1(new_n611_), .A2(new_n631_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n578_), .A2(new_n665_), .ZN(new_n666_));
  OR3_X1    g465(.A1(new_n666_), .A2(G29gat), .A3(new_n543_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n568_), .A2(new_n399_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n545_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT99), .B1(new_n670_), .B2(new_n536_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n569_), .A2(new_n540_), .A3(new_n570_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n538_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(new_n615_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n607_), .A2(new_n609_), .A3(new_n614_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n612_), .B2(new_n580_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n577_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n302_), .A2(new_n631_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT104), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n681_), .B(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n525_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n685_), .A2(KEYINPUT105), .A3(G29gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT105), .B1(new_n685_), .B2(G29gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n667_), .B1(new_n686_), .B2(new_n687_), .ZN(G1328gat));
  OR2_X1    g487(.A1(new_n646_), .A2(KEYINPUT106), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n646_), .A2(KEYINPUT106), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n666_), .A2(G36gat), .A3(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n684_), .A2(new_n495_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(G36gat), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT46), .ZN(G1329gat));
  NOR3_X1   g496(.A1(new_n666_), .A2(G43gat), .A3(new_n536_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n684_), .A2(new_n570_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(G43gat), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g500(.A1(new_n666_), .A2(G50gat), .A3(new_n399_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n684_), .A2(new_n400_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(G50gat), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(G1331gat));
  NOR3_X1   g505(.A1(new_n577_), .A2(new_n301_), .A3(new_n276_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(new_n633_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G57gat), .B1(new_n708_), .B2(new_n525_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n640_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT109), .Z(new_n711_));
  AND2_X1   g510(.A1(new_n525_), .A2(G57gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(G1332gat));
  INV_X1    g512(.A(G64gat), .ZN(new_n714_));
  INV_X1    g513(.A(new_n691_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n711_), .B2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT48), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n708_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1333gat));
  INV_X1    g518(.A(G71gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n708_), .A2(new_n720_), .A3(new_n570_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n711_), .B2(new_n570_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n722_), .A2(new_n723_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(G1334gat));
  INV_X1    g525(.A(G78gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n711_), .B2(new_n400_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT50), .Z(new_n729_));
  NAND3_X1  g528(.A1(new_n708_), .A2(new_n727_), .A3(new_n400_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1335gat));
  NAND2_X1  g530(.A1(new_n707_), .A2(new_n665_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n525_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735_));
  INV_X1    g534(.A(new_n301_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n275_), .A2(new_n736_), .A3(new_n632_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n275_), .A2(KEYINPUT111), .A3(new_n736_), .A4(new_n632_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n679_), .A2(new_n735_), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n735_), .B1(new_n679_), .B2(new_n741_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n525_), .A2(G85gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n734_), .B1(new_n744_), .B2(new_n745_), .ZN(G1336gat));
  AOI21_X1  g545(.A(G92gat), .B1(new_n733_), .B2(new_n495_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT113), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n715_), .A2(new_n217_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n744_), .B2(new_n749_), .ZN(G1337gat));
  NOR3_X1   g549(.A1(new_n742_), .A2(new_n743_), .A3(new_n536_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n570_), .A2(new_n215_), .ZN(new_n752_));
  OAI22_X1  g551(.A1(new_n751_), .A2(new_n225_), .B1(new_n732_), .B2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g553(.A1(new_n733_), .A2(new_n213_), .A3(new_n400_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n674_), .B1(new_n673_), .B2(new_n615_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n577_), .A2(KEYINPUT43), .A3(new_n677_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n400_), .B(new_n741_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n679_), .A2(KEYINPUT114), .A3(new_n400_), .A4(new_n741_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(G106gat), .A3(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(KEYINPUT115), .A3(KEYINPUT52), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n760_), .A2(new_n764_), .A3(G106gat), .A4(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT115), .B1(new_n762_), .B2(KEYINPUT52), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n755_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT53), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n770_), .B(new_n755_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1339gat));
  INV_X1    g571(.A(new_n210_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n253_), .B1(new_n252_), .B2(new_n259_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n260_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n252_), .A2(KEYINPUT55), .A3(new_n253_), .A4(new_n259_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  OR3_X1    g578(.A1(new_n778_), .A2(KEYINPUT119), .A3(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(KEYINPUT119), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n301_), .A2(new_n267_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT118), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n780_), .A2(new_n781_), .A3(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n289_), .A2(new_n293_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n292_), .A2(new_n290_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n299_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n299_), .B2(new_n295_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT120), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n272_), .A2(new_n273_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n784_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n611_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT57), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n267_), .B(new_n789_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n778_), .A2(new_n779_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n797_), .A2(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(KEYINPUT58), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n615_), .A3(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n791_), .A2(KEYINPUT57), .A3(new_n611_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n794_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n632_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n275_), .A2(new_n301_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(new_n631_), .A3(new_n677_), .ZN(new_n805_));
  XOR2_X1   g604(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(KEYINPUT117), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n806_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n633_), .A2(new_n808_), .A3(new_n804_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT117), .B1(new_n805_), .B2(new_n806_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n803_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n400_), .A2(new_n495_), .A3(new_n536_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n525_), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(G113gat), .B1(new_n815_), .B2(new_n301_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(KEYINPUT59), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n812_), .A2(new_n818_), .A3(new_n525_), .A4(new_n813_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n301_), .A2(G113gat), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n816_), .B1(new_n820_), .B2(new_n821_), .ZN(G1340gat));
  NAND3_X1  g621(.A1(new_n817_), .A2(new_n275_), .A3(new_n819_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(KEYINPUT121), .B(G120gat), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n824_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n276_), .B2(KEYINPUT60), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(KEYINPUT60), .B2(new_n826_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n825_), .B1(new_n814_), .B2(new_n828_), .ZN(G1341gat));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n632_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n817_), .A2(new_n819_), .A3(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n830_), .B1(new_n814_), .B2(new_n632_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n832_), .A2(KEYINPUT122), .A3(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1342gat));
  AOI21_X1  g637(.A(G134gat), .B1(new_n815_), .B2(new_n612_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n615_), .A2(G134gat), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n820_), .B2(new_n840_), .ZN(G1343gat));
  NOR2_X1   g640(.A1(new_n399_), .A2(new_n570_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n691_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n812_), .A2(new_n525_), .A3(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n736_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(new_n309_), .ZN(G1344gat));
  NOR2_X1   g645(.A1(new_n844_), .A2(new_n276_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT123), .B(G148gat), .Z(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1345gat));
  OR3_X1    g648(.A1(new_n844_), .A2(KEYINPUT124), .A3(new_n632_), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT124), .B1(new_n844_), .B2(new_n632_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT61), .B(G155gat), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1346gat));
  NOR3_X1   g654(.A1(new_n844_), .A2(new_n600_), .A3(new_n677_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n844_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n612_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n856_), .B1(new_n600_), .B2(new_n858_), .ZN(G1347gat));
  INV_X1    g658(.A(KEYINPUT62), .ZN(new_n860_));
  NOR4_X1   g659(.A1(new_n691_), .A2(new_n400_), .A3(new_n525_), .A4(new_n536_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n812_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n736_), .ZN(new_n863_));
  INV_X1    g662(.A(G169gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n860_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n443_), .B2(new_n442_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT62), .B(G169gat), .C1(new_n862_), .C2(new_n736_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .ZN(G1348gat));
  INV_X1    g667(.A(new_n862_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n869_), .A2(G176gat), .A3(new_n275_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n441_), .A2(new_n440_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n275_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n871_), .B2(new_n872_), .ZN(G1349gat));
  NOR2_X1   g672(.A1(new_n862_), .A2(new_n632_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n445_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n462_), .A2(new_n423_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n874_), .ZN(G1350gat));
  NAND3_X1  g676(.A1(new_n869_), .A2(new_n430_), .A3(new_n612_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n869_), .A2(new_n615_), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n879_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT125), .B1(new_n879_), .B2(G190gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n878_), .B1(new_n880_), .B2(new_n881_), .ZN(G1351gat));
  AND3_X1   g681(.A1(new_n842_), .A2(KEYINPUT126), .A3(new_n543_), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT126), .B1(new_n842_), .B2(new_n543_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n883_), .A2(new_n691_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n812_), .A2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n736_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n345_), .ZN(G1352gat));
  NOR2_X1   g687(.A1(new_n886_), .A2(new_n276_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT127), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n348_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT127), .B(G204gat), .Z(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n889_), .B2(new_n892_), .ZN(G1353gat));
  INV_X1    g692(.A(new_n886_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n631_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  AND2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n895_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n898_), .B1(new_n895_), .B2(new_n896_), .ZN(G1354gat));
  AND3_X1   g698(.A1(new_n894_), .A2(G218gat), .A3(new_n615_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G218gat), .B1(new_n894_), .B2(new_n612_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1355gat));
endmodule


