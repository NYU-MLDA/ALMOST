//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT96), .ZN(new_n206_));
  INV_X1    g005(.A(G197gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(G204gat), .ZN(new_n208_));
  INV_X1    g007(.A(G204gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(KEYINPUT96), .A3(G197gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT21), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n207_), .A2(G204gat), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .A4(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT97), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n209_), .A2(G197gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n211_), .B1(new_n216_), .B2(new_n212_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G211gat), .B(G218gat), .Z(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n208_), .A2(new_n212_), .A3(new_n210_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n218_), .A2(KEYINPUT21), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n215_), .A2(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT24), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT24), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n225_), .B1(new_n227_), .B2(new_n223_), .ZN(new_n228_));
  INV_X1    g027(.A(G190gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT26), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT26), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G190gat), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G183gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(KEYINPUT25), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(G183gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n228_), .B1(new_n233_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(KEYINPUT23), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT82), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n244_), .B1(G183gat), .B2(G190gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n240_), .A2(KEYINPUT82), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT23), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n239_), .A2(new_n243_), .A3(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n240_), .A2(KEYINPUT23), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n240_), .A2(KEYINPUT82), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n244_), .A2(G183gat), .A3(G190gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT23), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT83), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n251_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  AOI211_X1 g055(.A(KEYINPUT83), .B(KEYINPUT23), .C1(new_n252_), .C2(new_n253_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n250_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT98), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT22), .B(G169gat), .ZN(new_n260_));
  INV_X1    g059(.A(G176gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n226_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n258_), .A2(new_n259_), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n259_), .B1(new_n258_), .B2(new_n264_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n222_), .B(new_n248_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT19), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT20), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n247_), .A2(new_n243_), .A3(new_n250_), .ZN(new_n272_));
  INV_X1    g071(.A(G169gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT22), .ZN(new_n274_));
  AOI21_X1  g073(.A(G176gat), .B1(new_n274_), .B2(KEYINPUT84), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(KEYINPUT84), .B2(new_n260_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n272_), .A2(new_n226_), .A3(new_n276_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n230_), .B(new_n232_), .C1(new_n235_), .C2(KEYINPUT80), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT80), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n236_), .A2(G183gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n234_), .A2(KEYINPUT25), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n279_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT81), .B1(new_n278_), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT80), .B1(new_n235_), .B2(new_n237_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT81), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n279_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n233_), .A4(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n228_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n283_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n256_), .A2(new_n257_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n277_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n213_), .A2(new_n214_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n213_), .A2(new_n214_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n219_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n221_), .A2(new_n220_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n271_), .B1(new_n291_), .B2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n267_), .A2(new_n270_), .A3(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT20), .B1(new_n291_), .B2(new_n296_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n248_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n299_), .B1(new_n300_), .B2(new_n296_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n205_), .B(new_n298_), .C1(new_n301_), .C2(new_n270_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT99), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n276_), .A2(new_n226_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT23), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n305_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n306_), .A2(new_n242_), .A3(new_n249_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n283_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n251_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n305_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(KEYINPUT83), .ZN(new_n312_));
  INV_X1    g111(.A(new_n257_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n308_), .B1(new_n309_), .B2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n271_), .B1(new_n315_), .B2(new_n222_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n248_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n249_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT98), .B1(new_n318_), .B2(new_n263_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n258_), .A2(new_n259_), .A3(new_n264_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n317_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n316_), .B1(new_n321_), .B2(new_n222_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n269_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT99), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n205_), .A4(new_n298_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n298_), .B1(new_n301_), .B2(new_n270_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n205_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n303_), .A2(new_n325_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT33), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G1gat), .B(G29gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G85gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT0), .B(G57gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n336_));
  OR2_X1    g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT89), .B1(new_n335_), .B2(KEYINPUT1), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT90), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n335_), .A2(KEYINPUT1), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n335_), .A2(KEYINPUT1), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT89), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT90), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(new_n337_), .A4(new_n336_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n340_), .A2(new_n341_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G141gat), .ZN(new_n348_));
  INV_X1    g147(.A(G148gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354_));
  AND4_X1   g153(.A1(KEYINPUT91), .A2(new_n354_), .A3(new_n348_), .A4(new_n349_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G141gat), .A2(G148gat), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT91), .B1(new_n356_), .B2(new_n354_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT2), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(G141gat), .B2(G148gat), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n351_), .A2(KEYINPUT2), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n359_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT92), .B1(new_n358_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n351_), .A2(KEYINPUT2), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n360_), .A2(G141gat), .A3(G148gat), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n365_), .A2(new_n366_), .B1(new_n350_), .B2(KEYINPUT3), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT92), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n367_), .B(new_n368_), .C1(new_n357_), .C2(new_n355_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n337_), .A2(new_n335_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n364_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G127gat), .B(G134gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G113gat), .B(G120gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n353_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n373_), .A2(new_n374_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT87), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT87), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n373_), .A2(new_n374_), .A3(KEYINPUT86), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT86), .B1(new_n373_), .B2(new_n374_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n378_), .B(new_n380_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n353_), .B2(new_n372_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT4), .B1(new_n376_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n367_), .B1(new_n357_), .B2(new_n355_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n370_), .B1(new_n389_), .B2(KEYINPUT92), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n390_), .A2(new_n369_), .B1(new_n347_), .B2(new_n352_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n388_), .B1(new_n391_), .B2(new_n383_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n385_), .A2(new_n387_), .A3(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n386_), .B1(new_n376_), .B2(new_n384_), .ZN(new_n394_));
  AOI211_X1 g193(.A(new_n330_), .B(new_n334_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n394_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n334_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n376_), .A2(new_n384_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n334_), .B1(new_n399_), .B2(new_n386_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n387_), .B1(new_n385_), .B2(new_n392_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT33), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n395_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n404_), .B(new_n298_), .C1(new_n301_), .C2(new_n270_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT100), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n393_), .A2(new_n334_), .A3(new_n394_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n222_), .B(new_n248_), .C1(new_n318_), .C2(new_n263_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n297_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n269_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(new_n322_), .B2(new_n269_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n404_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n398_), .A2(new_n407_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n329_), .A2(new_n403_), .B1(new_n406_), .B2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n415_));
  NAND2_X1  g214(.A1(new_n353_), .A2(new_n372_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(KEYINPUT29), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT29), .ZN(new_n418_));
  INV_X1    g217(.A(new_n415_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n391_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G22gat), .B(G50gat), .Z(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n417_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n422_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n418_), .B1(new_n353_), .B2(new_n372_), .ZN(new_n427_));
  OAI21_X1  g226(.A(G78gat), .B1(new_n427_), .B2(new_n222_), .ZN(new_n428_));
  INV_X1    g227(.A(G78gat), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n429_), .B(new_n296_), .C1(new_n391_), .C2(new_n418_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n428_), .A2(new_n430_), .A3(G106gat), .ZN(new_n431_));
  AOI21_X1  g230(.A(G106gat), .B1(new_n428_), .B2(new_n430_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G228gat), .A2(G233gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT95), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n433_), .A2(KEYINPUT95), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n434_), .B(new_n435_), .C1(new_n222_), .C2(KEYINPUT94), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n431_), .A2(new_n432_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G106gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n416_), .A2(KEYINPUT29), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n429_), .B1(new_n440_), .B2(new_n296_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n427_), .A2(G78gat), .A3(new_n222_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n439_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n428_), .A2(new_n430_), .A3(G106gat), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n436_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n426_), .B1(new_n438_), .B2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n437_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n444_), .A3(new_n436_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(new_n425_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n303_), .A2(new_n325_), .A3(new_n328_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT27), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n302_), .A2(KEYINPUT27), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n205_), .B(KEYINPUT101), .Z(new_n455_));
  NAND2_X1  g254(.A1(new_n411_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n398_), .A2(new_n407_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n450_), .A2(new_n460_), .ZN(new_n461_));
  OAI22_X1  g260(.A1(new_n414_), .A2(new_n450_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G71gat), .B(G99gat), .ZN(new_n464_));
  INV_X1    g263(.A(G43gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT31), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G227gat), .A2(G233gat), .ZN(new_n469_));
  INV_X1    g268(.A(G15gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n291_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n471_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n277_), .B(new_n473_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n472_), .A2(new_n476_), .A3(new_n474_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n383_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n383_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n468_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n482_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n467_), .A3(new_n480_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n463_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n483_), .A2(new_n486_), .A3(KEYINPUT88), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n447_), .A2(new_n448_), .A3(new_n425_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n425_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n459_), .B1(new_n486_), .B2(new_n483_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n453_), .A4(new_n457_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT102), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n451_), .A2(new_n452_), .B1(new_n456_), .B2(new_n454_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT102), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(new_n494_), .A4(new_n495_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n462_), .A2(new_n491_), .B1(new_n497_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G99gat), .A2(G106gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT6), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(G99gat), .A3(G106gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT10), .B(G99gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT64), .ZN(new_n509_));
  OR2_X1    g308(.A1(G85gat), .A2(G92gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT9), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G85gat), .A2(G92gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n510_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  OAI221_X1 g312(.A(new_n506_), .B1(G106gat), .B2(new_n507_), .C1(new_n509_), .C2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT65), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n506_), .A2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT7), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n503_), .A2(new_n505_), .A3(KEYINPUT65), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n510_), .A2(new_n512_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n515_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n515_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n524_), .B1(new_n506_), .B2(new_n519_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n514_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT66), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G57gat), .B(G64gat), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n527_), .B1(new_n528_), .B2(KEYINPUT11), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n528_), .A2(KEYINPUT11), .ZN(new_n531_));
  XOR2_X1   g330(.A(G71gat), .B(G78gat), .Z(new_n532_));
  NAND3_X1  g331(.A1(new_n528_), .A2(new_n527_), .A3(KEYINPUT11), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .A4(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n532_), .B1(KEYINPUT11), .B2(new_n528_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n533_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n535_), .B1(new_n536_), .B2(new_n529_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n526_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT12), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT67), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n526_), .A2(new_n539_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT67), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n526_), .A2(new_n539_), .A3(new_n544_), .A4(KEYINPUT12), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n540_), .A2(new_n541_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n542_), .A2(new_n543_), .A3(new_n545_), .A4(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(G230gat), .A2(G233gat), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n543_), .A2(new_n540_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n548_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G120gat), .B(G148gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT69), .ZN(new_n554_));
  XOR2_X1   g353(.A(G176gat), .B(G204gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT70), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n554_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n552_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n549_), .A2(new_n551_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(KEYINPUT71), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n564_), .A2(KEYINPUT71), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n563_), .B1(new_n567_), .B2(new_n565_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G29gat), .B(G36gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G43gat), .B(G50gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT78), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G15gat), .B(G22gat), .ZN(new_n576_));
  INV_X1    g375(.A(G1gat), .ZN(new_n577_));
  INV_X1    g376(.A(G8gat), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT14), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G1gat), .B(G8gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n580_), .B(new_n581_), .Z(new_n582_));
  NAND2_X1  g381(.A1(new_n575_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n573_), .B(KEYINPUT15), .ZN(new_n584_));
  INV_X1    g383(.A(new_n582_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G229gat), .A2(G233gat), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  OR3_X1    g388(.A1(new_n587_), .A2(KEYINPUT79), .A3(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT79), .B1(new_n587_), .B2(new_n589_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n575_), .B(new_n582_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n589_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n590_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G169gat), .B(G197gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n590_), .A2(new_n591_), .A3(new_n593_), .A4(new_n597_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n582_), .B(KEYINPUT74), .Z(new_n602_));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(new_n538_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G183gat), .B(G211gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT76), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT77), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n607_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G127gat), .B(G155gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT17), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n612_), .A2(new_n613_), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n605_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n605_), .A2(new_n614_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n573_), .B(new_n514_), .C1(new_n523_), .C2(new_n525_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT34), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT35), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n526_), .A2(new_n584_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(KEYINPUT72), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(KEYINPUT72), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n620_), .B(new_n625_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n623_), .A2(new_n624_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(G190gat), .B(G218gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT73), .ZN(new_n633_));
  XOR2_X1   g432(.A(G134gat), .B(G162gat), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT36), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n629_), .A2(new_n630_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n631_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n635_), .B(new_n636_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n631_), .B2(new_n638_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT37), .B1(new_n640_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n642_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT37), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n645_), .A3(new_n639_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n619_), .A2(new_n647_), .ZN(new_n648_));
  NOR4_X1   g447(.A1(new_n501_), .A2(new_n570_), .A3(new_n601_), .A4(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(new_n577_), .A3(new_n459_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT103), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n640_), .A2(new_n642_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n501_), .A2(new_n655_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n570_), .A2(new_n601_), .A3(new_n618_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n460_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n653_), .A2(new_n654_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n653_), .A2(KEYINPUT104), .A3(new_n654_), .A4(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1324gat));
  NAND3_X1  g464(.A1(new_n649_), .A2(new_n578_), .A3(new_n458_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n658_), .A2(new_n667_), .A3(new_n458_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n668_), .A2(G8gat), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT39), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT105), .B1(new_n659_), .B2(new_n498_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n670_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n666_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT40), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  OAI211_X1 g475(.A(KEYINPUT40), .B(new_n666_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1325gat));
  AOI21_X1  g477(.A(new_n470_), .B1(new_n658_), .B2(new_n490_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT41), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n649_), .A2(new_n470_), .A3(new_n490_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1326gat));
  INV_X1    g481(.A(G22gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n658_), .B2(new_n450_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT42), .Z(new_n685_));
  NAND3_X1  g484(.A1(new_n649_), .A2(new_n683_), .A3(new_n450_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1327gat));
  NOR2_X1   g486(.A1(new_n458_), .A2(new_n461_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n329_), .A2(new_n403_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n406_), .A2(new_n413_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n450_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n491_), .B1(new_n688_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n497_), .A2(new_n500_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n601_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n655_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n619_), .A2(new_n696_), .ZN(new_n697_));
  AND4_X1   g496(.A1(new_n694_), .A2(new_n695_), .A3(new_n569_), .A4(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n459_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n569_), .A2(new_n695_), .A3(new_n618_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT43), .B1(new_n501_), .B2(new_n647_), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT43), .B(new_n647_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  INV_X1    g505(.A(new_n647_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n694_), .A2(new_n704_), .A3(new_n706_), .A4(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT44), .B(new_n701_), .C1(new_n705_), .C2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT107), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n694_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT106), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n708_), .A3(new_n702_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(KEYINPUT44), .A4(new_n701_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n711_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n701_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n717_), .A2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n459_), .A2(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n699_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  INV_X1    g522(.A(G36gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n698_), .A2(new_n724_), .A3(new_n458_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT45), .Z(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n706_), .B1(new_n694_), .B2(new_n707_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(KEYINPUT106), .B2(new_n712_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n700_), .B1(new_n730_), .B2(new_n708_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n458_), .B1(new_n731_), .B2(KEYINPUT44), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n711_), .B2(new_n716_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n727_), .B(new_n728_), .C1(new_n733_), .C2(new_n724_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n728_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n498_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n724_), .B1(new_n717_), .B2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n737_), .B2(new_n726_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n734_), .A2(new_n738_), .ZN(G1329gat));
  NOR2_X1   g538(.A1(new_n484_), .A2(new_n487_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(new_n465_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n717_), .A2(new_n720_), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(G43gat), .B1(new_n698_), .B2(new_n490_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n742_), .A2(new_n744_), .A3(new_n746_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1330gat));
  AOI21_X1  g549(.A(G50gat), .B1(new_n698_), .B2(new_n450_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n450_), .A2(G50gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n721_), .B2(new_n752_), .ZN(G1331gat));
  NOR4_X1   g552(.A1(new_n501_), .A2(new_n695_), .A3(new_n569_), .A4(new_n648_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G57gat), .B1(new_n754_), .B2(new_n459_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n570_), .A2(new_n601_), .ZN(new_n756_));
  NOR4_X1   g555(.A1(new_n756_), .A2(new_n501_), .A3(new_n618_), .A4(new_n655_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n460_), .A2(KEYINPUT110), .ZN(new_n758_));
  MUX2_X1   g557(.A(KEYINPUT110), .B(new_n758_), .S(G57gat), .Z(new_n759_));
  AOI21_X1  g558(.A(new_n755_), .B1(new_n757_), .B2(new_n759_), .ZN(G1332gat));
  INV_X1    g559(.A(G64gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n757_), .B2(new_n458_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT48), .Z(new_n763_));
  NAND3_X1  g562(.A1(new_n754_), .A2(new_n761_), .A3(new_n458_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT111), .ZN(G1333gat));
  INV_X1    g565(.A(G71gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n757_), .B2(new_n490_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT49), .Z(new_n769_));
  NAND3_X1  g568(.A1(new_n754_), .A2(new_n767_), .A3(new_n490_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1334gat));
  AOI21_X1  g570(.A(new_n429_), .B1(new_n757_), .B2(new_n450_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n494_), .A2(G78gat), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT113), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n754_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n774_), .A2(new_n777_), .ZN(G1335gat));
  AND4_X1   g577(.A1(new_n694_), .A2(new_n601_), .A3(new_n570_), .A4(new_n697_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G85gat), .B1(new_n779_), .B2(new_n459_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n756_), .A2(new_n619_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n714_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n714_), .A2(KEYINPUT114), .A3(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n459_), .A2(G85gat), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT115), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n780_), .B1(new_n786_), .B2(new_n788_), .ZN(G1336gat));
  INV_X1    g588(.A(G92gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n779_), .A2(new_n790_), .A3(new_n458_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n498_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n790_), .ZN(G1337gat));
  NOR2_X1   g592(.A1(new_n740_), .A2(new_n507_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n779_), .A2(new_n794_), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT116), .Z(new_n796_));
  AOI21_X1  g595(.A(new_n491_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n797_));
  INV_X1    g596(.A(G99gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g599(.A1(new_n779_), .A2(new_n439_), .A3(new_n450_), .ZN(new_n801_));
  OAI21_X1  g600(.A(G106gat), .B1(new_n782_), .B2(new_n494_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n802_), .A2(KEYINPUT52), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(KEYINPUT52), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n801_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT53), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n801_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1339gat));
  NAND4_X1  g608(.A1(new_n569_), .A2(new_n601_), .A3(new_n619_), .A4(new_n647_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n810_), .B(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n597_), .B1(new_n592_), .B2(new_n588_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n588_), .B2(new_n587_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n600_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n563_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n547_), .A2(new_n548_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n547_), .A2(new_n817_), .A3(new_n548_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n559_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(KEYINPUT56), .ZN(new_n824_));
  INV_X1    g623(.A(new_n562_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n601_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT56), .B1(new_n822_), .B2(new_n823_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n816_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n696_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n822_), .A2(KEYINPUT56), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT56), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n559_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n815_), .A2(new_n562_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n647_), .B1(new_n832_), .B2(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n833_), .A2(KEYINPUT58), .A3(new_n836_), .A4(new_n835_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n830_), .A2(new_n831_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n547_), .A2(new_n548_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT55), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n549_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n821_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT117), .B1(new_n846_), .B2(new_n559_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n824_), .B(new_n826_), .C1(new_n847_), .C2(KEYINPUT56), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n655_), .B1(new_n848_), .B2(new_n816_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n841_), .B1(new_n849_), .B2(KEYINPUT57), .ZN(new_n850_));
  AND4_X1   g649(.A1(new_n841_), .A2(new_n829_), .A3(KEYINPUT57), .A4(new_n696_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n840_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n812_), .B1(new_n852_), .B2(new_n618_), .ZN(new_n853_));
  OR4_X1    g652(.A1(new_n460_), .A2(new_n458_), .A3(new_n450_), .A4(new_n740_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT119), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT59), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n837_), .A2(new_n832_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n707_), .A3(new_n839_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n849_), .B2(KEYINPUT57), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT118), .B1(new_n830_), .B2(new_n831_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n849_), .A2(new_n841_), .A3(KEYINPUT57), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n857_), .B1(new_n863_), .B2(new_n619_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n852_), .A2(KEYINPUT121), .A3(new_n618_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n812_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n855_), .A2(KEYINPUT120), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n855_), .A2(KEYINPUT120), .ZN(new_n868_));
  OR3_X1    g667(.A1(new_n867_), .A2(new_n868_), .A3(KEYINPUT59), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n856_), .B1(new_n866_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT122), .B(new_n856_), .C1(new_n866_), .C2(new_n869_), .ZN(new_n873_));
  INV_X1    g672(.A(G113gat), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n601_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n872_), .A2(new_n873_), .A3(new_n875_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n853_), .A2(new_n855_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n874_), .B1(new_n877_), .B2(new_n601_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1340gat));
  OAI21_X1  g678(.A(G120gat), .B1(new_n870_), .B2(new_n569_), .ZN(new_n880_));
  INV_X1    g679(.A(G120gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n569_), .B2(KEYINPUT60), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(KEYINPUT60), .B2(new_n881_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n880_), .B1(new_n877_), .B2(new_n883_), .ZN(G1341gat));
  INV_X1    g683(.A(G127gat), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n618_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n872_), .A2(new_n873_), .A3(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n885_), .B1(new_n877_), .B2(new_n618_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1342gat));
  INV_X1    g688(.A(G134gat), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n647_), .A2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n872_), .A2(new_n873_), .A3(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n877_), .B2(new_n696_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1343gat));
  INV_X1    g693(.A(new_n853_), .ZN(new_n895_));
  NOR4_X1   g694(.A1(new_n490_), .A2(new_n458_), .A3(new_n460_), .A4(new_n494_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n601_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n348_), .ZN(G1344gat));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n569_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n349_), .ZN(G1345gat));
  NAND3_X1  g700(.A1(new_n895_), .A2(new_n619_), .A3(new_n896_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT61), .B(G155gat), .Z(new_n903_));
  OR2_X1    g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT123), .B(KEYINPUT124), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n903_), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n904_), .A2(new_n905_), .A3(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n904_), .B2(new_n906_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1346gat));
  OAI21_X1  g708(.A(G162gat), .B1(new_n897_), .B2(new_n647_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n696_), .A2(G162gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n897_), .B2(new_n911_), .ZN(G1347gat));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n864_), .A2(new_n865_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n812_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n490_), .A2(new_n460_), .A3(new_n458_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT125), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n450_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n913_), .B1(new_n916_), .B2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n919_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n866_), .A2(KEYINPUT126), .A3(new_n921_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n260_), .B(new_n695_), .C1(new_n920_), .C2(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n916_), .A2(new_n695_), .A3(new_n919_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n924_), .A2(new_n925_), .A3(G169gat), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n924_), .B2(G169gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n923_), .B1(new_n926_), .B2(new_n927_), .ZN(G1348gat));
  NOR2_X1   g727(.A1(new_n853_), .A2(new_n450_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n918_), .A2(new_n261_), .A3(new_n569_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n916_), .A2(new_n913_), .A3(new_n919_), .ZN(new_n932_));
  OAI21_X1  g731(.A(KEYINPUT126), .B1(new_n866_), .B2(new_n921_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n570_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n931_), .B1(new_n935_), .B2(new_n261_), .ZN(G1349gat));
  NOR2_X1   g735(.A1(new_n918_), .A2(new_n618_), .ZN(new_n937_));
  AOI21_X1  g736(.A(G183gat), .B1(new_n929_), .B2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n618_), .A2(new_n238_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n934_), .B2(new_n939_), .ZN(G1350gat));
  OAI211_X1 g739(.A(new_n233_), .B(new_n655_), .C1(new_n920_), .C2(new_n922_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n647_), .B1(new_n932_), .B2(new_n933_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n229_), .B2(new_n942_), .ZN(G1351gat));
  NOR3_X1   g742(.A1(new_n490_), .A2(new_n461_), .A3(new_n498_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n895_), .A2(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n601_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(new_n207_), .ZN(G1352gat));
  NOR2_X1   g746(.A1(new_n945_), .A2(new_n569_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(new_n209_), .ZN(G1353gat));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n950_));
  NOR2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n951_), .B1(new_n945_), .B2(new_n618_), .ZN(new_n952_));
  XOR2_X1   g751(.A(KEYINPUT63), .B(G211gat), .Z(new_n953_));
  NAND4_X1  g752(.A1(new_n895_), .A2(new_n619_), .A3(new_n944_), .A4(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n950_), .B1(new_n952_), .B2(new_n954_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n955_), .B1(new_n950_), .B2(new_n954_), .ZN(G1354gat));
  OAI21_X1  g755(.A(G218gat), .B1(new_n945_), .B2(new_n647_), .ZN(new_n957_));
  OR2_X1    g756(.A1(new_n696_), .A2(G218gat), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n945_), .B2(new_n958_), .ZN(G1355gat));
endmodule


