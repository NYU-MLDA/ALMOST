//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_;
  INV_X1    g000(.A(G204gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G197gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT88), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n202_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT21), .ZN(new_n207_));
  INV_X1    g006(.A(G197gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G204gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n207_), .B1(new_n203_), .B2(new_n209_), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n212_), .A2(KEYINPUT87), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(KEYINPUT87), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n210_), .B(new_n211_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT89), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n211_), .A2(new_n207_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n205_), .A2(new_n209_), .A3(new_n206_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n216_), .B1(new_n215_), .B2(new_n219_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G228gat), .A2(G233gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT85), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G141gat), .ZN(new_n233_));
  INV_X1    g032(.A(G148gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G141gat), .A2(G148gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT86), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT2), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n242_), .B(new_n243_), .C1(new_n235_), .C2(KEYINPUT3), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n228_), .B(new_n229_), .C1(new_n240_), .C2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n237_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n225_), .B1(new_n246_), .B2(KEYINPUT29), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n223_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n215_), .A2(new_n219_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT91), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT91), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n215_), .A2(new_n251_), .A3(new_n219_), .ZN(new_n252_));
  XOR2_X1   g051(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n253_));
  AOI22_X1  g052(.A1(new_n250_), .A2(new_n252_), .B1(new_n246_), .B2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n248_), .B1(new_n254_), .B2(new_n224_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G78gat), .B(G106gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT92), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n248_), .B(new_n257_), .C1(new_n224_), .C2(new_n254_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT93), .A3(new_n260_), .ZN(new_n261_));
  OR3_X1    g060(.A1(new_n255_), .A2(KEYINPUT93), .A3(new_n258_), .ZN(new_n262_));
  OR3_X1    g061(.A1(new_n246_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT28), .B1(new_n246_), .B2(KEYINPUT29), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G22gat), .B(G50gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n263_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n261_), .A2(new_n262_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n254_), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n272_), .A2(new_n225_), .B1(new_n223_), .B2(new_n247_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n256_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT94), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT95), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n270_), .B1(new_n260_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT94), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n255_), .A2(new_n278_), .A3(new_n256_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n273_), .A2(KEYINPUT95), .A3(new_n257_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n275_), .A2(new_n277_), .A3(new_n279_), .A4(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n271_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT81), .B(G190gat), .ZN(new_n284_));
  INV_X1    g083(.A(G183gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT23), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(G169gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT25), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(G183gat), .ZN(new_n294_));
  INV_X1    g093(.A(G190gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n285_), .A2(KEYINPUT25), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT80), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT80), .B1(new_n285_), .B2(KEYINPUT25), .ZN(new_n299_));
  OAI221_X1 g098(.A(new_n294_), .B1(KEYINPUT26), .B2(new_n295_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n284_), .A2(KEYINPUT26), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n301_), .A2(KEYINPUT82), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(KEYINPUT82), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n300_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n287_), .A2(KEYINPUT23), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT23), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(G183gat), .A3(G190gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT24), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n305_), .A2(new_n307_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n310_), .A2(KEYINPUT83), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(KEYINPUT83), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n308_), .B1(G169gat), .B2(G176gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n313_), .B1(G169gat), .B2(G176gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n292_), .B1(new_n304_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n223_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT20), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G226gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT19), .ZN(new_n320_));
  INV_X1    g119(.A(new_n249_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n288_), .B1(G183gat), .B2(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n291_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n296_), .A2(new_n294_), .ZN(new_n324_));
  XOR2_X1   g123(.A(KEYINPUT26), .B(G190gat), .Z(new_n325_));
  OAI211_X1 g124(.A(new_n314_), .B(new_n310_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  AOI211_X1 g126(.A(new_n318_), .B(new_n320_), .C1(new_n321_), .C2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n317_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n249_), .A2(KEYINPUT89), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n316_), .B1(new_n330_), .B2(new_n220_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT96), .B1(new_n331_), .B2(new_n318_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT96), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n333_), .B(KEYINPUT20), .C1(new_n223_), .C2(new_n316_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n321_), .A2(new_n327_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n332_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n329_), .B1(new_n336_), .B2(new_n320_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT18), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  NOR2_X1   g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n341_), .ZN(new_n343_));
  AOI211_X1 g142(.A(new_n343_), .B(new_n329_), .C1(new_n336_), .C2(new_n320_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT33), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G127gat), .B(G134gat), .Z(new_n348_));
  XOR2_X1   g147(.A(G113gat), .B(G120gat), .Z(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G127gat), .B(G134gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G113gat), .B(G120gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT84), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n350_), .A2(KEYINPUT84), .A3(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n246_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n237_), .A2(new_n245_), .A3(new_n354_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n347_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT4), .B1(new_n358_), .B2(new_n246_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n360_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n363_), .B2(KEYINPUT4), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n361_), .B1(new_n364_), .B2(new_n347_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G1gat), .B(G29gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(G85gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT0), .B(G57gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n345_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n369_), .ZN(new_n371_));
  AOI211_X1 g170(.A(new_n346_), .B(new_n362_), .C1(new_n363_), .C2(KEYINPUT4), .ZN(new_n372_));
  OAI211_X1 g171(.A(KEYINPUT33), .B(new_n371_), .C1(new_n372_), .C2(new_n361_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n359_), .A2(new_n360_), .A3(new_n347_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n374_), .A2(new_n369_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(new_n364_), .B2(new_n347_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT97), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n375_), .B(KEYINPUT97), .C1(new_n364_), .C2(new_n347_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n370_), .A2(new_n373_), .A3(new_n378_), .A4(new_n379_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n342_), .A2(new_n344_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n341_), .A2(KEYINPUT32), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI211_X1 g182(.A(new_n383_), .B(new_n329_), .C1(new_n336_), .C2(new_n320_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n250_), .A2(new_n252_), .A3(new_n327_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT99), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n317_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n320_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n320_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n332_), .A2(new_n334_), .A3(new_n392_), .A4(new_n335_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n382_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n365_), .B(new_n371_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n384_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n283_), .B1(new_n381_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT100), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n391_), .A2(new_n393_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n343_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n337_), .A2(new_n341_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT27), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT101), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT27), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT101), .A4(KEYINPUT27), .ZN(new_n407_));
  INV_X1    g206(.A(new_n395_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n408_), .B1(new_n271_), .B2(new_n281_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n404_), .A2(new_n406_), .A3(new_n407_), .A4(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT100), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n411_), .B(new_n283_), .C1(new_n381_), .C2(new_n396_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n398_), .A2(new_n410_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414_));
  INV_X1    g213(.A(G15gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT30), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n316_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n358_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G71gat), .B(G99gat), .ZN(new_n421_));
  INV_X1    g220(.A(G43gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT31), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n420_), .B(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n413_), .A2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n406_), .A2(new_n407_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n425_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n395_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  AND4_X1   g229(.A1(new_n283_), .A2(new_n427_), .A3(new_n430_), .A4(new_n404_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n426_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G229gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G36gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G29gat), .ZN(new_n437_));
  INV_X1    g236(.A(G29gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(G36gat), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n437_), .A2(new_n439_), .A3(KEYINPUT70), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT70), .B1(new_n437_), .B2(new_n439_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT71), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n439_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT70), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT71), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n437_), .A2(new_n439_), .A3(KEYINPUT70), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G43gat), .B(G50gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n442_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n449_), .B1(new_n442_), .B2(new_n448_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G1gat), .B(G8gat), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n454_), .A2(KEYINPUT76), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(KEYINPUT76), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G15gat), .B(G22gat), .ZN(new_n458_));
  INV_X1    g257(.A(G1gat), .ZN(new_n459_));
  INV_X1    g258(.A(G8gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT14), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n457_), .A2(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n455_), .A2(new_n461_), .A3(new_n458_), .A4(new_n456_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n453_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n442_), .A2(new_n448_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n449_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n450_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n471_), .A2(new_n465_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n435_), .B1(new_n467_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT15), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n470_), .A2(KEYINPUT15), .A3(new_n450_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n466_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n453_), .A2(new_n466_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n434_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n473_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G113gat), .B(G141gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G169gat), .B(G197gat), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n481_), .B(new_n482_), .Z(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n473_), .B(new_n483_), .C1(new_n477_), .C2(new_n479_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n433_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G57gat), .B(G64gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT11), .ZN(new_n490_));
  XOR2_X1   g289(.A(G71gat), .B(G78gat), .Z(new_n491_));
  OR2_X1    g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n489_), .A2(KEYINPUT11), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n491_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G231gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(new_n466_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT78), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G127gat), .B(G155gat), .Z(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G183gat), .B(G211gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT17), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n500_), .B(new_n506_), .ZN(new_n507_));
  OR3_X1    g306(.A1(new_n498_), .A2(KEYINPUT17), .A3(new_n505_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n509_), .B(KEYINPUT79), .Z(new_n510_));
  XNOR2_X1  g309(.A(G190gat), .B(G218gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G134gat), .B(G162gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT36), .Z(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT67), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G99gat), .A2(G106gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT6), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT6), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(G99gat), .A3(G106gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT7), .ZN(new_n525_));
  INV_X1    g324(.A(G99gat), .ZN(new_n526_));
  INV_X1    g325(.A(G106gat), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT67), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(new_n516_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n519_), .A2(new_n524_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G85gat), .ZN(new_n532_));
  INV_X1    g331(.A(G92gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n515_), .B1(new_n531_), .B2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n536_), .A2(KEYINPUT8), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n521_), .A2(new_n523_), .A3(KEYINPUT66), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT66), .B1(new_n521_), .B2(new_n523_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n528_), .A2(new_n516_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n540_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT68), .B1(new_n538_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT66), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n524_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n521_), .A2(new_n523_), .A3(KEYINPUT66), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n545_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n539_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT68), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n544_), .A2(KEYINPUT67), .B1(new_n521_), .B2(new_n523_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n536_), .B1(new_n554_), .B2(new_n530_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n552_), .B(new_n553_), .C1(new_n555_), .C2(new_n515_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n547_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n549_), .A2(new_n550_), .ZN(new_n558_));
  OR2_X1    g357(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n527_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n534_), .A2(KEYINPUT9), .A3(new_n535_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT65), .B(G92gat), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n532_), .A2(KEYINPUT9), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n561_), .B(new_n562_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n558_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n557_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n475_), .A2(new_n476_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT35), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n531_), .A2(new_n537_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT8), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n566_), .B1(new_n577_), .B2(new_n552_), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n578_), .A2(new_n453_), .B1(new_n574_), .B2(new_n573_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n570_), .A2(KEYINPUT72), .A3(new_n575_), .A4(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(KEYINPUT72), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n575_), .A2(KEYINPUT72), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n557_), .A2(new_n567_), .B1(new_n476_), .B2(new_n475_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n573_), .A2(new_n574_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n552_), .B1(new_n555_), .B2(new_n515_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n567_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n584_), .B1(new_n586_), .B2(new_n471_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n581_), .B(new_n582_), .C1(new_n583_), .C2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT73), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n580_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n580_), .B2(new_n588_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n514_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT74), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT37), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n580_), .A2(new_n588_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n513_), .A2(KEYINPUT36), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  OAI211_X1 g397(.A(KEYINPUT74), .B(new_n514_), .C1(new_n590_), .C2(new_n591_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n594_), .A2(new_n595_), .A3(new_n598_), .A4(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT75), .ZN(new_n601_));
  INV_X1    g400(.A(new_n514_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n598_), .B1(new_n602_), .B2(new_n596_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n603_), .B2(KEYINPUT37), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G120gat), .B(G148gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT5), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G176gat), .B(G204gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n607_), .B(new_n608_), .Z(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n585_), .A2(new_n495_), .A3(new_n567_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT12), .ZN(new_n613_));
  INV_X1    g412(.A(new_n495_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n586_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n612_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(KEYINPUT12), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n568_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT64), .Z(new_n621_));
  NAND3_X1  g420(.A1(new_n616_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n615_), .B2(new_n611_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n610_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n622_), .A2(new_n624_), .A3(new_n610_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT13), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n599_), .A2(new_n598_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n630_), .A2(new_n601_), .A3(new_n595_), .A4(new_n594_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n510_), .A2(new_n605_), .A3(new_n629_), .A4(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n488_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n459_), .A3(new_n408_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT38), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n431_), .B1(new_n413_), .B2(new_n425_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n599_), .A2(new_n598_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n596_), .A2(KEYINPUT73), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n580_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT74), .B1(new_n641_), .B2(new_n514_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT102), .B1(new_n638_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n594_), .A2(new_n644_), .A3(new_n598_), .A4(new_n599_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n637_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n629_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n487_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n509_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n647_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G1gat), .B1(new_n653_), .B2(new_n395_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n634_), .A2(new_n635_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n636_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT103), .ZN(G1324gat));
  NAND2_X1  g456(.A1(new_n427_), .A2(new_n404_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n633_), .A2(new_n460_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n652_), .A2(new_n658_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(G8gat), .ZN(new_n662_));
  AOI211_X1 g461(.A(KEYINPUT39), .B(new_n460_), .C1(new_n652_), .C2(new_n658_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g464(.A(new_n415_), .B1(new_n652_), .B2(new_n428_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT105), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n633_), .A2(new_n415_), .A3(new_n428_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n666_), .A2(new_n668_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(G1326gat));
  INV_X1    g471(.A(G22gat), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n282_), .B(KEYINPUT106), .Z(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n652_), .B2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT42), .Z(new_n677_));
  NAND3_X1  g476(.A1(new_n633_), .A2(new_n673_), .A3(new_n675_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1327gat));
  AOI21_X1  g478(.A(new_n649_), .B1(new_n426_), .B2(new_n432_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n510_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n629_), .A3(new_n646_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT107), .B1(new_n680_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n685_));
  NOR4_X1   g484(.A1(new_n637_), .A2(new_n682_), .A3(new_n685_), .A4(new_n649_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n438_), .B1(new_n688_), .B2(new_n395_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n605_), .A2(new_n631_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n433_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n510_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n648_), .A2(new_n649_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n433_), .A2(KEYINPUT43), .A3(new_n690_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n693_), .A2(KEYINPUT44), .A3(new_n694_), .A4(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n690_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n692_), .B1(new_n637_), .B2(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n695_), .A2(new_n698_), .A3(new_n681_), .A4(new_n694_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n696_), .A2(new_n701_), .A3(G29gat), .A4(new_n408_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n689_), .A2(new_n702_), .ZN(G1328gat));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n685_), .B1(new_n488_), .B2(new_n682_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n680_), .A2(KEYINPUT107), .A3(new_n683_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n658_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n708_), .A2(G36gat), .ZN(new_n709_));
  AND4_X1   g508(.A1(new_n705_), .A2(new_n706_), .A3(new_n707_), .A4(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n705_), .B1(new_n687_), .B2(new_n709_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n704_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n696_), .A2(new_n701_), .A3(new_n658_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G36gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n706_), .A2(new_n707_), .A3(new_n709_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT108), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n687_), .A2(new_n705_), .A3(new_n709_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(KEYINPUT45), .A3(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n712_), .A2(new_n714_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n712_), .A2(new_n714_), .A3(KEYINPUT46), .A4(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  OAI21_X1  g522(.A(new_n422_), .B1(new_n688_), .B2(new_n425_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n696_), .A2(new_n701_), .A3(G43gat), .A4(new_n428_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT47), .ZN(G1330gat));
  AND4_X1   g526(.A1(G50gat), .A2(new_n696_), .A3(new_n282_), .A4(new_n701_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G50gat), .B1(new_n687_), .B2(new_n675_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1331gat));
  AND3_X1   g529(.A1(new_n510_), .A2(new_n605_), .A3(new_n631_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n433_), .A2(new_n649_), .A3(new_n648_), .A4(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT109), .ZN(new_n733_));
  AOI21_X1  g532(.A(G57gat), .B1(new_n733_), .B2(new_n408_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n629_), .A2(new_n487_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n647_), .A2(new_n510_), .A3(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n395_), .A2(KEYINPUT110), .ZN(new_n737_));
  MUX2_X1   g536(.A(KEYINPUT110), .B(new_n737_), .S(G57gat), .Z(new_n738_));
  AOI21_X1  g537(.A(new_n734_), .B1(new_n736_), .B2(new_n738_), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n736_), .B2(new_n658_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT48), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n733_), .A2(new_n740_), .A3(new_n658_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n736_), .B2(new_n428_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT49), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n733_), .A2(new_n745_), .A3(new_n428_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n736_), .A2(new_n675_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G78gat), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT111), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n751_), .B(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT50), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n674_), .A2(G78gat), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT112), .Z(new_n759_));
  NAND2_X1  g558(.A1(new_n733_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n754_), .A2(new_n757_), .A3(new_n760_), .ZN(G1335gat));
  AND3_X1   g560(.A1(new_n646_), .A2(new_n648_), .A3(new_n681_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n433_), .A2(new_n649_), .A3(new_n762_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n763_), .A2(KEYINPUT113), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(KEYINPUT113), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(new_n532_), .A3(new_n408_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n695_), .A2(new_n698_), .A3(new_n681_), .A4(new_n735_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768_), .B2(new_n395_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1336gat));
  NOR3_X1   g569(.A1(new_n768_), .A2(new_n708_), .A3(new_n563_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n766_), .A2(new_n658_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(new_n533_), .ZN(G1337gat));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n559_), .A2(new_n560_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n428_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n774_), .B1(new_n766_), .B2(new_n777_), .ZN(new_n778_));
  AOI211_X1 g577(.A(KEYINPUT114), .B(new_n776_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G99gat), .B1(new_n768_), .B2(new_n425_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT115), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT51), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n782_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n784_), .B(new_n785_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n783_), .A2(new_n786_), .ZN(G1338gat));
  NAND3_X1  g586(.A1(new_n766_), .A2(new_n527_), .A3(new_n282_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n768_), .A2(new_n283_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(G106gat), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n789_), .B(G106gat), .C1(new_n768_), .C2(new_n283_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n788_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT53), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n796_), .B(new_n788_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1339gat));
  INV_X1    g597(.A(new_n627_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n649_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n613_), .B1(new_n578_), .B2(new_n495_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n566_), .B1(new_n547_), .B2(new_n556_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n802_), .B(new_n611_), .C1(new_n803_), .C2(new_n617_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n621_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n801_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n805_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n616_), .A2(new_n619_), .A3(KEYINPUT55), .A4(new_n621_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n809_), .A2(KEYINPUT56), .A3(new_n609_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT56), .B1(new_n809_), .B2(new_n609_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n800_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n434_), .B1(new_n467_), .B2(new_n472_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n478_), .A2(new_n435_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n814_), .B(new_n484_), .C1(new_n477_), .C2(new_n815_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n486_), .A2(new_n816_), .A3(KEYINPUT116), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT116), .B1(new_n486_), .B2(new_n816_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n628_), .B(new_n813_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n819_));
  OAI22_X1  g618(.A1(new_n799_), .A2(new_n625_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT117), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n812_), .A2(new_n819_), .A3(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n822_), .A2(new_n643_), .A3(KEYINPUT57), .A4(new_n645_), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n823_), .A2(KEYINPUT118), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(KEYINPUT118), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n486_), .A2(new_n816_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n486_), .A2(new_n816_), .A3(KEYINPUT116), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n799_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT58), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n822_), .A2(new_n643_), .A3(new_n645_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n833_), .A2(new_n690_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n509_), .B1(new_n826_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n731_), .A2(new_n838_), .A3(new_n649_), .A4(new_n629_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT54), .B1(new_n632_), .B2(new_n487_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n837_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n658_), .A2(new_n282_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(new_n408_), .A3(new_n428_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(G113gat), .B1(new_n845_), .B2(new_n487_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n842_), .A2(new_n844_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n690_), .A2(new_n833_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n834_), .A2(new_n835_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT119), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n836_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n851_), .A2(new_n853_), .A3(new_n826_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n841_), .B1(new_n854_), .B2(new_n681_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n844_), .A2(KEYINPUT59), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n847_), .A2(KEYINPUT59), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(G113gat), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n487_), .A2(KEYINPUT120), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(G113gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n846_), .B1(new_n858_), .B2(new_n862_), .ZN(G1340gat));
  INV_X1    g662(.A(KEYINPUT60), .ZN(new_n864_));
  AOI21_X1  g663(.A(G120gat), .B1(new_n648_), .B2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n864_), .B2(G120gat), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n845_), .A2(new_n866_), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(KEYINPUT121), .Z(new_n868_));
  NAND2_X1  g667(.A1(new_n858_), .A2(new_n648_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(G120gat), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1341gat));
  NAND2_X1  g670(.A1(new_n858_), .A2(new_n509_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G127gat), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n681_), .A2(G127gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n847_), .B2(new_n874_), .ZN(G1342gat));
  AOI21_X1  g674(.A(G134gat), .B1(new_n845_), .B2(new_n646_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT122), .B(G134gat), .Z(new_n877_));
  NOR2_X1   g676(.A1(new_n697_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n858_), .B2(new_n878_), .ZN(G1343gat));
  NOR2_X1   g678(.A1(new_n842_), .A2(new_n428_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n658_), .A2(new_n283_), .A3(new_n395_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n649_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n233_), .ZN(G1344gat));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n629_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n234_), .ZN(G1345gat));
  INV_X1    g685(.A(new_n882_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n510_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT61), .B(G155gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1346gat));
  OAI21_X1  g689(.A(G162gat), .B1(new_n882_), .B2(new_n697_), .ZN(new_n891_));
  INV_X1    g690(.A(G162gat), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n646_), .A2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n891_), .B1(new_n882_), .B2(new_n893_), .ZN(G1347gat));
  NOR2_X1   g693(.A1(new_n708_), .A2(new_n429_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n674_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n487_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n823_), .A2(KEYINPUT118), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n823_), .A2(KEYINPUT118), .ZN(new_n900_));
  OAI22_X1  g699(.A1(new_n836_), .A2(new_n852_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n850_), .A2(KEYINPUT119), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n681_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n841_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n898_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(G169gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT123), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n908_), .B(G169gat), .C1(new_n855_), .C2(new_n898_), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n907_), .A2(KEYINPUT62), .A3(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n911_), .B1(new_n855_), .B2(new_n896_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n850_), .A2(KEYINPUT119), .B1(new_n824_), .B2(new_n825_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n510_), .B1(new_n913_), .B2(new_n853_), .ZN(new_n914_));
  OAI211_X1 g713(.A(KEYINPUT124), .B(new_n897_), .C1(new_n914_), .C2(new_n841_), .ZN(new_n915_));
  XOR2_X1   g714(.A(KEYINPUT22), .B(G169gat), .Z(new_n916_));
  NOR2_X1   g715(.A1(new_n649_), .A2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n912_), .A2(new_n915_), .A3(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919_));
  OAI211_X1 g718(.A(KEYINPUT123), .B(new_n919_), .C1(new_n905_), .C2(new_n906_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(KEYINPUT125), .B1(new_n910_), .B2(new_n921_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n907_), .A2(KEYINPUT62), .A3(new_n909_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n923_), .A2(new_n924_), .A3(new_n920_), .A4(new_n918_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n922_), .A2(new_n925_), .ZN(G1348gat));
  NAND3_X1  g725(.A1(new_n895_), .A2(G176gat), .A3(new_n648_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n842_), .A2(new_n282_), .A3(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n912_), .A2(new_n915_), .A3(new_n648_), .ZN(new_n929_));
  INV_X1    g728(.A(G176gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n928_), .B1(new_n929_), .B2(new_n930_), .ZN(G1349gat));
  NAND2_X1  g730(.A1(new_n895_), .A2(new_n510_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n842_), .A2(new_n282_), .A3(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(G183gat), .B1(new_n933_), .B2(KEYINPUT126), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n934_), .B1(KEYINPUT126), .B2(new_n933_), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n912_), .A2(new_n915_), .A3(new_n324_), .A4(new_n509_), .ZN(new_n936_));
  AND2_X1   g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1350gat));
  NAND2_X1  g736(.A1(new_n912_), .A2(new_n915_), .ZN(new_n938_));
  OAI21_X1  g737(.A(G190gat), .B1(new_n938_), .B2(new_n697_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n325_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n646_), .A2(new_n940_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n939_), .B1(new_n938_), .B2(new_n941_), .ZN(G1351gat));
  AND2_X1   g741(.A1(new_n658_), .A2(new_n409_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n880_), .A2(new_n943_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n649_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(new_n208_), .ZN(G1352gat));
  INV_X1    g745(.A(new_n944_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n648_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n202_), .A2(KEYINPUT127), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n948_), .B(new_n949_), .ZN(G1353gat));
  AOI21_X1  g749(.A(new_n650_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n947_), .A2(new_n951_), .ZN(new_n952_));
  OR2_X1    g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n952_), .B(new_n953_), .ZN(G1354gat));
  OAI21_X1  g753(.A(G218gat), .B1(new_n944_), .B2(new_n697_), .ZN(new_n955_));
  INV_X1    g754(.A(G218gat), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n646_), .A2(new_n956_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n955_), .B1(new_n944_), .B2(new_n957_), .ZN(G1355gat));
endmodule


