//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT30), .Z(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT77), .B(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206_));
  OR3_X1    g005(.A1(new_n205_), .A2(KEYINPUT78), .A3(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(G169gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT79), .B(G176gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT78), .B1(new_n205_), .B2(new_n206_), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n212_), .B(KEYINPUT23), .Z(new_n213_));
  NOR2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT76), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n211_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  NOR3_X1   g018(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n213_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT25), .B(G183gat), .Z(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n218_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n221_), .B(new_n225_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G71gat), .B(G99gat), .Z(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n219_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G15gat), .B(G43gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n230_), .B1(new_n219_), .B2(new_n228_), .ZN(new_n235_));
  NOR3_X1   g034(.A1(new_n232_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n219_), .A2(new_n228_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n229_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n233_), .B1(new_n238_), .B2(new_n231_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n204_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n234_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n238_), .A2(new_n233_), .A3(new_n231_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(new_n203_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n240_), .A2(KEYINPUT82), .A3(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G113gat), .B(G120gat), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT80), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n246_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n245_), .A2(new_n246_), .A3(KEYINPUT80), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT81), .Z(new_n253_));
  NAND2_X1  g052(.A1(new_n244_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n253_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n240_), .A2(KEYINPUT82), .A3(new_n255_), .A4(new_n243_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n254_), .A2(new_n258_), .A3(new_n256_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT2), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(KEYINPUT85), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT85), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n265_), .B1(new_n266_), .B2(KEYINPUT2), .ZN(new_n267_));
  OR2_X1    g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n268_), .A2(KEYINPUT3), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(KEYINPUT3), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n263_), .A2(KEYINPUT85), .A3(new_n264_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n267_), .A2(new_n269_), .A3(new_n270_), .A4(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT1), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT84), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n274_), .A2(KEYINPUT1), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n274_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n273_), .A4(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(new_n263_), .A3(new_n268_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n275_), .A2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n284_));
  OR3_X1    g083(.A1(new_n283_), .A2(KEYINPUT29), .A3(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n284_), .B1(new_n283_), .B2(KEYINPUT29), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G22gat), .B(G50gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G211gat), .B(G218gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(G197gat), .B(G204gat), .Z(new_n291_));
  OAI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(KEYINPUT21), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(KEYINPUT21), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(new_n283_), .B2(KEYINPUT29), .ZN(new_n295_));
  AND2_X1   g094(.A1(G228gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G78gat), .B(G106gat), .Z(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n289_), .B1(KEYINPUT87), .B2(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n297_), .A2(new_n298_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n299_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n301_), .A2(new_n289_), .A3(KEYINPUT87), .A4(new_n299_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G1gat), .B(G29gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(G57gat), .B(G85gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  AND2_X1   g110(.A1(new_n247_), .A2(new_n249_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n283_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G225gat), .A2(G233gat), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n275_), .A2(new_n282_), .B1(new_n251_), .B2(new_n250_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n315_), .A2(KEYINPUT4), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n313_), .A2(new_n316_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n318_), .B1(new_n319_), .B2(KEYINPUT4), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n317_), .B(KEYINPUT92), .C1(new_n320_), .C2(new_n314_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n317_), .A2(KEYINPUT92), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n311_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n311_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n319_), .A2(new_n314_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n283_), .A2(new_n312_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT4), .B1(new_n327_), .B2(new_n315_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n318_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AOI211_X1 g129(.A(new_n325_), .B(new_n326_), .C1(new_n314_), .C2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT33), .B1(new_n324_), .B2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n314_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n317_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT92), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n325_), .B1(new_n336_), .B2(new_n322_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT33), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n340_), .B(KEYINPUT88), .Z(new_n341_));
  XOR2_X1   g140(.A(new_n341_), .B(KEYINPUT19), .Z(new_n342_));
  INV_X1    g141(.A(new_n217_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n224_), .B(KEYINPUT89), .ZN(new_n344_));
  OAI221_X1 g143(.A(new_n221_), .B1(new_n226_), .B2(new_n343_), .C1(new_n344_), .C2(new_n222_), .ZN(new_n345_));
  INV_X1    g144(.A(G169gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT22), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n209_), .A2(new_n208_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n218_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT90), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n345_), .B1(new_n350_), .B2(new_n215_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n294_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT20), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n294_), .B1(new_n219_), .B2(new_n228_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n342_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n352_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n342_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n219_), .A2(new_n228_), .A3(new_n294_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n356_), .A2(KEYINPUT20), .A3(new_n357_), .A4(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT18), .B(G64gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G92gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G8gat), .B(G36gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n364_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n355_), .A2(new_n366_), .A3(new_n359_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n332_), .A2(new_n339_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n364_), .A2(KEYINPUT32), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n360_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n357_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n356_), .A2(KEYINPUT20), .A3(new_n358_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n373_), .B1(new_n374_), .B2(new_n357_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n371_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n321_), .A2(new_n311_), .A3(new_n323_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n372_), .B(new_n377_), .C1(new_n379_), .C2(new_n324_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n306_), .B1(new_n370_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n365_), .A2(KEYINPUT93), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT27), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n375_), .B2(new_n366_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT93), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n360_), .A2(new_n385_), .A3(new_n364_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n382_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n368_), .A2(new_n383_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n303_), .A2(new_n304_), .A3(new_n378_), .A4(new_n337_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n262_), .B1(new_n381_), .B2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n379_), .A2(new_n324_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n260_), .A2(new_n393_), .A3(new_n261_), .A4(new_n305_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n394_), .A2(new_n389_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G120gat), .B(G148gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(G176gat), .B(G204gat), .Z(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G85gat), .B(G92gat), .Z(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(KEYINPUT9), .B2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(KEYINPUT10), .B(G99gat), .Z(new_n410_));
  INV_X1    g209(.A(G106gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT9), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(G85gat), .A3(G92gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n409_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT8), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT7), .ZN(new_n417_));
  INV_X1    g216(.A(G99gat), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(new_n411_), .A4(KEYINPUT64), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT64), .ZN(new_n420_));
  OAI22_X1  g219(.A1(new_n420_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(KEYINPUT7), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n416_), .B(new_n408_), .C1(new_n423_), .C2(new_n407_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AND3_X1   g224(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(new_n404_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n427_), .A2(new_n422_), .A3(new_n421_), .A4(new_n419_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n416_), .B1(new_n428_), .B2(new_n408_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n415_), .B1(new_n425_), .B2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G57gat), .B(G64gat), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n431_), .A2(KEYINPUT11), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(KEYINPUT11), .ZN(new_n433_));
  XOR2_X1   g232(.A(G71gat), .B(G78gat), .Z(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n433_), .A2(new_n434_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n430_), .A2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n437_), .B(new_n415_), .C1(new_n425_), .C2(new_n429_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(KEYINPUT12), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT12), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n430_), .A2(new_n442_), .A3(new_n438_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G230gat), .A2(G233gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT65), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n445_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n449_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT65), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n439_), .A2(new_n440_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n449_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n403_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT65), .B1(new_n444_), .B2(new_n445_), .ZN(new_n456_));
  AOI211_X1 g255(.A(new_n447_), .B(new_n449_), .C1(new_n441_), .C2(new_n443_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n454_), .B(new_n403_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT13), .ZN(new_n460_));
  OR3_X1    g259(.A1(new_n455_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n460_), .B1(new_n455_), .B2(new_n459_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G15gat), .B(G22gat), .ZN(new_n464_));
  INV_X1    g263(.A(G1gat), .ZN(new_n465_));
  INV_X1    g264(.A(G8gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT14), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G1gat), .B(G8gat), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n469_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(G29gat), .A2(G36gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G29gat), .A2(G36gat), .ZN(new_n474_));
  OAI21_X1  g273(.A(G43gat), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G29gat), .ZN(new_n476_));
  INV_X1    g275(.A(G36gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G43gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G29gat), .A2(G36gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n475_), .A2(new_n481_), .A3(G50gat), .ZN(new_n482_));
  AOI21_X1  g281(.A(G50gat), .B1(new_n475_), .B2(new_n481_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT68), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G50gat), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n473_), .A2(new_n474_), .A3(G43gat), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n479_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n485_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT68), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n475_), .A2(new_n481_), .A3(G50gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n484_), .A2(KEYINPUT15), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT15), .B1(new_n484_), .B2(new_n491_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n472_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G229gat), .A2(G233gat), .ZN(new_n495_));
  AND4_X1   g294(.A1(new_n490_), .A2(new_n470_), .A3(new_n488_), .A4(new_n471_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n482_), .A2(new_n483_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n499_), .B1(new_n471_), .B2(new_n470_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(new_n496_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT75), .B1(new_n501_), .B2(new_n495_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT75), .ZN(new_n503_));
  INV_X1    g302(.A(new_n495_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n503_), .B(new_n504_), .C1(new_n500_), .C2(new_n496_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n498_), .A2(new_n502_), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(new_n346_), .ZN(new_n508_));
  INV_X1    g307(.A(G197gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n510_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n498_), .A2(new_n502_), .A3(new_n505_), .A4(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n463_), .A2(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n397_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT74), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G231gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n472_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(new_n438_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT70), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n520_), .B(new_n437_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT70), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT16), .B(G183gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G211gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G127gat), .B(G155gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT71), .B(KEYINPUT17), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n531_), .B(KEYINPUT72), .Z(new_n532_));
  NAND3_X1  g331(.A1(new_n523_), .A2(new_n525_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT73), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n529_), .B(KEYINPUT17), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n524_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n534_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n518_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(KEYINPUT74), .A3(new_n537_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G190gat), .B(G218gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(G134gat), .ZN(new_n545_));
  INV_X1    g344(.A(G162gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(KEYINPUT36), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT67), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT34), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(KEYINPUT35), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n484_), .A2(new_n491_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT15), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n484_), .A2(new_n491_), .A3(KEYINPUT15), .ZN(new_n558_));
  INV_X1    g357(.A(new_n429_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n424_), .ZN(new_n560_));
  AOI22_X1  g359(.A1(new_n557_), .A2(new_n558_), .B1(new_n415_), .B2(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(KEYINPUT35), .B(new_n553_), .C1(new_n561_), .C2(KEYINPUT69), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n430_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n560_), .A2(new_n499_), .A3(new_n415_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT69), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n563_), .A2(new_n568_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n565_), .A2(new_n569_), .A3(KEYINPUT35), .A4(new_n553_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n554_), .B1(new_n567_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n548_), .A2(KEYINPUT36), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n550_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n571_), .A2(new_n550_), .A3(new_n572_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n574_), .A2(KEYINPUT37), .A3(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT37), .B1(new_n574_), .B2(new_n575_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n543_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n517_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT94), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n393_), .B(KEYINPUT95), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n517_), .A2(KEYINPUT94), .A3(new_n578_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n581_), .A2(new_n465_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT38), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n574_), .A2(new_n575_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n538_), .A2(new_n539_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n517_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(G1gat), .B1(new_n590_), .B2(new_n393_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n585_), .A2(new_n586_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n587_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT96), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n587_), .A2(KEYINPUT96), .A3(new_n591_), .A4(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(G1324gat));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n599_));
  INV_X1    g398(.A(new_n389_), .ZN(new_n600_));
  OAI221_X1 g399(.A(G8gat), .B1(new_n598_), .B2(new_n599_), .C1(new_n590_), .C2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(KEYINPUT97), .A2(KEYINPUT39), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n581_), .A2(new_n584_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n466_), .A3(new_n389_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n603_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT40), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n603_), .A2(KEYINPUT40), .A3(new_n605_), .A4(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1325gat));
  OAI21_X1  g410(.A(G15gat), .B1(new_n590_), .B2(new_n262_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT41), .ZN(new_n615_));
  INV_X1    g414(.A(G15gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n262_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n604_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(G1326gat));
  OAI21_X1  g418(.A(G22gat), .B1(new_n590_), .B2(new_n305_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT42), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n305_), .A2(G22gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT99), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n604_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(G1327gat));
  NOR2_X1   g424(.A1(new_n576_), .A2(new_n577_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT43), .B1(new_n627_), .B2(KEYINPUT100), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT43), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n368_), .B1(new_n338_), .B2(new_n337_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n337_), .A2(new_n378_), .B1(new_n376_), .B2(new_n375_), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n332_), .A2(new_n631_), .B1(new_n632_), .B2(new_n372_), .ZN(new_n633_));
  OAI22_X1  g432(.A1(new_n633_), .A2(new_n306_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n395_), .B1(new_n634_), .B2(new_n262_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n629_), .B(new_n630_), .C1(new_n635_), .C2(new_n626_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n628_), .A2(new_n636_), .A3(new_n516_), .A4(new_n543_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT102), .B1(KEYINPUT101), .B2(KEYINPUT44), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n638_), .B1(KEYINPUT102), .B2(KEYINPUT44), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n638_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n637_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n582_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n543_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n588_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n517_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n517_), .A2(KEYINPUT103), .A3(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n393_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n476_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT104), .ZN(new_n654_));
  OAI22_X1  g453(.A1(new_n644_), .A2(new_n476_), .B1(new_n651_), .B2(new_n654_), .ZN(G1328gat));
  INV_X1    g454(.A(KEYINPUT46), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n641_), .A2(new_n643_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n477_), .B1(new_n657_), .B2(new_n389_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n649_), .A2(new_n477_), .A3(new_n389_), .A4(new_n650_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT45), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n656_), .B1(new_n658_), .B2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n659_), .B(KEYINPUT45), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n600_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n663_), .B(KEYINPUT46), .C1(new_n477_), .C2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(G1329gat));
  INV_X1    g465(.A(KEYINPUT47), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n637_), .A2(new_n642_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n617_), .B1(new_n668_), .B2(new_n640_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G43gat), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n262_), .A2(G43gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n649_), .A2(new_n650_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n667_), .B1(new_n670_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n672_), .ZN(new_n674_));
  AOI211_X1 g473(.A(KEYINPUT47), .B(new_n674_), .C1(new_n669_), .C2(G43gat), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1330gat));
  OAI211_X1 g475(.A(G50gat), .B(new_n306_), .C1(new_n668_), .C2(new_n640_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n485_), .B1(new_n651_), .B2(new_n305_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(G1331gat));
  INV_X1    g480(.A(new_n463_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(new_n514_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n635_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n578_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G57gat), .B1(new_n687_), .B2(new_n583_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n588_), .ZN(new_n689_));
  NOR4_X1   g488(.A1(new_n635_), .A2(new_n684_), .A3(new_n689_), .A4(new_n543_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(new_n652_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n688_), .B1(G57gat), .B2(new_n691_), .ZN(G1332gat));
  OR3_X1    g491(.A1(new_n686_), .A2(G64gat), .A3(new_n600_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n389_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G64gat), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(KEYINPUT48), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(KEYINPUT48), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT106), .ZN(G1333gat));
  INV_X1    g498(.A(G71gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n690_), .B2(new_n617_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT49), .Z(new_n702_));
  NAND3_X1  g501(.A1(new_n687_), .A2(new_n700_), .A3(new_n617_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1334gat));
  OR3_X1    g503(.A1(new_n686_), .A2(G78gat), .A3(new_n305_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n690_), .A2(new_n306_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G78gat), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(KEYINPUT50), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(KEYINPUT50), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(G1335gat));
  NAND2_X1  g511(.A1(new_n685_), .A2(new_n646_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G85gat), .B1(new_n714_), .B2(new_n583_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n628_), .A2(new_n636_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n684_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n628_), .A2(new_n636_), .A3(KEYINPUT108), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n543_), .A3(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(new_n393_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n715_), .B1(new_n721_), .B2(G85gat), .ZN(G1336gat));
  NAND2_X1  g521(.A1(new_n389_), .A2(G92gat), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT109), .Z(new_n724_));
  NOR2_X1   g523(.A1(new_n713_), .A2(new_n600_), .ZN(new_n725_));
  OAI22_X1  g524(.A1(new_n720_), .A2(new_n724_), .B1(G92gat), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT110), .ZN(G1337gat));
  OAI21_X1  g526(.A(G99gat), .B1(new_n720_), .B2(new_n262_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n714_), .A2(new_n410_), .A3(new_n617_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT51), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n728_), .A2(new_n732_), .A3(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1338gat));
  NAND3_X1  g533(.A1(new_n714_), .A2(new_n411_), .A3(new_n306_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n628_), .A2(new_n636_), .A3(new_n306_), .A4(new_n543_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n737_), .A2(new_n684_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n738_), .B2(G106gat), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n736_), .B(G106gat), .C1(new_n737_), .C2(new_n684_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n735_), .B1(new_n739_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT53), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT53), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n744_), .B(new_n735_), .C1(new_n739_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1339gat));
  INV_X1    g545(.A(KEYINPUT54), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n463_), .A2(new_n514_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n578_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n578_), .B2(new_n748_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT115), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT56), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n441_), .A2(new_n449_), .A3(new_n443_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n446_), .B2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n452_), .B2(new_n755_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n752_), .B(new_n753_), .C1(new_n757_), .C2(new_n403_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n755_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n754_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(KEYINPUT55), .B2(new_n450_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n403_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT115), .B1(new_n762_), .B2(KEYINPUT56), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT56), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n758_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n510_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n766_), .A2(KEYINPUT114), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n494_), .A2(new_n504_), .A3(new_n497_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(KEYINPUT114), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n767_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(new_n513_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(new_n458_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n765_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n576_), .A2(new_n577_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n765_), .A2(KEYINPUT58), .A3(new_n772_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT58), .B1(new_n765_), .B2(new_n772_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT116), .B1(new_n780_), .B2(new_n626_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(new_n779_), .A3(new_n781_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n458_), .A2(new_n514_), .A3(KEYINPUT111), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT111), .B1(new_n458_), .B2(new_n514_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n762_), .A2(KEYINPUT112), .A3(new_n786_), .A4(new_n753_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT113), .B1(new_n753_), .B2(KEYINPUT112), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(new_n762_), .B2(KEYINPUT56), .ZN(new_n789_));
  AOI211_X1 g588(.A(KEYINPUT113), .B(new_n403_), .C1(new_n759_), .C2(new_n761_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n785_), .B(new_n787_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n771_), .B1(new_n455_), .B2(new_n459_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT57), .B1(new_n793_), .B2(new_n588_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n795_), .B(new_n689_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n782_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n589_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n751_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n617_), .A2(new_n305_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n801_), .A2(new_n389_), .A3(new_n582_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT117), .B1(new_n800_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n589_), .B1(new_n782_), .B2(new_n797_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n805_), .B(new_n802_), .C1(new_n806_), .C2(new_n751_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n514_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  INV_X1    g609(.A(G113gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n515_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT118), .B1(new_n813_), .B2(G113gat), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n798_), .B2(new_n543_), .ZN(new_n816_));
  AOI211_X1 g615(.A(KEYINPUT119), .B(new_n645_), .C1(new_n782_), .C2(new_n797_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n751_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT59), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n800_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n802_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n820_), .A2(new_n802_), .B1(KEYINPUT59), .B2(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n515_), .A2(new_n811_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n812_), .A2(new_n814_), .B1(new_n823_), .B2(new_n824_), .ZN(G1340gat));
  NAND2_X1  g624(.A1(new_n798_), .A2(new_n543_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT119), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n798_), .A2(new_n815_), .A3(new_n543_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n819_), .A3(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n802_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n822_), .A2(KEYINPUT59), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n463_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G120gat), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT60), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n804_), .A2(new_n807_), .B1(new_n836_), .B2(G120gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(G120gat), .B1(new_n463_), .B2(new_n836_), .ZN(new_n838_));
  XOR2_X1   g637(.A(new_n838_), .B(KEYINPUT120), .Z(new_n839_));
  AOI21_X1  g638(.A(new_n835_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n836_), .A2(G120gat), .ZN(new_n841_));
  AND4_X1   g640(.A1(new_n835_), .A2(new_n808_), .A3(new_n841_), .A4(new_n839_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n834_), .B1(new_n840_), .B2(new_n842_), .ZN(G1341gat));
  AOI21_X1  g642(.A(new_n543_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n844_), .A2(G127gat), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n831_), .A2(new_n832_), .A3(G127gat), .A4(new_n589_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1342gat));
  AOI21_X1  g646(.A(new_n588_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n848_), .A2(G134gat), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n831_), .A2(new_n832_), .A3(G134gat), .A4(new_n777_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1343gat));
  NOR2_X1   g650(.A1(new_n617_), .A2(new_n305_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(new_n583_), .A3(new_n600_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT122), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n800_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n514_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n463_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n645_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT61), .B(G155gat), .Z(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT123), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n860_), .B(new_n862_), .ZN(G1346gat));
  NOR4_X1   g662(.A1(new_n800_), .A2(new_n546_), .A3(new_n626_), .A4(new_n854_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n855_), .A2(new_n689_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n546_), .B2(new_n865_), .ZN(G1347gat));
  NOR3_X1   g665(.A1(new_n583_), .A2(new_n801_), .A3(new_n600_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n829_), .A2(new_n514_), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n868_), .A2(new_n869_), .A3(G169gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n868_), .B2(G169gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n208_), .A2(new_n347_), .ZN(new_n872_));
  OAI22_X1  g671(.A1(new_n870_), .A2(new_n871_), .B1(new_n868_), .B2(new_n872_), .ZN(G1348gat));
  AND2_X1   g672(.A1(new_n821_), .A2(new_n867_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n874_), .A2(KEYINPUT124), .A3(G176gat), .A4(new_n463_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n821_), .A2(G176gat), .A3(new_n867_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n682_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n878_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n829_), .A2(new_n867_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n463_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n209_), .B2(new_n881_), .ZN(G1349gat));
  AOI21_X1  g681(.A(G183gat), .B1(new_n874_), .B2(new_n645_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n799_), .A2(new_n223_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n880_), .B2(new_n884_), .ZN(G1350gat));
  NAND2_X1  g684(.A1(new_n880_), .A2(new_n777_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G190gat), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n588_), .A2(new_n344_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n880_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1351gat));
  NOR2_X1   g689(.A1(new_n600_), .A2(new_n652_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n821_), .A2(new_n852_), .A3(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n515_), .ZN(new_n893_));
  AOI21_X1  g692(.A(KEYINPUT125), .B1(new_n893_), .B2(G197gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(G197gat), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n896_));
  NOR4_X1   g695(.A1(new_n892_), .A2(new_n896_), .A3(new_n509_), .A4(new_n515_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n894_), .A2(new_n895_), .A3(new_n897_), .ZN(G1352gat));
  INV_X1    g697(.A(new_n892_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n463_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g700(.A1(new_n892_), .A2(new_n799_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT126), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT127), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n906_), .A2(new_n907_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n904_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n902_), .A2(new_n907_), .A3(new_n906_), .A4(new_n903_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1354gat));
  AOI21_X1  g711(.A(G218gat), .B1(new_n899_), .B2(new_n689_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n892_), .A2(new_n626_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(G218gat), .B2(new_n914_), .ZN(G1355gat));
endmodule


