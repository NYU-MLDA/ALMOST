//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT36), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G29gat), .B(G36gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  AOI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT9), .A2(G92gat), .ZN(new_n218_));
  INV_X1    g017(.A(G85gat), .ZN(new_n219_));
  INV_X1    g018(.A(G92gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n218_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n224_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n217_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230_));
  INV_X1    g029(.A(G99gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(new_n215_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n213_), .B1(G99gat), .B2(G106gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n229_), .B(new_n232_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n236_));
  AND2_X1   g035(.A1(G85gat), .A2(G92gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n221_), .A2(KEYINPUT66), .A3(new_n222_), .ZN(new_n240_));
  AND4_X1   g039(.A1(new_n228_), .A2(new_n235_), .A3(new_n239_), .A4(new_n240_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n239_), .A2(new_n240_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n228_), .B1(new_n242_), .B2(new_n235_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n227_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n211_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G232gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT34), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT35), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n232_), .A2(new_n229_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n214_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n239_), .A2(new_n240_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT8), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n242_), .A2(new_n228_), .A3(new_n235_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(new_n209_), .A3(new_n227_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n245_), .A2(new_n250_), .A3(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n248_), .A2(new_n249_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n259_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n206_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n260_), .A2(new_n261_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n263_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G127gat), .B(G155gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT16), .ZN(new_n270_));
  XOR2_X1   g069(.A(G183gat), .B(G211gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G1gat), .B(G8gat), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G1gat), .ZN(new_n277_));
  INV_X1    g076(.A(G8gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT14), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  OR2_X1    g078(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(G22gat), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(G22gat), .B1(new_n280_), .B2(new_n281_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n279_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n285_), .A2(KEYINPUT74), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT73), .B(G15gat), .ZN(new_n288_));
  INV_X1    g087(.A(G22gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n282_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n287_), .B1(new_n291_), .B2(new_n279_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n276_), .B1(new_n286_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n285_), .A2(KEYINPUT74), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n291_), .A2(new_n287_), .A3(new_n279_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n275_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G231gat), .A2(G233gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n298_), .B(KEYINPUT75), .Z(new_n299_));
  OR2_X1    g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n299_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G64gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G57gat), .ZN(new_n304_));
  INV_X1    g103(.A(G57gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G64gat), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n304_), .A2(new_n306_), .A3(KEYINPUT67), .ZN(new_n307_));
  AOI21_X1  g106(.A(KEYINPUT67), .B1(new_n304_), .B2(new_n306_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT11), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT67), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n305_), .A2(G64gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n303_), .A2(G57gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT11), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n304_), .A2(new_n306_), .A3(KEYINPUT67), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G78gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G71gat), .ZN(new_n318_));
  INV_X1    g117(.A(G71gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G78gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n309_), .A2(new_n316_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n313_), .A2(new_n315_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n321_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(KEYINPUT11), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n302_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n302_), .A2(new_n326_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n274_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OAI211_X1 g131(.A(KEYINPUT77), .B(new_n274_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n272_), .B(KEYINPUT17), .Z(new_n334_));
  OR3_X1    g133(.A1(new_n328_), .A2(new_n329_), .A3(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n332_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G127gat), .B(G134gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G113gat), .B(G120gat), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n338_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT31), .ZN(new_n342_));
  AND3_X1   g141(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT26), .B(G190gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n351_));
  INV_X1    g150(.A(G183gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT25), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n352_), .A2(KEYINPUT25), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n350_), .B(new_n353_), .C1(new_n354_), .C2(new_n351_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n346_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(KEYINPUT24), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT80), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n356_), .A2(new_n360_), .A3(KEYINPUT24), .A4(new_n357_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n349_), .A2(new_n355_), .A3(new_n359_), .A4(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G169gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT22), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT22), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G169gat), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n368_));
  INV_X1    g167(.A(G176gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n344_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n372_));
  INV_X1    g171(.A(G190gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n352_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n364_), .A2(new_n366_), .A3(new_n369_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT81), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n370_), .A2(new_n357_), .A3(new_n375_), .A4(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n362_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G71gat), .B(G99gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(G43gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n379_), .B(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G227gat), .A2(G233gat), .ZN(new_n383_));
  INV_X1    g182(.A(G15gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT30), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n382_), .B(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n342_), .B1(new_n388_), .B2(KEYINPUT82), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(KEYINPUT82), .B2(new_n388_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G1gat), .B(G29gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(G85gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT0), .B(G57gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n392_), .B(new_n393_), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G225gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT93), .ZN(new_n397_));
  XOR2_X1   g196(.A(G155gat), .B(G162gat), .Z(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT84), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT3), .ZN(new_n401_));
  INV_X1    g200(.A(G141gat), .ZN(new_n402_));
  INV_X1    g201(.A(G148gat), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .A4(KEYINPUT83), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT83), .ZN(new_n405_));
  OAI22_X1  g204(.A1(new_n405_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT2), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G141gat), .A2(G148gat), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n404_), .B(new_n406_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n398_), .B1(new_n400_), .B2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(G155gat), .A2(G162gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G155gat), .A2(G162gat), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n411_), .B1(KEYINPUT1), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(KEYINPUT1), .B2(new_n412_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n402_), .A2(new_n403_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n408_), .A3(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n410_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n341_), .A2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n397_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n341_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n410_), .A2(new_n416_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT92), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n341_), .A2(new_n410_), .A3(new_n416_), .A4(KEYINPUT92), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n420_), .B1(new_n426_), .B2(KEYINPUT4), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n397_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n395_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n397_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n418_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n431_), .B(new_n394_), .C1(new_n432_), .C2(new_n420_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n388_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT82), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n342_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n390_), .A2(new_n435_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT25), .B(G183gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n350_), .A2(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n349_), .A2(new_n358_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT89), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n376_), .A2(new_n444_), .A3(new_n357_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n444_), .B1(new_n376_), .B2(new_n357_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n375_), .A2(KEYINPUT90), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT90), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n345_), .A2(new_n449_), .A3(new_n374_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT91), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n376_), .A2(new_n357_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT89), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n376_), .A2(new_n444_), .A3(new_n357_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AND4_X1   g255(.A1(new_n449_), .A2(new_n371_), .A3(new_n372_), .A4(new_n374_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n449_), .B1(new_n345_), .B2(new_n374_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT91), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n456_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n443_), .B1(new_n452_), .B2(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G197gat), .B(G204gat), .Z(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT21), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G197gat), .B(G204gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT21), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G211gat), .B(G218gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  OR3_X1    g268(.A1(new_n465_), .A2(new_n468_), .A3(new_n466_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n462_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G226gat), .A2(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  AOI211_X1 g276(.A(new_n474_), .B(new_n477_), .C1(new_n379_), .C2(new_n471_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT20), .B1(new_n379_), .B2(new_n471_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n443_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n447_), .A2(new_n451_), .A3(KEYINPUT91), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n460_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n480_), .B1(new_n484_), .B2(new_n471_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n477_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n479_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G8gat), .B(G36gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT18), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G64gat), .B(G92gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n362_), .A2(new_n378_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n474_), .B1(new_n494_), .B2(new_n472_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n462_), .B2(new_n472_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n496_), .A2(new_n477_), .B1(new_n473_), .B2(new_n478_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n491_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n500_));
  AOI211_X1 g299(.A(new_n471_), .B(new_n443_), .C1(new_n456_), .C2(new_n459_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT20), .B1(new_n494_), .B2(new_n472_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n477_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n503_), .B1(new_n477_), .B2(new_n496_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n492_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT27), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n506_), .B1(new_n497_), .B2(new_n491_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n499_), .A2(new_n500_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G78gat), .B(G106gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(KEYINPUT87), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n471_), .A2(KEYINPUT85), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n422_), .A2(KEYINPUT29), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G228gat), .A2(G233gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n515_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n511_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n515_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n422_), .A2(KEYINPUT29), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n521_), .B2(new_n512_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n522_), .B(new_n516_), .C1(KEYINPUT87), .C2(new_n510_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n422_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT28), .B1(new_n422_), .B2(KEYINPUT29), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G22gat), .B(G50gat), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n526_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n529_), .B1(new_n530_), .B2(new_n524_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n519_), .A2(new_n523_), .A3(new_n528_), .A4(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(KEYINPUT86), .B(new_n510_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n528_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n509_), .B(KEYINPUT86), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n522_), .A2(new_n516_), .A3(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n532_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT96), .B1(new_n508_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n496_), .A2(new_n477_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n540_), .A2(new_n491_), .A3(new_n479_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n491_), .B1(new_n540_), .B2(new_n479_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n500_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n507_), .A2(new_n505_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n543_), .A2(new_n538_), .A3(new_n544_), .A4(KEYINPUT96), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n440_), .B1(new_n539_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n390_), .A2(new_n438_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n532_), .A2(new_n537_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n543_), .A2(new_n544_), .A3(new_n435_), .A4(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT33), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n426_), .A2(KEYINPUT4), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n417_), .A2(new_n419_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(new_n397_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n394_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT94), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n426_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n424_), .A2(KEYINPUT94), .A3(new_n425_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n397_), .A3(new_n559_), .ZN(new_n560_));
  AOI22_X1  g359(.A1(new_n552_), .A2(new_n433_), .B1(new_n556_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n420_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n553_), .A2(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n563_), .A2(KEYINPUT33), .A3(new_n431_), .A4(new_n394_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n561_), .A2(new_n498_), .A3(new_n493_), .A4(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n491_), .A2(KEYINPUT32), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n504_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n497_), .A2(new_n566_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n434_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n549_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n548_), .B1(new_n551_), .B2(new_n571_), .ZN(new_n572_));
  AOI211_X1 g371(.A(new_n268_), .B(new_n336_), .C1(new_n547_), .C2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT68), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G230gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT64), .ZN(new_n576_));
  AOI211_X1 g375(.A(new_n314_), .B(new_n321_), .C1(new_n313_), .C2(new_n315_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n324_), .B1(new_n323_), .B2(KEYINPUT11), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n577_), .B1(new_n578_), .B2(new_n316_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n244_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n326_), .A2(new_n256_), .A3(new_n227_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(KEYINPUT12), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT12), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n244_), .A2(new_n583_), .A3(new_n579_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n576_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n576_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n574_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G120gat), .B(G148gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(G176gat), .B(G204gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n588_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n582_), .A2(new_n584_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n587_), .B1(new_n595_), .B2(new_n586_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT68), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n586_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n587_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n593_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT70), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT70), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n596_), .A2(new_n603_), .A3(new_n600_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n594_), .A2(new_n597_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT13), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT13), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n597_), .A2(new_n593_), .A3(new_n588_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n603_), .B1(new_n596_), .B2(new_n600_), .ZN(new_n609_));
  NOR4_X1   g408(.A1(new_n585_), .A2(KEYINPUT70), .A3(new_n587_), .A4(new_n593_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n607_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n606_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G113gat), .B(G141gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G169gat), .B(G197gat), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n614_), .B(new_n615_), .Z(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n297_), .A2(new_n211_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT78), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n209_), .B(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n293_), .A3(new_n296_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G229gat), .A2(G233gat), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n618_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n297_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n622_), .B1(new_n625_), .B2(new_n621_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n617_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n622_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n620_), .A2(new_n293_), .A3(new_n296_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n620_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n628_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n618_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n632_), .A3(new_n616_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n627_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n613_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n573_), .A2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G1gat), .B1(new_n637_), .B2(new_n435_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT38), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n547_), .A2(new_n572_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n634_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n613_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT37), .B1(new_n262_), .B2(KEYINPUT72), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n268_), .A2(new_n644_), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n267_), .B(KEYINPUT37), .C1(KEYINPUT72), .C2(new_n262_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n336_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n643_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n642_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n435_), .A2(G1gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(KEYINPUT97), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n654_));
  INV_X1    g453(.A(new_n652_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n650_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n657_), .B2(new_n639_), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT98), .B(KEYINPUT38), .C1(new_n653_), .C2(new_n656_), .ZN(new_n660_));
  OAI221_X1 g459(.A(new_n638_), .B1(new_n639_), .B2(new_n657_), .C1(new_n659_), .C2(new_n660_), .ZN(G1324gat));
  OAI21_X1  g460(.A(G8gat), .B1(new_n637_), .B2(new_n508_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT39), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n543_), .A2(new_n544_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n651_), .A2(new_n278_), .A3(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g466(.A(G15gat), .B1(new_n637_), .B2(new_n548_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT41), .Z(new_n669_));
  AND2_X1   g468(.A1(new_n390_), .A2(new_n438_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n651_), .A2(new_n384_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT99), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n669_), .A2(new_n674_), .A3(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1326gat));
  OAI21_X1  g475(.A(G22gat), .B1(new_n637_), .B2(new_n538_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT42), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n651_), .A2(new_n289_), .A3(new_n549_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1327gat));
  INV_X1    g479(.A(new_n336_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n613_), .A2(new_n681_), .A3(new_n267_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n642_), .A2(new_n682_), .ZN(new_n683_));
  OR3_X1    g482(.A1(new_n683_), .A2(G29gat), .A3(new_n435_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n613_), .A2(new_n681_), .A3(new_n635_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n267_), .B(new_n644_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n640_), .B2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n543_), .A2(new_n538_), .A3(new_n544_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT96), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n439_), .B1(new_n691_), .B2(new_n545_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n433_), .A2(new_n552_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n556_), .A2(new_n560_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n564_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n570_), .B1(new_n499_), .B2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n538_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n670_), .B1(new_n697_), .B2(new_n550_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n686_), .B(new_n687_), .C1(new_n692_), .C2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n685_), .B1(new_n688_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT44), .B(new_n685_), .C1(new_n688_), .C2(new_n700_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n434_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT100), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n705_), .A2(new_n706_), .A3(G29gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n705_), .B2(G29gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n684_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT101), .B(new_n684_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1328gat));
  INV_X1    g512(.A(G36gat), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n703_), .A2(new_n704_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(new_n664_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n683_), .A2(G36gat), .A3(new_n508_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT103), .Z(new_n719_));
  XNOR2_X1  g518(.A(new_n717_), .B(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(KEYINPUT104), .ZN(new_n722_));
  OR3_X1    g521(.A1(new_n716_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n716_), .B2(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1329gat));
  NAND3_X1  g524(.A1(new_n715_), .A2(G43gat), .A3(new_n670_), .ZN(new_n726_));
  INV_X1    g525(.A(G43gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n727_), .B1(new_n683_), .B2(new_n548_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g529(.A(new_n683_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G50gat), .B1(new_n731_), .B2(new_n549_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n549_), .A2(G50gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n715_), .B2(new_n733_), .ZN(G1331gat));
  AND2_X1   g533(.A1(new_n647_), .A2(new_n613_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT105), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n634_), .B1(new_n547_), .B2(new_n572_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  OR3_X1    g537(.A1(new_n736_), .A2(KEYINPUT106), .A3(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT106), .B1(new_n736_), .B2(new_n738_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n739_), .A2(new_n305_), .A3(new_n434_), .A4(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n643_), .A2(new_n634_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n573_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G57gat), .B1(new_n743_), .B2(new_n435_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n741_), .A2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT107), .ZN(G1332gat));
  OAI21_X1  g545(.A(G64gat), .B1(new_n743_), .B2(new_n508_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT108), .Z(new_n748_));
  OR2_X1    g547(.A1(new_n748_), .A2(KEYINPUT48), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(KEYINPUT48), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n739_), .A2(new_n740_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n508_), .A2(G64gat), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT109), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n749_), .B(new_n750_), .C1(new_n751_), .C2(new_n753_), .ZN(G1333gat));
  OAI21_X1  g553(.A(G71gat), .B1(new_n743_), .B2(new_n548_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT49), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n670_), .A2(new_n319_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n751_), .B2(new_n757_), .ZN(G1334gat));
  OAI21_X1  g557(.A(G78gat), .B1(new_n743_), .B2(new_n538_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT50), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n549_), .A2(new_n317_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n751_), .B2(new_n761_), .ZN(G1335gat));
  OR2_X1    g561(.A1(new_n688_), .A2(new_n700_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n613_), .A2(new_n635_), .A3(new_n336_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT110), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766_), .B2(new_n435_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n737_), .A2(new_n268_), .A3(new_n336_), .A4(new_n613_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n219_), .A3(new_n434_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n770_), .ZN(G1336gat));
  OAI21_X1  g570(.A(G92gat), .B1(new_n766_), .B2(new_n508_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(new_n220_), .A3(new_n664_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1337gat));
  OAI21_X1  g573(.A(G99gat), .B1(new_n766_), .B2(new_n548_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n769_), .A2(new_n670_), .A3(new_n216_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g577(.A1(new_n769_), .A2(new_n215_), .A3(new_n549_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n763_), .A2(new_n549_), .A3(new_n765_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  AND4_X1   g580(.A1(KEYINPUT111), .A2(new_n780_), .A3(new_n781_), .A4(G106gat), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n215_), .B1(new_n783_), .B2(KEYINPUT52), .ZN(new_n784_));
  AOI22_X1  g583(.A1(new_n780_), .A2(new_n784_), .B1(KEYINPUT111), .B2(new_n781_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n779_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n779_), .B(new_n787_), .C1(new_n782_), .C2(new_n785_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1339gat));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n622_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n618_), .A2(new_n621_), .A3(new_n628_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n617_), .A3(new_n794_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n633_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n792_), .B1(new_n605_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n634_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT113), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n634_), .B(new_n801_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n582_), .A2(new_n576_), .A3(new_n584_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n598_), .A2(KEYINPUT55), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n600_), .B1(new_n585_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n806_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n800_), .A2(new_n802_), .A3(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(KEYINPUT114), .B(new_n796_), .C1(new_n608_), .C2(new_n611_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n798_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n267_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n814_), .A2(KEYINPUT57), .A3(new_n267_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n807_), .A2(KEYINPUT117), .A3(new_n808_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n809_), .A2(new_n821_), .A3(new_n810_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n602_), .A2(new_n604_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT116), .B1(new_n823_), .B2(new_n796_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n796_), .B(KEYINPUT116), .C1(new_n609_), .C2(new_n610_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n820_), .B(new_n822_), .C1(new_n824_), .C2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n611_), .B2(new_n797_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n825_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n832_), .A2(KEYINPUT58), .A3(new_n820_), .A4(new_n822_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n829_), .A2(new_n687_), .A3(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n818_), .A2(new_n819_), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n816_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n336_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n643_), .A2(new_n647_), .A3(new_n635_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n841_), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n435_), .B(new_n548_), .C1(new_n691_), .C2(new_n545_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(G113gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n634_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n843_), .A2(new_n848_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n815_), .A2(new_n817_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(new_n819_), .A3(new_n834_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n336_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n840_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(KEYINPUT118), .A3(new_n336_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n850_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n849_), .A2(new_n857_), .A3(new_n635_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n847_), .B1(new_n858_), .B2(new_n846_), .ZN(G1340gat));
  NOR3_X1   g658(.A1(new_n849_), .A2(new_n857_), .A3(new_n643_), .ZN(new_n860_));
  INV_X1    g659(.A(G120gat), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT60), .ZN(new_n862_));
  AOI21_X1  g661(.A(G120gat), .B1(new_n613_), .B2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n861_), .A2(KEYINPUT60), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT119), .B1(new_n845_), .B2(new_n865_), .ZN(new_n866_));
  AND4_X1   g665(.A1(KEYINPUT119), .A2(new_n842_), .A3(new_n843_), .A4(new_n865_), .ZN(new_n867_));
  OAI22_X1  g666(.A1(new_n860_), .A2(new_n861_), .B1(new_n866_), .B2(new_n867_), .ZN(G1341gat));
  INV_X1    g667(.A(G127gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n845_), .A2(new_n869_), .A3(new_n681_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n849_), .A2(new_n857_), .A3(new_n336_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n869_), .ZN(G1342gat));
  AOI21_X1  g671(.A(G134gat), .B1(new_n845_), .B2(new_n268_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n849_), .A2(new_n857_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n687_), .A2(G134gat), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT120), .Z(new_n876_));
  AOI21_X1  g675(.A(new_n873_), .B1(new_n874_), .B2(new_n876_), .ZN(G1343gat));
  NOR4_X1   g676(.A1(new_n670_), .A2(new_n664_), .A3(new_n435_), .A4(new_n538_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n837_), .B2(new_n841_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n634_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n613_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g683(.A1(new_n880_), .A2(new_n681_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT61), .B(G155gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1346gat));
  INV_X1    g686(.A(G162gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(new_n880_), .B2(new_n687_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n267_), .A2(G162gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n880_), .A2(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n890_), .A2(KEYINPUT121), .A3(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n894_));
  INV_X1    g693(.A(new_n892_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n889_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n893_), .A2(new_n896_), .ZN(G1347gat));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n439_), .A2(new_n508_), .A3(new_n549_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n635_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n898_), .B(new_n899_), .C1(new_n904_), .C2(new_n363_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n367_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n853_), .A2(new_n854_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n907_), .A2(new_n841_), .A3(new_n856_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n363_), .B1(new_n908_), .B2(new_n902_), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT62), .B1(new_n909_), .B2(KEYINPUT122), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n904_), .A2(new_n898_), .A3(new_n363_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n905_), .B(new_n906_), .C1(new_n910_), .C2(new_n911_), .ZN(G1348gat));
  AOI21_X1  g711(.A(new_n549_), .B1(new_n837_), .B2(new_n841_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n439_), .A2(new_n508_), .ZN(new_n914_));
  AND4_X1   g713(.A1(G176gat), .A2(new_n913_), .A3(new_n613_), .A4(new_n914_), .ZN(new_n915_));
  AOI211_X1 g714(.A(new_n643_), .B(new_n901_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n916_));
  OAI21_X1  g715(.A(KEYINPUT123), .B1(new_n916_), .B2(G176gat), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n901_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n613_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n919_), .A2(new_n920_), .A3(new_n369_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n915_), .B1(new_n917_), .B2(new_n921_), .ZN(G1349gat));
  NAND3_X1  g721(.A1(new_n913_), .A2(new_n681_), .A3(new_n914_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n336_), .A2(new_n441_), .ZN(new_n924_));
  AOI22_X1  g723(.A1(new_n923_), .A2(new_n352_), .B1(new_n918_), .B2(new_n924_), .ZN(G1350gat));
  NAND2_X1  g724(.A1(new_n268_), .A2(new_n350_), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT124), .Z(new_n927_));
  NAND2_X1  g726(.A1(new_n918_), .A2(new_n927_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n918_), .A2(new_n687_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n373_), .ZN(G1351gat));
  NAND4_X1  g729(.A1(new_n548_), .A2(new_n664_), .A3(new_n435_), .A4(new_n549_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n931_), .B1(new_n837_), .B2(new_n841_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n634_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n613_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g735(.A(new_n336_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n937_));
  XOR2_X1   g736(.A(new_n937_), .B(KEYINPUT125), .Z(new_n938_));
  NAND2_X1  g737(.A1(new_n932_), .A2(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(KEYINPUT126), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(KEYINPUT127), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n939_), .B(new_n942_), .ZN(G1354gat));
  INV_X1    g742(.A(G218gat), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n932_), .A2(new_n944_), .A3(new_n268_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n932_), .A2(new_n687_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n946_), .B2(new_n944_), .ZN(G1355gat));
endmodule


