//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT65), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(KEYINPUT9), .B2(G85gat), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n204_), .B(new_n209_), .C1(new_n211_), .C2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G99gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(new_n203_), .A3(KEYINPUT66), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT7), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n221_), .A2(new_n218_), .A3(new_n203_), .A4(KEYINPUT66), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n209_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n212_), .A2(G85gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n214_), .A2(G92gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n223_), .A2(new_n224_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n224_), .B1(new_n223_), .B2(new_n228_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n217_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G29gat), .B(G36gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G43gat), .B(G50gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n233_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(KEYINPUT15), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n235_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT15), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n231_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n223_), .A2(new_n228_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT8), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n223_), .A2(new_n224_), .A3(new_n228_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(new_n237_), .A3(new_n217_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G232gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT34), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT35), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT72), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n240_), .A2(new_n245_), .A3(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n248_), .A2(new_n249_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G190gat), .B(G218gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT71), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G134gat), .B(G162gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n255_), .A2(new_n257_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT36), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n252_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n240_), .A2(new_n264_), .A3(new_n245_), .A4(new_n250_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n253_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT73), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT73), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n253_), .A2(new_n268_), .A3(new_n263_), .A4(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT75), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n253_), .A2(new_n265_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n263_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n260_), .A2(KEYINPUT36), .A3(new_n262_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT74), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n274_), .A2(new_n275_), .A3(KEYINPUT74), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n273_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n270_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n272_), .A2(new_n281_), .A3(KEYINPUT37), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT37), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n270_), .B(new_n280_), .C1(new_n271_), .C2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G231gat), .A2(G233gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT17), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G127gat), .B(G155gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT16), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G183gat), .B(G211gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT16), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n289_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n291_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n288_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT77), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n287_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G57gat), .B(G64gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G71gat), .B(G78gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n302_), .A3(KEYINPUT11), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(KEYINPUT11), .ZN(new_n304_));
  INV_X1    g103(.A(new_n302_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n301_), .A2(KEYINPUT11), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n303_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n297_), .A2(new_n298_), .A3(new_n287_), .ZN(new_n309_));
  NOR3_X1   g108(.A1(new_n300_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n308_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n309_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(new_n299_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G1gat), .B(G8gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT76), .ZN(new_n315_));
  OR2_X1    g114(.A1(G15gat), .A2(G22gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G15gat), .A2(G22gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G1gat), .A2(G8gat), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n316_), .A2(new_n317_), .B1(KEYINPUT14), .B2(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(G1gat), .A2(G8gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(new_n318_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n315_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n319_), .B1(new_n315_), .B2(new_n322_), .ZN(new_n324_));
  OAI22_X1  g123(.A1(new_n310_), .A2(new_n313_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n308_), .B1(new_n300_), .B2(new_n309_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n312_), .A2(new_n311_), .A3(new_n299_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n323_), .A2(new_n324_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n292_), .A2(new_n296_), .A3(new_n288_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n325_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT78), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT78), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n325_), .A2(new_n329_), .A3(new_n333_), .A4(new_n330_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G120gat), .B(G148gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT5), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G176gat), .B(G204gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT12), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(KEYINPUT68), .A2(KEYINPUT12), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n231_), .A2(new_n311_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n217_), .B(new_n308_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G230gat), .A2(G233gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n349_), .B(KEYINPUT64), .Z(new_n350_));
  AOI21_X1  g149(.A(new_n343_), .B1(new_n231_), .B2(new_n311_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n350_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n353_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n340_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n308_), .B1(new_n244_), .B2(new_n217_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n347_), .ZN(new_n357_));
  OAI22_X1  g156(.A1(new_n356_), .A2(new_n357_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n351_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(new_n353_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n354_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n340_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT69), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n355_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(KEYINPUT69), .B(new_n340_), .C1(new_n352_), .C2(new_n354_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT70), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT13), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n365_), .A2(new_n366_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n369_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  AND4_X1   g173(.A1(new_n285_), .A2(new_n336_), .A3(new_n370_), .A4(new_n374_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n375_), .A2(KEYINPUT79), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n328_), .A2(new_n239_), .A3(new_n236_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G229gat), .A2(G233gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n237_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n322_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n321_), .B1(new_n320_), .B2(new_n318_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n316_), .A2(new_n317_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n318_), .A2(KEYINPUT14), .ZN(new_n386_));
  OAI22_X1  g185(.A1(new_n383_), .A2(new_n384_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n315_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n235_), .A4(new_n234_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n380_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n379_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n237_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n328_), .A2(KEYINPUT80), .A3(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n391_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n391_), .A2(KEYINPUT81), .A3(new_n394_), .A4(new_n392_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n382_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G113gat), .B(G141gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G169gat), .B(G197gat), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n400_), .B(new_n401_), .Z(new_n402_));
  AOI21_X1  g201(.A(new_n377_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n404_));
  OR3_X1    g203(.A1(new_n399_), .A2(KEYINPUT82), .A3(new_n402_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G78gat), .B(G106gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G211gat), .B(G218gat), .Z(new_n409_));
  AND2_X1   g208(.A1(new_n409_), .A2(KEYINPUT21), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT93), .ZN(new_n411_));
  INV_X1    g210(.A(G204gat), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n411_), .B1(new_n412_), .B2(G197gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(G197gat), .ZN(new_n414_));
  INV_X1    g213(.A(G197gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(KEYINPUT93), .A3(G204gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n413_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n410_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT21), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n413_), .A2(new_n416_), .A3(new_n419_), .A4(new_n414_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT94), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n415_), .A2(G204gat), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n419_), .B1(new_n423_), .B2(new_n414_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(new_n409_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n420_), .A2(new_n421_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n418_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT2), .ZN(new_n429_));
  INV_X1    g228(.A(G141gat), .ZN(new_n430_));
  INV_X1    g229(.A(G148gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(G141gat), .A2(G148gat), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT3), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n432_), .A2(new_n435_), .A3(new_n436_), .A4(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G155gat), .A2(G162gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(G155gat), .A2(G162gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n438_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(KEYINPUT1), .B2(new_n439_), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n439_), .A2(KEYINPUT1), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n430_), .A2(new_n431_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n446_), .A2(new_n433_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n442_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT29), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n428_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G228gat), .A2(G233gat), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n452_), .B(KEYINPUT92), .Z(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n428_), .A2(new_n450_), .A3(new_n453_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n408_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(new_n408_), .A3(new_n456_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n449_), .A2(KEYINPUT29), .ZN(new_n461_));
  XOR2_X1   g260(.A(G22gat), .B(G50gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT28), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n461_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT95), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n464_), .B1(new_n457_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n460_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n458_), .A2(new_n465_), .A3(new_n459_), .A4(new_n464_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT27), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT99), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G169gat), .A2(G176gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT87), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT22), .B(G169gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n475_), .A2(KEYINPUT88), .ZN(new_n476_));
  INV_X1    g275(.A(G169gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT88), .B1(new_n477_), .B2(KEYINPUT22), .ZN(new_n478_));
  INV_X1    g277(.A(G176gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n474_), .B1(new_n476_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT89), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G183gat), .A2(G190gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT23), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT83), .B(G183gat), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n488_), .A2(G190gat), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n481_), .A2(new_n482_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(KEYINPUT89), .B(new_n474_), .C1(new_n476_), .C2(new_n480_), .ZN(new_n491_));
  OAI21_X1  g290(.A(G183gat), .B1(KEYINPUT85), .B2(KEYINPUT25), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT25), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT86), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT26), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(new_n498_), .B2(G190gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(KEYINPUT26), .B(G190gat), .Z(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(new_n500_), .B2(new_n497_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT83), .B(G183gat), .Z(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT84), .B1(new_n502_), .B2(KEYINPUT25), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT84), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n488_), .A2(new_n504_), .A3(new_n495_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n496_), .B(new_n501_), .C1(new_n503_), .C2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n477_), .A2(new_n479_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n485_), .B(new_n486_), .C1(new_n507_), .C2(KEYINPUT24), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(KEYINPUT24), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n508_), .B1(new_n510_), .B2(new_n474_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n490_), .A2(new_n491_), .B1(new_n506_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n428_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n472_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n481_), .A2(new_n482_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n489_), .A2(new_n487_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n491_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n506_), .A2(new_n511_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(KEYINPUT99), .A3(new_n428_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G226gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT19), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT20), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n508_), .B(KEYINPUT97), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT26), .B(G190gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT25), .B(G183gat), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n510_), .A2(new_n473_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT98), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n475_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n475_), .A2(new_n529_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n479_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT87), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n473_), .B(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(G183gat), .A2(G190gat), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n487_), .B2(new_n535_), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n525_), .A2(new_n528_), .B1(new_n532_), .B2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n524_), .B1(new_n513_), .B2(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n514_), .A2(new_n520_), .A3(new_n523_), .A4(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n508_), .A2(KEYINPUT97), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n508_), .A2(KEYINPUT97), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n528_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n532_), .A2(new_n536_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n524_), .B1(new_n544_), .B2(new_n428_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n513_), .A2(new_n518_), .A3(new_n517_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n522_), .B(KEYINPUT96), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(G8gat), .B(G36gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT18), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G64gat), .B(G92gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n539_), .A2(new_n549_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n539_), .B2(new_n549_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n471_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n548_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n545_), .A2(new_n546_), .A3(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n514_), .A2(new_n520_), .A3(new_n538_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n559_), .B1(new_n560_), .B2(new_n522_), .ZN(new_n561_));
  OAI211_X1 g360(.A(KEYINPUT27), .B(new_n554_), .C1(new_n561_), .C2(new_n553_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n470_), .A2(new_n557_), .A3(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G71gat), .B(G99gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(G43gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G227gat), .A2(G233gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(G15gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n565_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n512_), .A2(KEYINPUT30), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT30), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n519_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT90), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n569_), .A2(new_n571_), .A3(KEYINPUT90), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n568_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n568_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n578_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G113gat), .B(G120gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G127gat), .B(G134gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT91), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n583_), .A2(KEYINPUT91), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n582_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n583_), .A2(KEYINPUT91), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n584_), .A3(new_n581_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT31), .Z(new_n591_));
  NAND3_X1  g390(.A1(new_n577_), .A2(new_n580_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n591_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n576_), .B2(new_n579_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G1gat), .B(G29gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(G85gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT0), .B(G57gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n596_), .B(new_n597_), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G225gat), .A2(G233gat), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n585_), .A2(new_n586_), .A3(new_n582_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n581_), .B1(new_n588_), .B2(new_n584_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n449_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n587_), .A2(new_n589_), .A3(new_n448_), .A4(new_n442_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n601_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n604_), .A2(new_n605_), .A3(KEYINPUT4), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT4), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n590_), .A2(new_n609_), .A3(new_n449_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n599_), .B(new_n607_), .C1(new_n611_), .C2(new_n600_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n600_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n598_), .B1(new_n613_), .B2(new_n606_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n592_), .A2(new_n594_), .A3(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n563_), .A2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n592_), .A2(new_n594_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n539_), .A2(new_n549_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n553_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  OAI211_X1 g421(.A(KEYINPUT33), .B(new_n598_), .C1(new_n613_), .C2(new_n606_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n608_), .A2(new_n600_), .A3(new_n610_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n604_), .A2(new_n605_), .A3(new_n601_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n599_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT33), .B1(new_n624_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n614_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n622_), .A2(new_n554_), .A3(new_n623_), .A4(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n553_), .A2(KEYINPUT32), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n539_), .A2(new_n549_), .A3(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n615_), .B(new_n631_), .C1(new_n561_), .C2(new_n630_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n470_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n615_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n557_), .A2(new_n635_), .A3(new_n562_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n619_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n618_), .B1(new_n637_), .B2(KEYINPUT100), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n592_), .A2(new_n594_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n557_), .A2(new_n635_), .A3(new_n562_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n469_), .B1(new_n629_), .B2(new_n632_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n639_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n406_), .B1(new_n638_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n375_), .A2(KEYINPUT79), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n376_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n647_), .A2(G1gat), .A3(new_n616_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(KEYINPUT38), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT102), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n370_), .A2(new_n374_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n331_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n651_), .A2(new_n406_), .A3(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT101), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n270_), .A2(new_n280_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n638_), .B2(new_n644_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n654_), .A2(new_n615_), .A3(new_n656_), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n648_), .A2(KEYINPUT38), .B1(new_n657_), .B2(G1gat), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n650_), .A2(new_n658_), .ZN(G1324gat));
  NAND2_X1  g458(.A1(new_n557_), .A2(new_n562_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n654_), .A2(new_n660_), .A3(new_n656_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n662_));
  INV_X1    g461(.A(G8gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(KEYINPUT103), .B2(KEYINPUT39), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n661_), .A2(new_n662_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n662_), .B1(new_n661_), .B2(new_n664_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n660_), .A2(new_n663_), .ZN(new_n668_));
  OAI22_X1  g467(.A1(new_n666_), .A2(new_n667_), .B1(new_n647_), .B2(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g469(.A1(new_n654_), .A2(new_n656_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G15gat), .B1(new_n671_), .B2(new_n639_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n673_), .ZN(new_n675_));
  OR3_X1    g474(.A1(new_n647_), .A2(G15gat), .A3(new_n639_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n674_), .A2(new_n675_), .A3(new_n676_), .ZN(G1326gat));
  OAI21_X1  g476(.A(G22gat), .B1(new_n671_), .B2(new_n470_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT42), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n470_), .A2(G22gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n647_), .B2(new_n680_), .ZN(G1327gat));
  AOI21_X1  g480(.A(new_n285_), .B1(new_n638_), .B2(new_n644_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n651_), .A2(new_n406_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n285_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT100), .B(new_n639_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n618_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n634_), .A2(new_n636_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT100), .B1(new_n690_), .B2(new_n639_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n686_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(KEYINPUT105), .A3(new_n693_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n684_), .A2(new_n335_), .A3(new_n685_), .A4(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n692_), .A2(KEYINPUT105), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n336_), .B1(new_n698_), .B2(KEYINPUT43), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n699_), .A2(KEYINPUT44), .A3(new_n685_), .A4(new_n694_), .ZN(new_n700_));
  AND4_X1   g499(.A1(G29gat), .A2(new_n697_), .A3(new_n615_), .A4(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n651_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n336_), .A2(new_n281_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n645_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G29gat), .B1(new_n705_), .B2(new_n615_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n701_), .A2(new_n706_), .ZN(G1328gat));
  NAND3_X1  g506(.A1(new_n697_), .A2(new_n660_), .A3(new_n700_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G36gat), .ZN(new_n709_));
  INV_X1    g508(.A(new_n660_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n704_), .A2(G36gat), .A3(new_n710_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT45), .Z(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n709_), .A2(new_n712_), .A3(KEYINPUT46), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  NAND4_X1  g516(.A1(new_n697_), .A2(new_n700_), .A3(G43gat), .A4(new_n619_), .ZN(new_n718_));
  INV_X1    g517(.A(G43gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n704_), .B2(new_n639_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT47), .ZN(G1330gat));
  AND4_X1   g521(.A1(G50gat), .A2(new_n697_), .A3(new_n469_), .A4(new_n700_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G50gat), .B1(new_n705_), .B2(new_n469_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1331gat));
  NAND4_X1  g524(.A1(new_n656_), .A2(new_n406_), .A3(new_n336_), .A4(new_n651_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G57gat), .B1(new_n726_), .B2(new_n616_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n406_), .ZN(new_n728_));
  AOI211_X1 g527(.A(new_n728_), .B(new_n702_), .C1(new_n638_), .C2(new_n644_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n335_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n616_), .A2(G57gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(G1332gat));
  OAI21_X1  g532(.A(G64gat), .B1(new_n726_), .B2(new_n710_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT48), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n710_), .A2(G64gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n731_), .B2(new_n736_), .ZN(G1333gat));
  OAI21_X1  g536(.A(G71gat), .B1(new_n726_), .B2(new_n639_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT49), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n639_), .A2(G71gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n731_), .B2(new_n740_), .ZN(G1334gat));
  OAI21_X1  g540(.A(G78gat), .B1(new_n726_), .B2(new_n470_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT50), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n470_), .A2(G78gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n731_), .B2(new_n744_), .ZN(G1335gat));
  NAND2_X1  g544(.A1(new_n729_), .A2(new_n703_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n214_), .A3(new_n615_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n702_), .A2(new_n728_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n684_), .A2(new_n335_), .A3(new_n694_), .A4(new_n749_), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n750_), .A2(KEYINPUT106), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(KEYINPUT106), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n751_), .A2(new_n615_), .A3(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n748_), .B1(new_n753_), .B2(new_n214_), .ZN(G1336gat));
  NAND2_X1  g553(.A1(new_n660_), .A2(G92gat), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT107), .Z(new_n756_));
  NAND3_X1  g555(.A1(new_n751_), .A2(new_n752_), .A3(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n212_), .B1(new_n746_), .B2(new_n710_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1337gat));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n619_), .A2(new_n202_), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n746_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n746_), .B2(new_n761_), .ZN(new_n763_));
  AOI22_X1  g562(.A1(new_n762_), .A2(new_n763_), .B1(KEYINPUT109), .B2(KEYINPUT51), .ZN(new_n764_));
  OR2_X1    g563(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n765_));
  OAI21_X1  g564(.A(G99gat), .B1(new_n750_), .B2(new_n639_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1338gat));
  NAND3_X1  g568(.A1(new_n747_), .A2(new_n203_), .A3(new_n469_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(G106gat), .C1(new_n750_), .C2(new_n470_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n699_), .A2(new_n469_), .A3(new_n694_), .A4(new_n749_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n771_), .B1(new_n774_), .B2(G106gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n770_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT53), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n770_), .C1(new_n773_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1339gat));
  INV_X1    g579(.A(G113gat), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n563_), .A2(new_n639_), .A3(new_n616_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n378_), .A2(new_n392_), .A3(new_n380_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n391_), .A2(new_n379_), .A3(new_n394_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n402_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n785_), .A2(KEYINPUT111), .A3(new_n786_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n784_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n791_), .A2(new_n792_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n363_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n353_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n360_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NOR4_X1   g598(.A1(new_n348_), .A2(new_n798_), .A3(new_n351_), .A4(new_n350_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n796_), .B(new_n362_), .C1(new_n799_), .C2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n350_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n352_), .B1(KEYINPUT55), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n340_), .B1(new_n804_), .B2(new_n800_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n796_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n802_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(KEYINPUT114), .A3(new_n796_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n795_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n783_), .B(new_n686_), .C1(new_n810_), .C2(KEYINPUT58), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n362_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n807_), .B1(new_n812_), .B2(KEYINPUT56), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(KEYINPUT56), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n809_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n795_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT58), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT115), .B1(new_n817_), .B2(new_n285_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n810_), .A2(KEYINPUT58), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n811_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n404_), .A2(new_n405_), .A3(new_n363_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n812_), .A2(KEYINPUT56), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n802_), .ZN(new_n824_));
  AND4_X1   g623(.A1(new_n366_), .A2(new_n793_), .A3(new_n794_), .A4(new_n365_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n655_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n821_), .B1(new_n827_), .B2(KEYINPUT113), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n806_), .A2(new_n814_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n825_), .B1(new_n830_), .B2(new_n822_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n829_), .B(KEYINPUT57), .C1(new_n831_), .C2(new_n655_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n828_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n331_), .B1(new_n820_), .B2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n730_), .A2(new_n406_), .A3(new_n370_), .A4(new_n374_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT110), .B1(new_n835_), .B2(KEYINPUT54), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT110), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n375_), .A2(new_n837_), .A3(new_n838_), .A4(new_n406_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n835_), .A2(KEYINPUT54), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n836_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n782_), .B1(new_n834_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n781_), .B1(new_n842_), .B2(new_n406_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n843_), .A2(KEYINPUT116), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n336_), .B1(new_n820_), .B2(new_n833_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n845_), .A2(new_n841_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .A4(new_n782_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n845_), .A2(new_n841_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n782_), .A2(new_n848_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT117), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n842_), .A2(KEYINPUT59), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n406_), .A2(new_n781_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n849_), .A2(new_n852_), .A3(new_n853_), .A4(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n843_), .A2(KEYINPUT116), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n844_), .A2(new_n855_), .A3(new_n856_), .ZN(G1340gat));
  XNOR2_X1  g656(.A(KEYINPUT118), .B(G120gat), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n849_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n842_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT60), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n702_), .B2(new_n859_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n651_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n859_), .B1(new_n860_), .B2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1341gat));
  OAI21_X1  g667(.A(G127gat), .B1(new_n860_), .B2(new_n652_), .ZN(new_n869_));
  OR3_X1    g668(.A1(new_n842_), .A2(G127gat), .A3(new_n335_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1342gat));
  INV_X1    g670(.A(new_n860_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n686_), .A2(G134gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT120), .ZN(new_n874_));
  INV_X1    g673(.A(G134gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n842_), .B2(new_n281_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n877_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n872_), .A2(new_n874_), .B1(new_n878_), .B2(new_n879_), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n619_), .A2(new_n470_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n660_), .A2(new_n616_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n881_), .B(new_n882_), .C1(new_n834_), .C2(new_n841_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n883_), .A2(KEYINPUT121), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(KEYINPUT121), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G141gat), .B1(new_n886_), .B2(new_n406_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n430_), .B(new_n728_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1344gat));
  OAI21_X1  g688(.A(G148gat), .B1(new_n886_), .B2(new_n702_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n431_), .B(new_n651_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1345gat));
  XNOR2_X1  g691(.A(KEYINPUT61), .B(G155gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n893_), .B1(new_n886_), .B2(new_n335_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n893_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n336_), .B(new_n895_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1346gat));
  OAI21_X1  g696(.A(G162gat), .B1(new_n886_), .B2(new_n285_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n281_), .A2(G162gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1347gat));
  NOR4_X1   g700(.A1(new_n710_), .A2(new_n639_), .A3(new_n615_), .A4(new_n469_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n902_), .A2(new_n728_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n845_), .B2(new_n841_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT122), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n906_), .B(new_n903_), .C1(new_n845_), .C2(new_n841_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n905_), .A2(G169gat), .A3(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n477_), .B1(new_n904_), .B2(KEYINPUT122), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(KEYINPUT123), .A3(new_n907_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n910_), .A2(KEYINPUT62), .A3(new_n912_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n846_), .A2(new_n530_), .A3(new_n531_), .A4(new_n903_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(KEYINPUT123), .B1(new_n911_), .B2(new_n907_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n913_), .A2(new_n918_), .ZN(G1348gat));
  OR2_X1    g718(.A1(new_n834_), .A2(new_n841_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n920_), .A2(new_n902_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n702_), .A2(new_n479_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n846_), .A2(new_n651_), .A3(new_n902_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n921_), .A2(new_n922_), .B1(new_n923_), .B2(new_n479_), .ZN(G1349gat));
  NAND3_X1  g723(.A1(new_n920_), .A2(new_n336_), .A3(new_n902_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n502_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n652_), .A2(new_n527_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n846_), .A2(new_n902_), .A3(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n926_), .A2(KEYINPUT124), .A3(new_n928_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1350gat));
  NAND3_X1  g732(.A1(new_n846_), .A2(new_n686_), .A3(new_n902_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(G190gat), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n846_), .A2(new_n526_), .A3(new_n655_), .A4(new_n902_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n935_), .A2(KEYINPUT125), .A3(new_n936_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1351gat));
  NOR2_X1   g740(.A1(new_n710_), .A2(new_n615_), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n881_), .B(new_n942_), .C1(new_n834_), .C2(new_n841_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n943_), .A2(new_n406_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(new_n415_), .ZN(G1352gat));
  NOR2_X1   g744(.A1(new_n943_), .A2(new_n702_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(new_n412_), .ZN(G1353gat));
  AOI21_X1  g746(.A(new_n652_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  OR3_X1    g748(.A1(new_n943_), .A2(KEYINPUT126), .A3(new_n949_), .ZN(new_n950_));
  OAI21_X1  g749(.A(KEYINPUT126), .B1(new_n943_), .B2(new_n949_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n953_));
  INV_X1    g752(.A(G211gat), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n952_), .A2(new_n955_), .ZN(new_n956_));
  NAND4_X1  g755(.A1(new_n950_), .A2(new_n953_), .A3(new_n954_), .A4(new_n951_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1354gat));
  OR3_X1    g757(.A1(new_n943_), .A2(G218gat), .A3(new_n281_), .ZN(new_n959_));
  OAI21_X1  g758(.A(G218gat), .B1(new_n943_), .B2(new_n285_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(KEYINPUT127), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n959_), .A2(new_n963_), .A3(new_n960_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n962_), .A2(new_n964_), .ZN(G1355gat));
endmodule


