//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n910_, new_n912_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  INV_X1    g002(.A(G113gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G120gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G141gat), .ZN(new_n208_));
  INV_X1    g007(.A(G148gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT87), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT1), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n210_), .B(new_n211_), .C1(new_n214_), .C2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n210_), .A2(KEYINPUT3), .ZN(new_n218_));
  OR3_X1    g017(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n211_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n218_), .A2(new_n219_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n212_), .B(KEYINPUT87), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n215_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n207_), .A2(new_n217_), .A3(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n205_), .B(G120gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n217_), .A2(new_n225_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n226_), .A2(new_n229_), .A3(KEYINPUT4), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G225gat), .A2(G233gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n230_), .B(new_n232_), .C1(KEYINPUT4), .C2(new_n229_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n226_), .A2(new_n229_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(KEYINPUT93), .A3(new_n231_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n226_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT93), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n233_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT0), .B(G57gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G85gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(G1gat), .B(G29gat), .Z(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n243_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n233_), .A2(new_n235_), .A3(new_n238_), .A4(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G85gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(G92gat), .ZN(new_n249_));
  INV_X1    g048(.A(G92gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(G85gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT7), .ZN(new_n253_));
  INV_X1    g052(.A(G99gat), .ZN(new_n254_));
  INV_X1    g053(.A(G106gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AND3_X1   g057(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n252_), .B1(new_n258_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT8), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n256_), .A2(new_n257_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT66), .B1(new_n259_), .B2(new_n260_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G99gat), .A2(G106gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n269_));
  NAND3_X1  g068(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n264_), .B1(new_n265_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n250_), .A2(G85gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n248_), .A2(G92gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n263_), .ZN(new_n276_));
  OAI22_X1  g075(.A1(new_n262_), .A2(new_n263_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(KEYINPUT10), .B(G99gat), .Z(new_n278_));
  AOI22_X1  g077(.A1(new_n265_), .A2(new_n271_), .B1(new_n278_), .B2(new_n255_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT9), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(KEYINPUT64), .A3(G85gat), .ZN(new_n281_));
  OR2_X1    g080(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n250_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n280_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT65), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n286_), .A2(KEYINPUT9), .ZN(new_n287_));
  NOR2_X1   g086(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(G92gat), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT9), .B1(new_n249_), .B2(new_n251_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n279_), .A2(new_n285_), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G57gat), .ZN(new_n294_));
  INV_X1    g093(.A(G64gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT11), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G57gat), .A2(G64gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT67), .ZN(new_n300_));
  INV_X1    g099(.A(G71gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G78gat), .ZN(new_n302_));
  INV_X1    g101(.A(G78gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G71gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n299_), .A2(new_n300_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n300_), .B1(new_n299_), .B2(new_n305_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n297_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n307_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(G57gat), .A2(G64gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G57gat), .A2(G64gat), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT11), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G71gat), .B(G78gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT67), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n309_), .B1(new_n316_), .B2(new_n306_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n277_), .B(new_n293_), .C1(new_n311_), .C2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G230gat), .A2(G233gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(KEYINPUT69), .A3(new_n319_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n316_), .A2(new_n309_), .A3(new_n306_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n310_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n279_), .A2(new_n285_), .A3(new_n292_), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n259_), .A2(new_n260_), .A3(KEYINPUT66), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n269_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n258_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n276_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n268_), .A2(new_n270_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n275_), .B1(new_n264_), .B2(new_n332_), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n330_), .A2(new_n331_), .B1(new_n333_), .B2(KEYINPUT8), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n325_), .B(new_n326_), .C1(new_n327_), .C2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(new_n327_), .B2(new_n334_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(KEYINPUT12), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n326_), .A2(new_n325_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n277_), .A2(new_n293_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT12), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n340_), .B(new_n341_), .C1(new_n336_), .C2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n338_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n324_), .A2(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n335_), .A2(new_n318_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n345_), .B1(new_n319_), .B2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G120gat), .B(G148gat), .ZN(new_n348_));
  INV_X1    g147(.A(G204gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT5), .ZN(new_n351_));
  INV_X1    g150(.A(G176gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n347_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT13), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT37), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G232gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT34), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT35), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT70), .B(G43gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G50gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(G29gat), .B(G36gat), .Z(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(G50gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n363_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n365_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n371_), .A2(new_n341_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n366_), .A2(new_n370_), .ZN(new_n374_));
  XOR2_X1   g173(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n366_), .A2(new_n370_), .A3(new_n375_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n379_), .A2(KEYINPUT72), .A3(new_n341_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT72), .B1(new_n379_), .B2(new_n341_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n362_), .B(new_n373_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n360_), .A2(new_n361_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n379_), .A2(new_n341_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT72), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n379_), .A2(KEYINPUT72), .A3(new_n341_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n383_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(new_n362_), .A4(new_n373_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT73), .B(G190gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G218gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(G134gat), .B(G162gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n396_));
  NAND4_X1  g195(.A1(new_n384_), .A2(new_n391_), .A3(new_n395_), .A4(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n357_), .B1(new_n397_), .B2(KEYINPUT75), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n395_), .B(KEYINPUT36), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n372_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n390_), .B1(new_n400_), .B2(new_n362_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n382_), .A2(new_n383_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n399_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n397_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n398_), .A2(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n403_), .B(new_n397_), .C1(KEYINPUT75), .C2(new_n357_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT16), .B(G183gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(G211gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G127gat), .B(G155gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n411_), .A2(KEYINPUT17), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT78), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(KEYINPUT17), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n413_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(G231gat), .A2(G233gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n339_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G1gat), .B(G8gat), .Z(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G1gat), .A2(G8gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT14), .ZN(new_n424_));
  INV_X1    g223(.A(G15gat), .ZN(new_n425_));
  INV_X1    g224(.A(G22gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(G15gat), .A2(G22gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n424_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT76), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n429_), .A2(KEYINPUT76), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n422_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n432_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(new_n421_), .A3(new_n430_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n339_), .A2(new_n418_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n420_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n437_), .B1(new_n420_), .B2(new_n438_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n417_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT79), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT79), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n417_), .B(new_n443_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  OR3_X1    g244(.A1(new_n439_), .A2(new_n440_), .A3(KEYINPUT68), .ZN(new_n446_));
  INV_X1    g245(.A(new_n414_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT68), .B1(new_n439_), .B2(new_n440_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT77), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT77), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n446_), .A2(new_n451_), .A3(new_n447_), .A4(new_n448_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n445_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT80), .B1(new_n407_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT80), .ZN(new_n456_));
  AOI211_X1 g255(.A(new_n456_), .B(new_n453_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n457_));
  OAI211_X1 g256(.A(KEYINPUT81), .B(new_n356_), .C1(new_n455_), .C2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G183gat), .A2(G190gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT23), .ZN(new_n460_));
  OR2_X1    g259(.A1(G169gat), .A2(G176gat), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n461_), .A2(KEYINPUT24), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G169gat), .A2(G176gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n461_), .A2(KEYINPUT24), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT84), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT25), .B(G183gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT26), .B(G190gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n465_), .A2(new_n466_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n463_), .A2(new_n467_), .A3(new_n470_), .A4(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n460_), .B1(G183gat), .B2(G190gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT22), .B(G169gat), .Z(new_n474_));
  OAI211_X1 g273(.A(new_n473_), .B(new_n464_), .C1(G176gat), .C2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT85), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT30), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n472_), .A2(new_n475_), .A3(KEYINPUT85), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n479_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT30), .B1(new_n481_), .B2(new_n476_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n207_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n482_), .A3(new_n207_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G15gat), .B(G43gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT86), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT31), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n485_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n488_), .B1(new_n491_), .B2(new_n483_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G71gat), .B(G99gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G227gat), .A2(G233gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  AND3_X1   g294(.A1(new_n490_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n495_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G78gat), .B(G106gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(new_n367_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT88), .B(G204gat), .ZN(new_n501_));
  INV_X1    g300(.A(G197gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n503_), .B(KEYINPUT21), .C1(new_n502_), .C2(new_n349_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G211gat), .B(G218gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(G197gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n506_), .B1(G197gat), .B2(new_n349_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n504_), .B(new_n505_), .C1(new_n507_), .C2(KEYINPUT21), .ZN(new_n508_));
  INV_X1    g307(.A(new_n505_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(KEYINPUT21), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n228_), .A2(KEYINPUT29), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G228gat), .A2(G233gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n514_), .A2(KEYINPUT89), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(KEYINPUT89), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n513_), .A2(new_n516_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n500_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n500_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n518_), .B(new_n522_), .C1(new_n513_), .C2(new_n516_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  OR3_X1    g323(.A1(new_n228_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT28), .B1(new_n228_), .B2(KEYINPUT29), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT90), .B(G22gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n525_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n528_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n524_), .B(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n463_), .A2(new_n470_), .A3(new_n465_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT91), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n475_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n511_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n511_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n477_), .A2(new_n538_), .A3(new_n479_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(KEYINPUT20), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G226gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT19), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n511_), .B1(new_n481_), .B2(new_n476_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n544_), .A2(KEYINPUT20), .ZN(new_n545_));
  INV_X1    g344(.A(new_n542_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n535_), .A2(new_n475_), .A3(new_n538_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n545_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n543_), .A2(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(G8gat), .B(G36gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(G64gat), .B(G92gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n552_), .B(new_n553_), .Z(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT33), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT94), .B1(new_n246_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n554_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n543_), .A2(new_n548_), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n246_), .A2(new_n556_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n555_), .A2(new_n557_), .A3(new_n559_), .A4(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n230_), .B1(KEYINPUT4), .B2(new_n229_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(new_n232_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n234_), .B(KEYINPUT95), .ZN(new_n564_));
  AOI211_X1 g363(.A(new_n245_), .B(new_n563_), .C1(new_n232_), .C2(new_n564_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n246_), .A2(KEYINPUT94), .A3(new_n556_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n561_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n540_), .A2(new_n542_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n538_), .A2(new_n475_), .A3(new_n533_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n546_), .B1(new_n545_), .B2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(KEYINPUT32), .B(new_n558_), .C1(new_n568_), .C2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n558_), .A2(KEYINPUT32), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n543_), .A2(new_n548_), .A3(new_n572_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n247_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n498_), .B(new_n532_), .C1(new_n567_), .C2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT27), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n543_), .A2(new_n558_), .A3(new_n548_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n558_), .B1(new_n543_), .B2(new_n548_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n576_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  OAI211_X1 g380(.A(KEYINPUT96), .B(new_n576_), .C1(new_n577_), .C2(new_n578_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n532_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n490_), .A2(new_n492_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n495_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n524_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n521_), .A2(new_n531_), .A3(new_n523_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n490_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n587_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n584_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n247_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n554_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(KEYINPUT27), .A3(new_n559_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n583_), .A2(new_n593_), .A3(new_n594_), .A4(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n575_), .A2(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n458_), .A2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n356_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT81), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n371_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n436_), .A2(new_n374_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G229gat), .A2(G233gat), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n377_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n605_), .B2(new_n375_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n609_), .B1(new_n611_), .B2(new_n608_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G169gat), .B(G197gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(G141gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT82), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(G113gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n612_), .B(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT83), .Z(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n599_), .A2(KEYINPUT97), .A3(new_n602_), .A4(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n458_), .A2(new_n598_), .A3(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n407_), .A2(new_n454_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n456_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n453_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT80), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT81), .B1(new_n628_), .B2(new_n356_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n622_), .B1(new_n623_), .B2(new_n629_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n620_), .A2(new_n621_), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n621_), .B1(new_n620_), .B2(new_n630_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n202_), .B(new_n247_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n404_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(new_n453_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n575_), .B2(new_n597_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n356_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n617_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n594_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n633_), .A2(new_n634_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n635_), .A2(new_n645_), .A3(new_n646_), .ZN(G1324gat));
  INV_X1    g446(.A(G8gat), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n583_), .A2(new_n596_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n648_), .B(new_n649_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n598_), .A2(new_n642_), .A3(new_n649_), .A4(new_n637_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT99), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n639_), .A2(new_n655_), .A3(new_n642_), .A4(new_n649_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n653_), .A2(new_n654_), .A3(G8gat), .A4(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT39), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n653_), .A2(G8gat), .A3(new_n656_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT100), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n658_), .B(new_n660_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n650_), .A2(new_n651_), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n651_), .B1(new_n650_), .B2(new_n661_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  INV_X1    g463(.A(new_n498_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n425_), .B1(new_n643_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT41), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n620_), .A2(new_n630_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(new_n425_), .A3(new_n665_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n669_), .A2(new_n670_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n667_), .B1(new_n671_), .B2(new_n672_), .ZN(G1326gat));
  AOI21_X1  g472(.A(new_n426_), .B1(new_n643_), .B2(new_n590_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT103), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT42), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n668_), .A2(new_n426_), .A3(new_n590_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1327gat));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  INV_X1    g478(.A(new_n407_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n598_), .B2(new_n680_), .ZN(new_n681_));
  AOI211_X1 g480(.A(KEYINPUT43), .B(new_n407_), .C1(new_n575_), .C2(new_n597_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n640_), .A2(new_n454_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n683_), .A2(KEYINPUT44), .A3(new_n617_), .A4(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n617_), .B(new_n684_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G29gat), .B1(new_n689_), .B2(new_n594_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n404_), .B1(new_n575_), .B2(new_n597_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n691_), .A2(new_n619_), .A3(new_n684_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n594_), .A2(G29gat), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT104), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n690_), .A2(new_n695_), .ZN(G1328gat));
  INV_X1    g495(.A(new_n649_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G36gat), .B1(new_n689_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(G36gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n692_), .A2(new_n699_), .A3(new_n649_), .ZN(new_n700_));
  XOR2_X1   g499(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n698_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n698_), .A2(KEYINPUT46), .A3(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n665_), .A2(G43gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n689_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n709_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n685_), .A2(KEYINPUT106), .A3(new_n688_), .A4(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n692_), .A2(new_n665_), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT107), .B(G43gat), .Z(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n710_), .A2(new_n712_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT47), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n710_), .A2(new_n718_), .A3(new_n712_), .A4(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1330gat));
  NOR3_X1   g519(.A1(new_n689_), .A2(new_n367_), .A3(new_n532_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G50gat), .B1(new_n692_), .B2(new_n590_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1331gat));
  AND3_X1   g522(.A1(new_n639_), .A2(new_n640_), .A3(new_n618_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(G57gat), .A3(new_n247_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT109), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n628_), .A2(new_n641_), .A3(new_n640_), .A4(new_n598_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n594_), .B1(new_n728_), .B2(KEYINPUT108), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n729_), .B1(KEYINPUT108), .B2(new_n728_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n726_), .B1(new_n294_), .B2(new_n730_), .ZN(G1332gat));
  AOI21_X1  g530(.A(new_n295_), .B1(new_n724_), .B2(new_n649_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT48), .Z(new_n733_));
  NAND3_X1  g532(.A1(new_n728_), .A2(new_n295_), .A3(new_n649_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1333gat));
  AOI21_X1  g534(.A(new_n301_), .B1(new_n724_), .B2(new_n665_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT49), .Z(new_n737_));
  NAND3_X1  g536(.A1(new_n728_), .A2(new_n301_), .A3(new_n665_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(G1334gat));
  AOI21_X1  g540(.A(new_n303_), .B1(new_n724_), .B2(new_n590_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT50), .Z(new_n743_));
  NAND3_X1  g542(.A1(new_n728_), .A2(new_n303_), .A3(new_n590_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1335gat));
  NOR3_X1   g544(.A1(new_n356_), .A2(new_n617_), .A3(new_n454_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n691_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G85gat), .B1(new_n748_), .B2(new_n247_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n683_), .A2(new_n746_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n594_), .B1(new_n282_), .B2(new_n286_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(G1336gat));
  NAND3_X1  g551(.A1(new_n750_), .A2(G92gat), .A3(new_n649_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n250_), .B1(new_n747_), .B2(new_n697_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT111), .Z(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT112), .Z(G1337gat));
  NAND2_X1  g556(.A1(new_n750_), .A2(new_n665_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G99gat), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n760_), .A2(KEYINPUT113), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n748_), .A2(new_n278_), .A3(new_n665_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n760_), .A2(KEYINPUT113), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT114), .Z(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n763_), .B(new_n766_), .ZN(G1338gat));
  OAI211_X1 g566(.A(new_n590_), .B(new_n746_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(G106gat), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n691_), .A2(new_n746_), .A3(new_n255_), .A4(new_n590_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT115), .Z(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n772_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT116), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n771_), .A2(new_n774_), .A3(new_n777_), .A4(new_n772_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n776_), .A2(KEYINPUT53), .A3(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1339gat));
  NAND2_X1  g582(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n626_), .A2(new_n356_), .A3(new_n618_), .A4(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n785_), .B(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n612_), .A2(new_n616_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n616_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n606_), .A2(new_n608_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n789_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(new_n355_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT120), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n324_), .A2(new_n796_), .A3(KEYINPUT55), .A4(new_n344_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n322_), .A2(new_n323_), .B1(new_n338_), .B2(new_n343_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n796_), .B1(new_n799_), .B2(KEYINPUT55), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n344_), .A2(new_n318_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n319_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n345_), .A2(new_n802_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n353_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n795_), .B1(new_n806_), .B2(KEYINPUT56), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n324_), .A2(KEYINPUT55), .A3(new_n344_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT119), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n345_), .A2(new_n802_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n803_), .A2(new_n804_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .A4(new_n797_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n354_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT121), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n812_), .B2(new_n354_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT120), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n812_), .A2(KEYINPUT121), .A3(KEYINPUT56), .A4(new_n354_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n807_), .A2(new_n815_), .A3(new_n817_), .A4(new_n818_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n347_), .A2(new_n354_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n617_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n617_), .A2(new_n820_), .A3(KEYINPUT118), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n794_), .B1(new_n819_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n788_), .B1(new_n826_), .B2(new_n636_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n823_), .A2(new_n824_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n815_), .A2(new_n818_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n812_), .A2(new_n354_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT120), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  AOI211_X1 g631(.A(new_n795_), .B(KEYINPUT56), .C1(new_n812_), .C2(new_n354_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n828_), .B1(new_n829_), .B2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT57), .B(new_n404_), .C1(new_n835_), .C2(new_n794_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n813_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n793_), .B(new_n820_), .C1(new_n837_), .C2(new_n816_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n407_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n820_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n816_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n813_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n845_), .A2(KEYINPUT122), .A3(KEYINPUT58), .A4(new_n793_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n840_), .A2(new_n842_), .A3(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n827_), .A2(new_n836_), .A3(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n787_), .B1(new_n848_), .B2(new_n453_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n649_), .A2(new_n594_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n584_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n849_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(G113gat), .B1(new_n853_), .B2(new_n617_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n848_), .A2(new_n453_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n787_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n852_), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT59), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n849_), .A2(new_n861_), .A3(new_n852_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n204_), .B1(new_n860_), .B2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n854_), .B1(new_n864_), .B2(new_n619_), .ZN(G1340gat));
  OAI21_X1  g664(.A(new_n640_), .B1(new_n859_), .B2(new_n862_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT123), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n868_), .B(new_n640_), .C1(new_n859_), .C2(new_n862_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n867_), .A2(G120gat), .A3(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n206_), .B1(new_n356_), .B2(KEYINPUT60), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n853_), .B(new_n871_), .C1(KEYINPUT60), .C2(new_n206_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(G1341gat));
  AOI21_X1  g672(.A(G127gat), .B1(new_n853_), .B2(new_n454_), .ZN(new_n874_));
  INV_X1    g673(.A(G127gat), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n454_), .B2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n860_), .B2(new_n863_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n875_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n874_), .B1(new_n878_), .B2(new_n879_), .ZN(G1342gat));
  AOI21_X1  g679(.A(G134gat), .B1(new_n853_), .B2(new_n636_), .ZN(new_n881_));
  INV_X1    g680(.A(G134gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n860_), .B2(new_n863_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n883_), .B2(new_n680_), .ZN(G1343gat));
  NOR2_X1   g683(.A1(new_n849_), .A2(new_n592_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n850_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n641_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n208_), .ZN(G1344gat));
  NOR2_X1   g687(.A1(new_n886_), .A2(new_n356_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(new_n209_), .ZN(G1345gat));
  NOR2_X1   g689(.A1(new_n886_), .A2(new_n453_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT61), .B(G155gat), .Z(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT125), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n891_), .B(new_n893_), .ZN(G1346gat));
  INV_X1    g693(.A(G162gat), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n886_), .A2(new_n895_), .A3(new_n407_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n885_), .A2(new_n636_), .A3(new_n850_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n895_), .B2(new_n897_), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n697_), .A2(new_n247_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n849_), .A2(new_n584_), .A3(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n617_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G169gat), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n902_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n905_), .B(new_n906_), .C1(new_n474_), .C2(new_n902_), .ZN(G1348gat));
  NAND2_X1  g706(.A1(new_n901_), .A2(new_n640_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g708(.A1(new_n901_), .A2(new_n454_), .ZN(new_n910_));
  MUX2_X1   g709(.A(new_n468_), .B(G183gat), .S(new_n910_), .Z(G1350gat));
  INV_X1    g710(.A(new_n901_), .ZN(new_n912_));
  OAI21_X1  g711(.A(G190gat), .B1(new_n912_), .B2(new_n407_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n901_), .A2(new_n469_), .A3(new_n636_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1351gat));
  NAND2_X1  g714(.A1(new_n885_), .A2(new_n899_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n641_), .ZN(new_n917_));
  XOR2_X1   g716(.A(KEYINPUT126), .B(G197gat), .Z(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1352gat));
  NOR2_X1   g718(.A1(new_n916_), .A2(new_n356_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n501_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n921_), .B1(new_n920_), .B2(new_n349_), .ZN(G1353gat));
  NOR4_X1   g721(.A1(new_n849_), .A2(new_n592_), .A3(new_n453_), .A4(new_n900_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT63), .B(G211gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n923_), .B2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT127), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n925_), .B(new_n929_), .C1(new_n923_), .C2(new_n926_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1354gat));
  INV_X1    g730(.A(G218gat), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n916_), .A2(new_n932_), .A3(new_n407_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n885_), .A2(new_n636_), .A3(new_n899_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n932_), .B2(new_n934_), .ZN(G1355gat));
endmodule


