//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n203_), .B(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT10), .B(G99gat), .Z(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT64), .ZN(new_n211_));
  NAND2_X1  g010(.A1(KEYINPUT9), .A2(G85gat), .ZN(new_n212_));
  INV_X1    g011(.A(G92gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(KEYINPUT9), .B2(G85gat), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n206_), .B(new_n209_), .C1(new_n211_), .C2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  INV_X1    g016(.A(G99gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n218_), .B(new_n208_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n219_), .A2(new_n220_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n223_));
  OAI22_X1  g022(.A1(new_n222_), .A2(new_n223_), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n206_), .A2(new_n221_), .A3(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G85gat), .B(G92gat), .Z(new_n226_));
  AOI21_X1  g025(.A(new_n217_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n203_), .B(new_n204_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n221_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n226_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(KEYINPUT8), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n216_), .B1(new_n227_), .B2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n235_));
  XOR2_X1   g034(.A(G71gat), .B(G78gat), .Z(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n235_), .A2(new_n236_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(new_n240_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n216_), .B(new_n239_), .C1(new_n227_), .C2(new_n231_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(KEYINPUT12), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT12), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n232_), .A2(new_n244_), .A3(new_n240_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G230gat), .A2(G233gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n241_), .A2(new_n242_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n247_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(KEYINPUT67), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n250_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n248_), .A2(new_n251_), .A3(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G120gat), .B(G148gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT5), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G176gat), .B(G204gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  AND2_X1   g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n255_), .A2(new_n259_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n202_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n260_), .A2(new_n261_), .A3(new_n202_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n263_), .A2(new_n264_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT68), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G127gat), .B(G155gat), .Z(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT16), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G183gat), .B(G211gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT17), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT76), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G15gat), .B(G22gat), .ZN(new_n279_));
  INV_X1    g078(.A(G1gat), .ZN(new_n280_));
  INV_X1    g079(.A(G8gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT14), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G1gat), .B(G8gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G231gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(new_n239_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n278_), .A2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n289_), .A2(KEYINPUT77), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n288_), .A2(new_n276_), .A3(new_n275_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT75), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(KEYINPUT77), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n290_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT78), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n290_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT78), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n232_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G29gat), .B(G36gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G43gat), .B(G50gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(new_n306_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n301_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n309_), .B(KEYINPUT15), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n311_), .B1(new_n301_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G232gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT34), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n315_), .B(KEYINPUT35), .Z(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(KEYINPUT35), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n313_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n313_), .A2(KEYINPUT73), .A3(new_n316_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(G190gat), .B(G218gat), .Z(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT71), .ZN(new_n325_));
  XOR2_X1   g124(.A(G134gat), .B(G162gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT36), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n330_));
  AND2_X1   g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n319_), .A2(new_n321_), .A3(new_n322_), .A4(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT37), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n334_), .B1(new_n332_), .B2(KEYINPUT74), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n329_), .B(new_n332_), .C1(KEYINPUT74), .C2(new_n334_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n300_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n271_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G1gat), .B(G29gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G57gat), .B(G85gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G134gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G127gat), .ZN(new_n348_));
  INV_X1    g147(.A(G127gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G134gat), .ZN(new_n350_));
  INV_X1    g149(.A(G120gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G113gat), .ZN(new_n352_));
  INV_X1    g151(.A(G113gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(G120gat), .ZN(new_n354_));
  AND4_X1   g153(.A1(new_n348_), .A2(new_n350_), .A3(new_n352_), .A4(new_n354_), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n348_), .A2(new_n350_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT86), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n360_), .A2(new_n361_), .A3(KEYINPUT1), .ZN(new_n362_));
  INV_X1    g161(.A(G141gat), .ZN(new_n363_));
  INV_X1    g162(.A(G148gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G141gat), .A2(G148gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n365_), .B(new_n366_), .C1(new_n367_), .C2(new_n359_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n358_), .B1(new_n362_), .B2(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n365_), .A2(new_n366_), .ZN(new_n370_));
  OR2_X1    g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(new_n367_), .A3(new_n359_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n360_), .A2(KEYINPUT1), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n370_), .A2(new_n372_), .A3(KEYINPUT86), .A4(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n360_), .A2(new_n361_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT87), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT87), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n379_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n366_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n363_), .A2(new_n364_), .A3(KEYINPUT3), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(G141gat), .B2(G148gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n381_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n376_), .B1(new_n388_), .B2(KEYINPUT88), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n384_), .A2(new_n386_), .B1(new_n382_), .B2(new_n366_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT88), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n381_), .ZN(new_n392_));
  AOI221_X4 g191(.A(new_n357_), .B1(new_n369_), .B2(new_n374_), .C1(new_n389_), .C2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n357_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n388_), .A2(KEYINPUT88), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(new_n375_), .A3(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n369_), .A2(new_n374_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n394_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT98), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n401_), .B(KEYINPUT96), .Z(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n399_), .A2(new_n400_), .A3(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n390_), .A2(new_n391_), .A3(new_n381_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n391_), .B1(new_n390_), .B2(new_n381_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n376_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n397_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n357_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n396_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n403_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT98), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n404_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n403_), .B1(new_n398_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n409_), .A2(KEYINPUT4), .A3(new_n410_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT95), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n409_), .A2(KEYINPUT95), .A3(KEYINPUT4), .A4(new_n410_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n416_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n346_), .B1(new_n413_), .B2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT95), .B1(new_n399_), .B2(KEYINPUT4), .ZN(new_n423_));
  INV_X1    g222(.A(new_n420_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n415_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n404_), .A2(new_n412_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n345_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G78gat), .B(G106gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n429_), .B(KEYINPUT90), .Z(new_n430_));
  NAND2_X1  g229(.A1(G228gat), .A2(G233gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT29), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G211gat), .B(G218gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(G197gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(G204gat), .ZN(new_n438_));
  INV_X1    g237(.A(G204gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(G197gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n436_), .B1(KEYINPUT21), .B2(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n438_), .A2(KEYINPUT89), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n438_), .A2(KEYINPUT89), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT21), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .A4(new_n440_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n444_), .A3(new_n440_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n435_), .A2(new_n445_), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n442_), .A2(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n432_), .B1(new_n434_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n449_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n389_), .A2(new_n392_), .B1(new_n369_), .B2(new_n374_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n431_), .B(new_n451_), .C1(new_n452_), .C2(new_n433_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n430_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(new_n430_), .A3(new_n453_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n452_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT28), .B1(new_n457_), .B2(KEYINPUT29), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT28), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n452_), .A2(new_n459_), .A3(new_n433_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G22gat), .B(G50gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n458_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n455_), .A2(new_n456_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT91), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT92), .ZN(new_n468_));
  OAI22_X1  g267(.A1(new_n454_), .A2(new_n467_), .B1(new_n456_), .B2(new_n468_), .ZN(new_n469_));
  AOI211_X1 g268(.A(KEYINPUT91), .B(new_n430_), .C1(new_n450_), .C2(new_n453_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n456_), .A2(new_n468_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n472_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n466_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G8gat), .B(G36gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT18), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G64gat), .B(G92gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  NOR2_X1   g278(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(G169gat), .ZN(new_n481_));
  INV_X1    g280(.A(G183gat), .ZN(new_n482_));
  INV_X1    g281(.A(G190gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT23), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT23), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(G183gat), .A3(G190gat), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(G183gat), .A2(G190gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n481_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(KEYINPUT83), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT83), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n491_), .A2(new_n485_), .A3(G183gat), .A4(G190gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n484_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G169gat), .A2(G176gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT81), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT24), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  OR3_X1    g300(.A1(new_n483_), .A2(KEYINPUT80), .A3(KEYINPUT26), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT25), .B(G183gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT26), .B1(new_n483_), .B2(KEYINPUT80), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n494_), .A2(new_n501_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n500_), .B1(G169gat), .B2(G176gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT82), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT82), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n507_), .A2(new_n497_), .A3(new_n510_), .A4(new_n498_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n489_), .B1(new_n506_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT84), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n515_), .B(new_n489_), .C1(new_n506_), .C2(new_n512_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n449_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT94), .ZN(new_n518_));
  INV_X1    g317(.A(new_n488_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n494_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n485_), .B1(G183gat), .B2(G190gat), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT94), .B1(new_n522_), .B2(new_n488_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n481_), .A3(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT26), .B(G190gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n503_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n508_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT93), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n487_), .B1(new_n500_), .B2(new_n495_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n526_), .A2(new_n508_), .A3(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n528_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n524_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n451_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n517_), .A2(KEYINPUT20), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G226gat), .A2(G233gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT19), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n524_), .A2(new_n449_), .A3(new_n532_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT20), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT100), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n514_), .A2(new_n516_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n451_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n540_), .A2(KEYINPUT100), .A3(KEYINPUT20), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n543_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n537_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n479_), .B1(new_n539_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n535_), .A2(new_n537_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n537_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n541_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n545_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n550_), .A2(new_n553_), .A3(new_n479_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT27), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n549_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n550_), .A2(new_n553_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n479_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n554_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT101), .B(KEYINPUT27), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT102), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n550_), .A2(new_n479_), .A3(new_n553_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n479_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n565_));
  OAI211_X1 g364(.A(KEYINPUT102), .B(new_n562_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n557_), .B1(new_n563_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT103), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n562_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT102), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n566_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT103), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n574_), .A3(new_n557_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n475_), .B1(new_n569_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G71gat), .B(G99gat), .ZN(new_n577_));
  INV_X1    g376(.A(G43gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n544_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n544_), .A2(new_n579_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G227gat), .A2(G233gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(G15gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT30), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n580_), .A2(new_n585_), .A3(new_n581_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT85), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT85), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n587_), .A2(new_n591_), .A3(new_n588_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n357_), .B(KEYINPUT31), .Z(new_n593_));
  NAND3_X1  g392(.A1(new_n590_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n593_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(KEYINPUT85), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n597_), .A2(new_n428_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n402_), .B1(new_n398_), .B2(new_n414_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n599_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n345_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n345_), .A2(KEYINPUT33), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n404_), .B2(new_n412_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n425_), .A2(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n560_), .A2(new_n602_), .A3(new_n605_), .A4(new_n554_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n413_), .A2(new_n421_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT33), .B1(new_n607_), .B2(new_n345_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT99), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n564_), .A2(new_n565_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n427_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n600_), .A2(new_n601_), .B1(new_n425_), .B2(new_n604_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n610_), .A2(new_n612_), .A3(new_n613_), .A4(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n558_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n479_), .A2(KEYINPUT32), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n422_), .A2(new_n427_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n539_), .A2(new_n548_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(KEYINPUT32), .A3(new_n479_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n609_), .A2(new_n615_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n474_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n474_), .A2(new_n428_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n624_), .B(new_n557_), .C1(new_n563_), .C2(new_n567_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  AOI22_X1  g425(.A1(new_n576_), .A2(new_n598_), .B1(new_n626_), .B2(new_n597_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n312_), .A2(new_n285_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n310_), .A2(new_n285_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G229gat), .A2(G233gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n309_), .B(new_n285_), .Z(new_n632_));
  INV_X1    g431(.A(new_n630_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G113gat), .B(G141gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT79), .ZN(new_n637_));
  XOR2_X1   g436(.A(G169gat), .B(G197gat), .Z(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n635_), .B(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n627_), .A2(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n340_), .A2(new_n280_), .A3(new_n428_), .A4(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT38), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n643_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n333_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n627_), .A2(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n265_), .A2(new_n296_), .A3(new_n640_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(new_n428_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G1gat), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n651_), .A2(KEYINPUT104), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(KEYINPUT104), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n644_), .B(new_n645_), .C1(new_n652_), .C2(new_n653_), .ZN(G1324gat));
  AOI21_X1  g453(.A(new_n574_), .B1(new_n573_), .B2(new_n557_), .ZN(new_n655_));
  AOI211_X1 g454(.A(KEYINPUT103), .B(new_n556_), .C1(new_n572_), .C2(new_n566_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n647_), .A2(new_n657_), .A3(new_n648_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(KEYINPUT105), .A2(KEYINPUT39), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n281_), .B1(KEYINPUT105), .B2(KEYINPUT39), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n658_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n659_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n340_), .A2(new_n281_), .A3(new_n657_), .A4(new_n641_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(G1325gat));
  INV_X1    g466(.A(new_n597_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n649_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G15gat), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT107), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(new_n672_), .A3(G15gat), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(KEYINPUT41), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(KEYINPUT41), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n340_), .A2(new_n641_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n677_), .A2(G15gat), .A3(new_n597_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT108), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n676_), .A3(new_n679_), .ZN(G1326gat));
  OR3_X1    g479(.A1(new_n677_), .A2(G22gat), .A3(new_n474_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n649_), .A2(new_n475_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G22gat), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT42), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(KEYINPUT42), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(G1327gat));
  NAND2_X1  g485(.A1(new_n299_), .A2(new_n646_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(new_n265_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n641_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G29gat), .B1(new_n690_), .B2(new_n428_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT110), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n692_), .B(new_n694_), .C1(new_n627_), .C2(new_n338_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n610_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n696_));
  AOI22_X1  g495(.A1(new_n696_), .A2(KEYINPUT99), .B1(new_n620_), .B2(new_n618_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n475_), .B1(new_n697_), .B2(new_n615_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n625_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n597_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n474_), .B(new_n598_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n338_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT110), .B1(new_n702_), .B2(new_n693_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n695_), .A2(new_n703_), .A3(new_n705_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n300_), .A2(new_n265_), .A3(new_n640_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n706_), .A2(KEYINPUT44), .A3(new_n707_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n428_), .A2(G29gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n691_), .B1(new_n711_), .B2(new_n712_), .ZN(G1328gat));
  INV_X1    g512(.A(new_n657_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n689_), .A2(G36gat), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n708_), .A2(new_n710_), .A3(new_n714_), .ZN(new_n718_));
  INV_X1    g517(.A(G36gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n717_), .B(KEYINPUT46), .C1(new_n718_), .C2(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1329gat));
  NAND3_X1  g523(.A1(new_n706_), .A2(KEYINPUT44), .A3(new_n707_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n597_), .A2(new_n578_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n706_), .A2(new_n707_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n725_), .B(new_n726_), .C1(new_n727_), .C2(new_n709_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n578_), .B1(new_n689_), .B2(new_n597_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(G1330gat));
  AOI21_X1  g531(.A(G50gat), .B1(new_n690_), .B2(new_n475_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n475_), .A2(G50gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n711_), .B2(new_n734_), .ZN(G1331gat));
  INV_X1    g534(.A(new_n640_), .ZN(new_n736_));
  NOR4_X1   g535(.A1(new_n627_), .A2(new_n339_), .A3(new_n736_), .A4(new_n268_), .ZN(new_n737_));
  INV_X1    g536(.A(G57gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n428_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n299_), .A2(new_n736_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n647_), .A2(new_n271_), .A3(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(new_n428_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n739_), .B1(new_n742_), .B2(new_n738_), .ZN(G1332gat));
  INV_X1    g542(.A(G64gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n737_), .A2(new_n744_), .A3(new_n657_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n741_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G64gat), .B1(new_n746_), .B2(new_n714_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(KEYINPUT48), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(KEYINPUT48), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1333gat));
  INV_X1    g549(.A(G71gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n737_), .A2(new_n751_), .A3(new_n668_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G71gat), .B1(new_n746_), .B2(new_n597_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(KEYINPUT49), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(KEYINPUT49), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n752_), .B1(new_n754_), .B2(new_n755_), .ZN(G1334gat));
  NOR2_X1   g555(.A1(new_n474_), .A2(G78gat), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT113), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n737_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G78gat), .B1(new_n746_), .B2(new_n474_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(KEYINPUT50), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(KEYINPUT50), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n761_), .B2(new_n762_), .ZN(G1335gat));
  NOR4_X1   g562(.A1(new_n270_), .A2(new_n627_), .A3(new_n736_), .A4(new_n687_), .ZN(new_n764_));
  AOI21_X1  g563(.A(G85gat), .B1(new_n764_), .B2(new_n428_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n300_), .A2(new_n736_), .A3(new_n268_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n706_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n428_), .A2(G85gat), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT114), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n765_), .B1(new_n767_), .B2(new_n769_), .ZN(G1336gat));
  NAND3_X1  g569(.A1(new_n764_), .A2(new_n213_), .A3(new_n657_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n767_), .A2(new_n657_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(new_n213_), .ZN(G1337gat));
  NAND3_X1  g572(.A1(new_n706_), .A2(new_n668_), .A3(new_n766_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(G99gat), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n764_), .A2(new_n668_), .A3(new_n207_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g577(.A1(new_n764_), .A2(new_n208_), .A3(new_n475_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT115), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n706_), .A2(new_n475_), .A3(new_n766_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(G106gat), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n780_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT53), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n780_), .A2(new_n784_), .A3(new_n788_), .A4(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1339gat));
  NAND3_X1  g589(.A1(new_n740_), .A2(new_n268_), .A3(new_n338_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n248_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n250_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT116), .B1(new_n797_), .B2(KEYINPUT55), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n243_), .A2(new_n250_), .A3(new_n245_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(KEYINPUT55), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n796_), .A2(new_n798_), .A3(new_n799_), .A4(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(KEYINPUT56), .A3(new_n259_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n801_), .A2(KEYINPUT117), .A3(KEYINPUT56), .A4(new_n259_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n801_), .A2(new_n259_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT56), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n804_), .A2(new_n805_), .A3(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n631_), .A2(new_n634_), .A3(new_n639_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n628_), .A2(new_n629_), .A3(new_n633_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n639_), .B1(new_n632_), .B2(new_n630_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n261_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n809_), .A2(KEYINPUT58), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT58), .B1(new_n809_), .B2(new_n815_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n338_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n640_), .A2(new_n261_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n808_), .B2(new_n802_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n260_), .A2(new_n261_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n822_), .A2(new_n814_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n333_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(KEYINPUT57), .B(new_n333_), .C1(new_n821_), .C2(new_n823_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n299_), .B1(new_n819_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n793_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT119), .B(new_n299_), .C1(new_n819_), .C2(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n576_), .A2(new_n428_), .A3(new_n668_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n826_), .A2(new_n827_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n818_), .A2(new_n338_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n816_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n294_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n793_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT59), .B1(new_n842_), .B2(new_n835_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n837_), .A2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n640_), .A2(new_n353_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT120), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n736_), .B(new_n836_), .C1(new_n841_), .C2(new_n793_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(KEYINPUT118), .A3(new_n353_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n353_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n844_), .A2(new_n846_), .B1(new_n848_), .B2(new_n851_), .ZN(G1340gat));
  NAND3_X1  g651(.A1(new_n837_), .A2(new_n271_), .A3(new_n843_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(G120gat), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n842_), .A2(new_n835_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n351_), .B1(new_n268_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n855_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n351_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(new_n857_), .ZN(G1341gat));
  NAND3_X1  g657(.A1(new_n837_), .A2(new_n294_), .A3(new_n843_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(G127gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n855_), .A2(new_n349_), .A3(new_n300_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1342gat));
  INV_X1    g661(.A(new_n338_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n837_), .A2(new_n863_), .A3(new_n843_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G134gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n855_), .A2(new_n347_), .A3(new_n646_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1343gat));
  NAND4_X1  g666(.A1(new_n714_), .A2(new_n428_), .A3(new_n475_), .A4(new_n597_), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(KEYINPUT121), .Z(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n841_), .B2(new_n793_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n640_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n363_), .ZN(G1344gat));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n270_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT122), .B(G148gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1345gat));
  NOR2_X1   g674(.A1(new_n870_), .A2(new_n299_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT61), .B(G155gat), .Z(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1346gat));
  OAI21_X1  g677(.A(G162gat), .B1(new_n870_), .B2(new_n338_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n333_), .A2(G162gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n870_), .B2(new_n880_), .ZN(G1347gat));
  AND2_X1   g680(.A1(new_n657_), .A2(new_n598_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n475_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n887_));
  AND2_X1   g686(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n886_), .B(new_n736_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(G169gat), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n882_), .A2(new_n736_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT123), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n475_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n890_), .B1(new_n833_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n895_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n889_), .B1(new_n896_), .B2(new_n897_), .ZN(G1348gat));
  NAND3_X1  g697(.A1(new_n833_), .A2(new_n265_), .A3(new_n884_), .ZN(new_n899_));
  INV_X1    g698(.A(G176gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n271_), .A2(G176gat), .A3(new_n882_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n842_), .A2(new_n475_), .A3(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n901_), .A2(new_n902_), .A3(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G176gat), .B1(new_n886_), .B2(new_n265_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT124), .B1(new_n907_), .B2(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1349gat));
  INV_X1    g708(.A(new_n842_), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n910_), .A2(new_n474_), .A3(new_n300_), .A4(new_n882_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n296_), .A2(new_n503_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n911_), .A2(new_n482_), .B1(new_n886_), .B2(new_n912_), .ZN(G1350gat));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n483_), .B1(new_n886_), .B2(new_n863_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n646_), .A2(new_n525_), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n833_), .A2(new_n884_), .A3(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n914_), .B1(new_n915_), .B2(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n833_), .A2(new_n863_), .A3(new_n884_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(G190gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n886_), .A2(new_n916_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n920_), .A2(KEYINPUT125), .A3(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n918_), .A2(new_n922_), .ZN(G1351gat));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n657_), .A2(new_n624_), .A3(new_n597_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n842_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n925_), .ZN(new_n927_));
  OAI211_X1 g726(.A(KEYINPUT126), .B(new_n927_), .C1(new_n841_), .C2(new_n793_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n640_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(new_n437_), .ZN(G1352gat));
  AOI21_X1  g729(.A(new_n270_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(new_n439_), .ZN(G1353gat));
  XNOR2_X1  g731(.A(KEYINPUT63), .B(G211gat), .ZN(new_n933_));
  AOI211_X1 g732(.A(new_n296_), .B(new_n933_), .C1(new_n926_), .C2(new_n928_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n926_), .A2(new_n928_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n294_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n934_), .B1(new_n936_), .B2(new_n937_), .ZN(G1354gat));
  NAND2_X1  g737(.A1(new_n935_), .A2(new_n646_), .ZN(new_n939_));
  INV_X1    g738(.A(G218gat), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n863_), .A2(G218gat), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(KEYINPUT127), .ZN(new_n942_));
  AOI22_X1  g741(.A1(new_n939_), .A2(new_n940_), .B1(new_n935_), .B2(new_n942_), .ZN(G1355gat));
endmodule


