//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT20), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G197gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT85), .B1(new_n214_), .B2(G204gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT85), .ZN(new_n216_));
  INV_X1    g015(.A(G204gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(G197gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(G204gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n213_), .B1(new_n220_), .B2(KEYINPUT21), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT86), .B1(new_n217_), .B2(G197gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT86), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(new_n214_), .A3(G204gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT21), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n214_), .A2(G204gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AND4_X1   g027(.A1(KEYINPUT87), .A2(new_n225_), .A3(new_n226_), .A4(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n227_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT87), .B1(new_n230_), .B2(new_n226_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n221_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n230_), .A2(new_n226_), .A3(new_n212_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G169gat), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n241_));
  INV_X1    g040(.A(G183gat), .ZN(new_n242_));
  INV_X1    g041(.A(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G169gat), .A2(G176gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n238_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n243_), .A2(KEYINPUT26), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT26), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G190gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n242_), .A2(KEYINPUT25), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G183gat), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n248_), .A2(new_n250_), .A3(new_n251_), .A4(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(new_n239_), .ZN(new_n256_));
  INV_X1    g055(.A(G169gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n237_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(KEYINPUT24), .A3(new_n246_), .ZN(new_n259_));
  NOR3_X1   g058(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n254_), .A2(new_n256_), .A3(new_n259_), .A4(new_n261_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n247_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n211_), .B1(new_n235_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n246_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n266_), .B1(new_n256_), .B2(new_n244_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT22), .ZN(new_n268_));
  OAI21_X1  g067(.A(G169gat), .B1(new_n268_), .B2(KEYINPUT78), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT78), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(new_n257_), .A3(KEYINPUT22), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n271_), .A3(new_n237_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT79), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT79), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n269_), .A2(new_n271_), .A3(new_n274_), .A4(new_n237_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n267_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n260_), .B1(new_n278_), .B2(new_n246_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT25), .B(G183gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT77), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n248_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n279_), .B(new_n256_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n276_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT80), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n223_), .B1(new_n214_), .B2(G204gat), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n217_), .A2(KEYINPUT86), .A3(G197gat), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n226_), .B(new_n228_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT87), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n230_), .A2(KEYINPUT87), .A3(new_n226_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n233_), .B1(new_n294_), .B2(new_n221_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT80), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n276_), .A2(new_n285_), .A3(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n287_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n210_), .B1(new_n265_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n209_), .A2(new_n211_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n287_), .A2(new_n297_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(new_n235_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n232_), .A2(new_n234_), .A3(new_n263_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT91), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n295_), .A2(KEYINPUT91), .A3(new_n263_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n304_), .A2(new_n309_), .A3(KEYINPUT92), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT92), .B1(new_n304_), .B2(new_n309_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n206_), .B(new_n300_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT98), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT27), .ZN(new_n315_));
  XOR2_X1   g114(.A(KEYINPUT96), .B(KEYINPUT20), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n263_), .B(KEYINPUT97), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n316_), .B1(new_n317_), .B2(new_n235_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n276_), .A2(new_n296_), .A3(new_n285_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n296_), .B1(new_n276_), .B2(new_n285_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n235_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n209_), .B1(new_n318_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n265_), .A2(new_n298_), .A3(new_n210_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n315_), .B1(new_n325_), .B2(new_n205_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT92), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT91), .B1(new_n295_), .B2(new_n263_), .ZN(new_n328_));
  AND4_X1   g127(.A1(KEYINPUT91), .A2(new_n232_), .A3(new_n234_), .A4(new_n263_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n321_), .A2(new_n301_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n327_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n304_), .A2(new_n309_), .A3(KEYINPUT92), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n334_), .A2(KEYINPUT98), .A3(new_n206_), .A4(new_n300_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n314_), .A2(new_n326_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n206_), .B1(new_n334_), .B2(new_n300_), .ZN(new_n337_));
  AOI211_X1 g136(.A(new_n205_), .B(new_n299_), .C1(new_n332_), .C2(new_n333_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n315_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G78gat), .B(G106gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT88), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344_));
  OR3_X1    g143(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  OR3_X1    g146(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT2), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n348_), .A2(new_n351_), .A3(new_n352_), .A4(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n347_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(KEYINPUT1), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(G155gat), .A3(G162gat), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n345_), .A2(new_n357_), .A3(new_n359_), .A4(new_n346_), .ZN(new_n360_));
  INV_X1    g159(.A(G141gat), .ZN(new_n361_));
  INV_X1    g160(.A(G148gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n363_), .A3(new_n349_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n344_), .B1(new_n356_), .B2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT84), .B1(new_n295_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(G228gat), .ZN(new_n367_));
  INV_X1    g166(.A(G233gat), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n356_), .A2(new_n364_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT29), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n220_), .A2(KEYINPUT21), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n212_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n371_), .B(new_n372_), .C1(new_n375_), .C2(new_n233_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n366_), .A2(new_n369_), .A3(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n369_), .B1(new_n366_), .B2(new_n376_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n343_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n366_), .A2(new_n376_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n366_), .A2(new_n376_), .A3(new_n369_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n342_), .A3(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n385_));
  OR3_X1    g184(.A1(new_n370_), .A2(KEYINPUT29), .A3(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G22gat), .B(G50gat), .Z(new_n387_));
  OAI21_X1  g186(.A(new_n385_), .B1(new_n370_), .B2(KEYINPUT29), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n379_), .A2(new_n384_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT89), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n379_), .A2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(KEYINPUT89), .B(new_n343_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n395_));
  OR3_X1    g194(.A1(new_n377_), .A2(new_n378_), .A3(new_n343_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n391_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n392_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(G127gat), .B(G134gat), .Z(new_n401_));
  XOR2_X1   g200(.A(G113gat), .B(G120gat), .Z(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G127gat), .B(G134gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G113gat), .B(G120gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT81), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n403_), .A2(KEYINPUT81), .A3(new_n406_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT93), .B(KEYINPUT4), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n370_), .A2(new_n409_), .A3(new_n410_), .A4(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n370_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n356_), .A2(new_n407_), .A3(new_n364_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(KEYINPUT4), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT94), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n416_), .A2(new_n417_), .A3(new_n413_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT94), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n415_), .A2(new_n422_), .A3(new_n418_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(G85gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT0), .B(G57gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n426_), .B(new_n427_), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n424_), .A2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n420_), .A2(new_n421_), .A3(new_n423_), .A4(new_n428_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n341_), .A2(new_n400_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT95), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n435_), .A2(KEYINPUT33), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n431_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n418_), .A2(new_n413_), .A3(new_n412_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n416_), .A2(new_n417_), .A3(new_n414_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n429_), .A3(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(new_n431_), .B2(new_n436_), .ZN(new_n441_));
  NOR4_X1   g240(.A1(new_n337_), .A2(new_n437_), .A3(new_n441_), .A4(new_n338_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n300_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n325_), .A2(new_n444_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n433_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n399_), .B1(new_n442_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n434_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G227gat), .A2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(G15gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT30), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n303_), .B(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n409_), .A2(new_n410_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G71gat), .B(G99gat), .Z(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(G43gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT31), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n456_), .A2(new_n459_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n449_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n399_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT99), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n399_), .A2(new_n336_), .A3(new_n339_), .A4(KEYINPUT99), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n462_), .A2(new_n433_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT100), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT100), .ZN(new_n473_));
  AOI211_X1 g272(.A(new_n473_), .B(new_n470_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n464_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G29gat), .B(G36gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G43gat), .B(G50gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT74), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G15gat), .B(G22gat), .ZN(new_n480_));
  INV_X1    g279(.A(G1gat), .ZN(new_n481_));
  INV_X1    g280(.A(G8gat), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT14), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G1gat), .B(G8gat), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n484_), .B(new_n485_), .Z(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT74), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n478_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n486_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n487_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G229gat), .A2(G233gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT75), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n478_), .B(KEYINPUT15), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n490_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n487_), .A2(new_n498_), .A3(new_n493_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G113gat), .B(G141gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G169gat), .B(G197gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n496_), .A2(new_n499_), .A3(new_n503_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(KEYINPUT76), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT76), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n500_), .A2(new_n508_), .A3(new_n504_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n475_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT6), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT64), .ZN(new_n515_));
  INV_X1    g314(.A(G85gat), .ZN(new_n516_));
  INV_X1    g315(.A(G92gat), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n516_), .A2(new_n517_), .A3(KEYINPUT9), .ZN(new_n518_));
  XOR2_X1   g317(.A(G85gat), .B(G92gat), .Z(new_n519_));
  AOI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(KEYINPUT9), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT10), .B(G99gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(G106gat), .B2(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n515_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT8), .ZN(new_n524_));
  NOR3_X1   g323(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT7), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n524_), .B(new_n519_), .C1(new_n515_), .C2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n514_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n519_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT8), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n523_), .B1(new_n528_), .B2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G57gat), .B(G64gat), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n533_), .A2(KEYINPUT11), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(KEYINPUT11), .ZN(new_n535_));
  XOR2_X1   g334(.A(G71gat), .B(G78gat), .Z(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n535_), .A2(new_n536_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n532_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G230gat), .A2(G233gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT67), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n540_), .A2(KEYINPUT67), .A3(new_n541_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT12), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n528_), .A2(new_n531_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n523_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n539_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n546_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n532_), .A2(KEYINPUT12), .A3(new_n539_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n544_), .B(new_n545_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n541_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n540_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n532_), .A2(new_n539_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n554_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT66), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n557_), .A2(new_n558_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n553_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G120gat), .B(G148gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT5), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G176gat), .B(G204gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n563_), .B(new_n564_), .Z(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n565_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n553_), .B(new_n567_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT13), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n566_), .A2(KEYINPUT13), .A3(new_n568_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT72), .ZN(new_n575_));
  XOR2_X1   g374(.A(KEYINPUT71), .B(KEYINPUT16), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G127gat), .B(G155gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT17), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n486_), .B(new_n539_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(KEYINPUT17), .A3(new_n579_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT73), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n549_), .A2(new_n497_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n532_), .A2(new_n478_), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n589_), .B(new_n590_), .C1(KEYINPUT35), .C2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(KEYINPUT35), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G190gat), .B(G218gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT69), .ZN(new_n599_));
  XOR2_X1   g398(.A(G134gat), .B(G162gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n596_), .A2(new_n597_), .A3(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n597_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n602_), .B1(new_n596_), .B2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT70), .B(KEYINPUT37), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AND4_X1   g406(.A1(new_n512_), .A2(new_n573_), .A3(new_n588_), .A4(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(new_n481_), .A3(new_n432_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT38), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n604_), .B(KEYINPUT101), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n475_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n573_), .A2(new_n511_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n614_), .A2(new_n586_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n481_), .B1(new_n616_), .B2(new_n432_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n611_), .A2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n618_), .B1(new_n610_), .B2(new_n609_), .ZN(G1324gat));
  AOI21_X1  g418(.A(new_n482_), .B1(new_n616_), .B2(new_n340_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT39), .Z(new_n621_));
  NAND3_X1  g420(.A1(new_n608_), .A2(new_n482_), .A3(new_n340_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n621_), .A2(KEYINPUT40), .A3(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1325gat));
  INV_X1    g426(.A(KEYINPUT41), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n616_), .A2(new_n462_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(G15gat), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n630_), .B1(new_n629_), .B2(G15gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n628_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n633_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(KEYINPUT41), .A3(new_n631_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n608_), .A2(new_n451_), .A3(new_n462_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT103), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n634_), .A2(new_n636_), .A3(new_n640_), .A4(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(G1326gat));
  INV_X1    g441(.A(G22gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n399_), .B(KEYINPUT104), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n616_), .B2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT42), .Z(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n643_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT105), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n608_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(G1327gat));
  NAND2_X1  g449(.A1(new_n612_), .A2(new_n587_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n573_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n512_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n433_), .A2(G29gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT107), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n615_), .A2(new_n588_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n475_), .A2(new_n660_), .A3(new_n606_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n475_), .B2(new_n606_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT44), .B(new_n659_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n432_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G29gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G29gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n658_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT108), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n673_), .B(new_n658_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1328gat));
  NOR3_X1   g474(.A1(new_n654_), .A2(G36gat), .A3(new_n341_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT45), .Z(new_n677_));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n665_), .A2(new_n666_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(new_n340_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n665_), .A2(new_n678_), .A3(new_n340_), .A4(new_n666_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G36gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n677_), .B1(new_n680_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT46), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(KEYINPUT46), .B(new_n677_), .C1(new_n680_), .C2(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1329gat));
  NAND3_X1  g486(.A1(new_n679_), .A2(G43gat), .A3(new_n462_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT110), .B(G43gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n654_), .B2(new_n463_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g491(.A(G50gat), .B1(new_n655_), .B2(new_n644_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n400_), .A2(G50gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n679_), .B2(new_n694_), .ZN(G1331gat));
  NOR2_X1   g494(.A1(new_n511_), .A2(new_n587_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n614_), .A2(new_n573_), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G57gat), .B1(new_n699_), .B2(new_n433_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n475_), .A2(new_n510_), .ZN(new_n701_));
  NOR4_X1   g500(.A1(new_n701_), .A2(new_n573_), .A3(new_n587_), .A4(new_n606_), .ZN(new_n702_));
  INV_X1    g501(.A(G57gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n432_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n700_), .A2(new_n704_), .ZN(G1332gat));
  INV_X1    g504(.A(G64gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n698_), .B2(new_n340_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT48), .Z(new_n708_));
  NAND3_X1  g507(.A1(new_n702_), .A2(new_n706_), .A3(new_n340_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1333gat));
  INV_X1    g509(.A(G71gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n698_), .B2(new_n462_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n702_), .A2(new_n711_), .A3(new_n462_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1334gat));
  INV_X1    g515(.A(G78gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n698_), .B2(new_n644_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT50), .Z(new_n719_));
  NAND3_X1  g518(.A1(new_n702_), .A2(new_n717_), .A3(new_n644_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1335gat));
  NOR3_X1   g520(.A1(new_n701_), .A2(new_n573_), .A3(new_n651_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(new_n516_), .A3(new_n432_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n661_), .A2(new_n662_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n573_), .A2(new_n511_), .A3(new_n588_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(new_n432_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n727_), .B2(new_n516_), .ZN(G1336gat));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n340_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n341_), .A2(G92gat), .ZN(new_n730_));
  AOI22_X1  g529(.A1(new_n729_), .A2(G92gat), .B1(new_n722_), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT112), .ZN(G1337gat));
  INV_X1    g531(.A(new_n521_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n722_), .A2(new_n462_), .A3(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT113), .Z(new_n735_));
  INV_X1    g534(.A(G99gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n726_), .B2(new_n462_), .ZN(new_n737_));
  OR3_X1    g536(.A1(new_n735_), .A2(KEYINPUT51), .A3(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT51), .B1(new_n735_), .B2(new_n737_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1338gat));
  NAND3_X1  g539(.A1(new_n724_), .A2(new_n400_), .A3(new_n725_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G106gat), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n741_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n745_));
  INV_X1    g544(.A(G106gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n722_), .A2(new_n746_), .A3(new_n400_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT114), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n744_), .A2(new_n745_), .A3(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g549(.A1(new_n469_), .A2(new_n432_), .A3(new_n462_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n751_), .A2(KEYINPUT59), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT57), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n545_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT67), .B1(new_n540_), .B2(new_n541_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT118), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT55), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n553_), .A2(KEYINPUT118), .A3(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n540_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT119), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n554_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n554_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT119), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n757_), .A2(new_n759_), .A3(new_n762_), .A4(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n565_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n565_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n507_), .A2(new_n509_), .A3(new_n568_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n507_), .A2(KEYINPUT117), .A3(new_n509_), .A4(new_n568_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n506_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n487_), .A2(new_n498_), .A3(new_n494_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n503_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n569_), .A2(new_n779_), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n753_), .B(new_n612_), .C1(new_n775_), .C2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n773_), .A2(new_n774_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n769_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n565_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n780_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT57), .B1(new_n786_), .B2(new_n613_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n781_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n779_), .A2(new_n568_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n606_), .B1(new_n790_), .B2(KEYINPUT58), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(KEYINPUT58), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n606_), .B(KEYINPUT120), .C1(new_n790_), .C2(KEYINPUT58), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n588_), .B1(new_n788_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n573_), .A2(new_n798_), .A3(new_n696_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n607_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n573_), .B2(new_n696_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  OR3_X1    g602(.A1(new_n800_), .A2(new_n801_), .A3(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n752_), .B1(new_n797_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n786_), .A2(new_n613_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n753_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n786_), .A2(KEYINPUT57), .A3(new_n613_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n586_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n804_), .A2(new_n805_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n751_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT59), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n807_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(G113gat), .B1(new_n817_), .B2(new_n510_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n751_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n586_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n788_), .B2(new_n796_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n821_), .B2(new_n806_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n510_), .A2(G113gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n818_), .B1(new_n822_), .B2(new_n823_), .ZN(G1340gat));
  NOR2_X1   g623(.A1(new_n817_), .A2(new_n573_), .ZN(new_n825_));
  XOR2_X1   g624(.A(KEYINPUT121), .B(G120gat), .Z(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n573_), .B2(KEYINPUT60), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(KEYINPUT60), .B2(new_n826_), .ZN(new_n828_));
  OAI22_X1  g627(.A1(new_n825_), .A2(new_n826_), .B1(new_n822_), .B2(new_n828_), .ZN(G1341gat));
  INV_X1    g628(.A(KEYINPUT122), .ZN(new_n830_));
  INV_X1    g629(.A(G127gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n587_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n814_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n822_), .A2(KEYINPUT59), .B1(new_n833_), .B2(new_n752_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n831_), .B1(new_n834_), .B2(new_n820_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n822_), .A2(G127gat), .A3(new_n587_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n830_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(G127gat), .B1(new_n817_), .B2(new_n586_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n836_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(KEYINPUT122), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(G1342gat));
  AOI21_X1  g640(.A(G134gat), .B1(new_n815_), .B2(new_n612_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n606_), .A2(G134gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(KEYINPUT123), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n842_), .B1(new_n834_), .B2(new_n844_), .ZN(G1343gat));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n821_), .A2(new_n806_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n341_), .A2(new_n400_), .A3(new_n432_), .A4(new_n463_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n847_), .A2(new_n846_), .A3(new_n848_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G141gat), .B1(new_n852_), .B2(new_n510_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n361_), .B(new_n511_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1344gat));
  OAI21_X1  g654(.A(G148gat), .B1(new_n852_), .B2(new_n573_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n362_), .B(new_n652_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1345gat));
  XNOR2_X1  g657(.A(KEYINPUT61), .B(G155gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n852_), .B2(new_n587_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n859_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n588_), .B(new_n861_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1346gat));
  INV_X1    g662(.A(new_n851_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n607_), .B1(new_n864_), .B2(new_n849_), .ZN(new_n865_));
  INV_X1    g664(.A(G162gat), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n612_), .A2(new_n866_), .ZN(new_n867_));
  OAI22_X1  g666(.A1(new_n865_), .A2(new_n866_), .B1(new_n852_), .B2(new_n867_), .ZN(G1347gat));
  NOR2_X1   g667(.A1(new_n341_), .A2(new_n470_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  AOI211_X1 g669(.A(new_n644_), .B(new_n870_), .C1(new_n832_), .C2(new_n814_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n257_), .B1(new_n871_), .B2(new_n511_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n872_), .A2(KEYINPUT62), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n871_), .A2(new_n236_), .A3(new_n511_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(KEYINPUT62), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n873_), .A2(new_n874_), .A3(new_n875_), .ZN(G1348gat));
  AOI21_X1  g675(.A(G176gat), .B1(new_n871_), .B2(new_n652_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n847_), .A2(new_n400_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n573_), .A2(new_n870_), .A3(new_n237_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n878_), .B2(new_n879_), .ZN(G1349gat));
  NAND3_X1  g679(.A1(new_n878_), .A2(new_n588_), .A3(new_n869_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n586_), .A2(new_n280_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n881_), .A2(new_n242_), .B1(new_n871_), .B2(new_n882_), .ZN(G1350gat));
  NAND4_X1  g682(.A1(new_n871_), .A2(new_n248_), .A3(new_n250_), .A4(new_n612_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n871_), .A2(new_n606_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n243_), .ZN(G1351gat));
  NAND4_X1  g685(.A1(new_n463_), .A2(new_n340_), .A3(new_n400_), .A4(new_n433_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n847_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n511_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n214_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT125), .B(G197gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n889_), .B2(new_n892_), .ZN(G1352gat));
  NAND2_X1  g692(.A1(new_n888_), .A2(new_n652_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g694(.A(KEYINPUT126), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n586_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n888_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n896_), .B1(new_n888_), .B2(new_n897_), .ZN(new_n900_));
  OAI22_X1  g699(.A1(new_n899_), .A2(new_n900_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n901_));
  INV_X1    g700(.A(new_n900_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n902_), .A2(new_n903_), .A3(new_n898_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n904_), .ZN(G1354gat));
  INV_X1    g704(.A(G218gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n888_), .A2(new_n906_), .A3(new_n612_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n847_), .A2(new_n607_), .A3(new_n887_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n906_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n907_), .B(KEYINPUT127), .C1(new_n906_), .C2(new_n908_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1355gat));
endmodule


