//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_;
  INV_X1    g000(.A(KEYINPUT107), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  INV_X1    g003(.A(G8gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G29gat), .B(G36gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n209_), .B(new_n212_), .Z(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G229gat), .A3(G233gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n212_), .B(KEYINPUT15), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(new_n209_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n209_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(new_n212_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G229gat), .A2(G233gat), .ZN(new_n219_));
  XOR2_X1   g018(.A(new_n219_), .B(KEYINPUT81), .Z(new_n220_));
  NAND3_X1  g019(.A1(new_n216_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n214_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(G113gat), .B(G141gat), .Z(new_n223_));
  XNOR2_X1  g022(.A(G169gat), .B(G197gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n222_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT71), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(G85gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G92gat), .ZN(new_n230_));
  OR3_X1    g029(.A1(new_n229_), .A2(KEYINPUT9), .A3(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G85gat), .B(G92gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT9), .ZN(new_n234_));
  XOR2_X1   g033(.A(KEYINPUT10), .B(G99gat), .Z(new_n235_));
  INV_X1    g034(.A(G106gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G99gat), .A2(G106gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT6), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n231_), .A2(new_n234_), .A3(new_n237_), .A4(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244_));
  NOR2_X1   g043(.A1(G99gat), .A2(G106gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT7), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT7), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT65), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n245_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  AOI211_X1 g049(.A(G99gat), .B(G106gat), .C1(new_n246_), .C2(KEYINPUT7), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n244_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(new_n245_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT65), .B(KEYINPUT7), .ZN(new_n254_));
  OAI211_X1 g053(.A(KEYINPUT66), .B(new_n253_), .C1(new_n254_), .C2(new_n245_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n252_), .A2(new_n241_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n233_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(KEYINPUT67), .A3(new_n233_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT8), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT8), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n253_), .B1(new_n254_), .B2(new_n245_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n262_), .B(new_n233_), .C1(new_n263_), .C2(new_n240_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n243_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n215_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n227_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n264_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n240_), .B1(new_n263_), .B2(new_n244_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n232_), .B1(new_n269_), .B2(new_n255_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n262_), .B1(new_n270_), .B2(KEYINPUT67), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n268_), .B1(new_n271_), .B2(new_n259_), .ZN(new_n272_));
  OAI211_X1 g071(.A(KEYINPUT71), .B(new_n215_), .C1(new_n272_), .C2(new_n243_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n265_), .A2(new_n212_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n267_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT35), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n267_), .A2(new_n273_), .A3(new_n278_), .A4(new_n274_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G232gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(new_n279_), .A3(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n279_), .A2(new_n282_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G190gat), .B(G218gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G134gat), .B(G162gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT74), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n283_), .A2(new_n284_), .A3(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n279_), .A2(new_n282_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n279_), .A2(new_n282_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n293_), .B1(new_n294_), .B2(new_n277_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n287_), .B(KEYINPUT36), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n292_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT85), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT2), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n299_), .A2(KEYINPUT85), .A3(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n301_), .A2(new_n303_), .A3(new_n306_), .A4(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G155gat), .B(G162gat), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n304_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n313_), .A2(new_n299_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT28), .B1(new_n317_), .B2(KEYINPUT29), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n308_), .A2(new_n309_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT28), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT29), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT86), .ZN(new_n324_));
  XOR2_X1   g123(.A(G22gat), .B(G50gat), .Z(new_n325_));
  INV_X1    g124(.A(KEYINPUT86), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n318_), .A2(new_n326_), .A3(new_n322_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n327_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n325_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G78gat), .B(G106gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G218gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(G211gat), .ZN(new_n335_));
  INV_X1    g134(.A(G211gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G218gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT87), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G211gat), .B(G218gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT87), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(G197gat), .A2(G204gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G197gat), .A2(G204gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(KEYINPUT21), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n343_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n345_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT21), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n351_), .A2(new_n339_), .A3(new_n342_), .A4(new_n346_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(G228gat), .ZN(new_n354_));
  INV_X1    g153(.A(G233gat), .ZN(new_n355_));
  OAI221_X1 g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .C1(new_n321_), .C2(new_n319_), .ZN(new_n356_));
  XOR2_X1   g155(.A(KEYINPUT88), .B(KEYINPUT29), .Z(new_n357_));
  OAI21_X1  g156(.A(new_n353_), .B1(new_n319_), .B2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n354_), .A2(new_n355_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(KEYINPUT89), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT89), .B1(new_n358_), .B2(new_n359_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n333_), .B(new_n356_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n328_), .A2(new_n331_), .B1(new_n363_), .B2(KEYINPUT91), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n363_), .A2(KEYINPUT91), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n356_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(KEYINPUT90), .A3(new_n332_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT90), .ZN(new_n368_));
  INV_X1    g167(.A(new_n356_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n362_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n360_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n368_), .B1(new_n371_), .B2(new_n333_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n364_), .A2(new_n365_), .A3(new_n367_), .A4(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n371_), .A2(new_n333_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n363_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n328_), .B(new_n331_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G71gat), .B(G99gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G43gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT31), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G127gat), .B(G134gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G113gat), .B(G120gat), .Z(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G113gat), .B(G120gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n383_), .A2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n382_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n382_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n381_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G15gat), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n395_), .B(KEYINPUT30), .Z(new_n396_));
  XNOR2_X1  g195(.A(new_n393_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT25), .B(G183gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT26), .B(G190gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT24), .ZN(new_n400_));
  NOR2_X1   g199(.A1(G169gat), .A2(G176gat), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n398_), .A2(new_n399_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G169gat), .ZN(new_n403_));
  INV_X1    g202(.A(G176gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  OR3_X1    g204(.A1(new_n405_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G183gat), .A2(G190gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT82), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(G183gat), .A3(G190gat), .ZN(new_n411_));
  AOI21_X1  g210(.A(KEYINPUT23), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT23), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(G183gat), .B2(G190gat), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n407_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G169gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n408_), .A2(new_n413_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n409_), .A2(new_n411_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(KEYINPUT23), .ZN(new_n423_));
  NOR2_X1   g222(.A1(G183gat), .A2(G190gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n419_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n416_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT84), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n397_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n397_), .A2(new_n429_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n383_), .B(new_n387_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n319_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G225gat), .A2(G233gat), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n434_), .B(new_n435_), .C1(new_n392_), .C2(new_n319_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT99), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n390_), .B1(new_n433_), .B2(new_n382_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n317_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT99), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n435_), .A4(new_n434_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT4), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n438_), .A2(new_n443_), .A3(new_n317_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT98), .ZN(new_n445_));
  INV_X1    g244(.A(new_n435_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n434_), .B(KEYINPUT4), .C1(new_n392_), .C2(new_n319_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT98), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n438_), .A2(new_n448_), .A3(new_n317_), .A4(new_n443_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .A4(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n442_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G1gat), .B(G29gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(G85gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT0), .B(G57gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n453_), .B(new_n454_), .Z(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n451_), .A2(new_n456_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n450_), .A2(new_n455_), .A3(new_n437_), .A4(new_n441_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n432_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT96), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n422_), .A2(KEYINPUT23), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n420_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n407_), .A2(new_n463_), .ZN(new_n464_));
  OAI211_X1 g263(.A(KEYINPUT95), .B(new_n425_), .C1(new_n412_), .C2(new_n414_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n425_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT95), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n419_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n464_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n348_), .A2(new_n352_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n461_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n465_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n464_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(KEYINPUT96), .A3(new_n353_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n418_), .B1(new_n463_), .B2(new_n424_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n402_), .B(new_n406_), .C1(new_n414_), .C2(new_n412_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n476_), .A2(new_n352_), .A3(new_n348_), .A4(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(KEYINPUT20), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n479_), .B1(new_n478_), .B2(KEYINPUT20), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n471_), .B(new_n475_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G226gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n486_), .B(KEYINPUT93), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n472_), .A2(new_n473_), .A3(new_n470_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n490_), .A2(KEYINPUT20), .A3(new_n486_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT97), .B1(new_n427_), .B2(new_n470_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT97), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n493_), .B(new_n353_), .C1(new_n416_), .C2(new_n426_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n489_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G8gat), .B(G36gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT18), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G64gat), .B(G92gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n489_), .A2(new_n501_), .A3(new_n496_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT27), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(KEYINPUT27), .ZN(new_n506_));
  INV_X1    g305(.A(new_n486_), .ZN(new_n507_));
  XOR2_X1   g306(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n509_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n495_), .B1(new_n510_), .B2(KEYINPUT102), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n490_), .A2(new_n508_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT102), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n507_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n471_), .A2(new_n475_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n516_), .B(new_n487_), .C1(new_n482_), .C2(new_n481_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n501_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT103), .B1(new_n506_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT27), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n483_), .A2(new_n488_), .B1(new_n495_), .B2(new_n491_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n520_), .B1(new_n521_), .B2(new_n501_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n483_), .A2(new_n488_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n512_), .A2(new_n513_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n510_), .A2(KEYINPUT102), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n486_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n502_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT103), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n522_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  AOI211_X1 g328(.A(KEYINPUT104), .B(new_n505_), .C1(new_n519_), .C2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT104), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n519_), .A2(new_n529_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n505_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n378_), .B(new_n460_), .C1(new_n530_), .C2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n459_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n529_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n528_), .B1(new_n522_), .B2(new_n527_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n533_), .B(new_n536_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n445_), .A2(new_n435_), .A3(new_n447_), .A4(new_n449_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n439_), .A2(new_n446_), .A3(new_n434_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n541_), .A2(new_n456_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n458_), .A2(KEYINPUT33), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT33), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n442_), .A2(new_n545_), .A3(new_n455_), .A4(new_n450_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n543_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n503_), .A2(new_n547_), .A3(new_n504_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT100), .ZN(new_n549_));
  OAI211_X1 g348(.A(KEYINPUT32), .B(new_n501_), .C1(new_n523_), .C2(new_n526_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n501_), .A2(KEYINPUT32), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n458_), .A2(new_n457_), .B1(new_n521_), .B2(new_n551_), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n548_), .A2(new_n549_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n503_), .A2(new_n547_), .A3(KEYINPUT100), .A4(new_n504_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n377_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n432_), .B1(new_n540_), .B2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n298_), .B1(new_n535_), .B2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G57gat), .B(G64gat), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n558_), .A2(KEYINPUT11), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(KEYINPUT11), .ZN(new_n560_));
  XOR2_X1   g359(.A(G71gat), .B(G78gat), .Z(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n560_), .A2(new_n561_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n260_), .A2(KEYINPUT8), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT67), .B1(new_n256_), .B2(new_n233_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n264_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n570_), .A2(new_n564_), .A3(new_n242_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n564_), .B1(new_n570_), .B2(new_n242_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n567_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n565_), .B1(new_n272_), .B2(new_n243_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(KEYINPUT68), .A3(new_n566_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT68), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n572_), .B2(KEYINPUT12), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n573_), .A2(new_n575_), .A3(new_n577_), .A4(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n570_), .A2(new_n564_), .A3(new_n242_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n574_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n578_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G120gat), .B(G148gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(G176gat), .B(G204gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n584_), .A2(KEYINPUT69), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n584_), .B1(KEYINPUT69), .B2(new_n589_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT13), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT13), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n564_), .B(new_n597_), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT77), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(new_n217_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G183gat), .B(G211gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT79), .ZN(new_n602_));
  XOR2_X1   g401(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(G127gat), .B(G155gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT17), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n606_), .A2(new_n607_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n600_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n608_), .B2(new_n600_), .ZN(new_n611_));
  AND4_X1   g410(.A1(new_n226_), .A2(new_n557_), .A3(new_n596_), .A4(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n459_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(G1gat), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n297_), .A2(KEYINPUT37), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT76), .B1(new_n295_), .B2(new_n296_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n296_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT76), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n292_), .A2(KEYINPUT75), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT75), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n295_), .A2(new_n621_), .A3(new_n291_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n616_), .A2(new_n619_), .A3(new_n620_), .A4(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n615_), .B1(new_n623_), .B2(KEYINPUT37), .ZN(new_n624_));
  INV_X1    g423(.A(new_n611_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT80), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n226_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n593_), .A2(new_n595_), .ZN(new_n630_));
  AOI211_X1 g429(.A(new_n629_), .B(new_n630_), .C1(new_n535_), .C2(new_n556_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT105), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(KEYINPUT105), .A3(new_n631_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n459_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(G1gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(new_n635_), .A3(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n614_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n628_), .A2(KEYINPUT105), .A3(new_n631_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT105), .B1(new_n628_), .B2(new_n631_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n639_), .B1(new_n644_), .B2(new_n637_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n202_), .B1(new_n641_), .B2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n638_), .A2(new_n640_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n647_), .A2(new_n648_), .A3(KEYINPUT107), .A4(new_n614_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(G1324gat));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n530_), .A2(new_n534_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n612_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G8gat), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT39), .Z(new_n655_));
  NAND2_X1  g454(.A1(new_n634_), .A2(new_n635_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(new_n205_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n651_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n654_), .B(KEYINPUT39), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n660_), .B(KEYINPUT40), .C1(new_n656_), .C2(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(G1325gat));
  INV_X1    g461(.A(new_n432_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n612_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G15gat), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT41), .Z(new_n666_));
  OR2_X1    g465(.A1(new_n432_), .A2(G15gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n656_), .B2(new_n667_), .ZN(G1326gat));
  NAND2_X1  g467(.A1(new_n612_), .A2(new_n377_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G22gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT42), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n378_), .A2(G22gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n656_), .B2(new_n672_), .ZN(G1327gat));
  NAND2_X1  g472(.A1(new_n535_), .A2(new_n556_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(new_n624_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n674_), .A2(KEYINPUT108), .A3(new_n675_), .A4(new_n624_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n674_), .A2(new_n624_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT43), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n678_), .A2(new_n679_), .A3(new_n681_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n630_), .A2(new_n629_), .A3(new_n611_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(KEYINPUT44), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT44), .B1(new_n682_), .B2(new_n683_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G29gat), .B1(new_n687_), .B2(new_n636_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n611_), .A2(new_n297_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n631_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n636_), .A2(G29gat), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT109), .Z(new_n693_));
  OAI21_X1  g492(.A(new_n688_), .B1(new_n691_), .B2(new_n693_), .ZN(G1328gat));
  INV_X1    g493(.A(G36gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n690_), .A2(new_n695_), .A3(new_n652_), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n652_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n684_), .A2(new_n685_), .A3(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n700_), .B2(new_n695_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT46), .B(new_n698_), .C1(new_n700_), .C2(new_n695_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1329gat));
  NAND2_X1  g504(.A1(new_n663_), .A2(G43gat), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n684_), .A2(new_n685_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G43gat), .B1(new_n690_), .B2(new_n663_), .ZN(new_n708_));
  OR3_X1    g507(.A1(new_n707_), .A2(KEYINPUT47), .A3(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT47), .B1(new_n707_), .B2(new_n708_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n690_), .B2(new_n377_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n377_), .A2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n686_), .B2(new_n713_), .ZN(G1331gat));
  NAND2_X1  g513(.A1(new_n630_), .A2(new_n629_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n556_), .B2(new_n535_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n628_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(G57gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n459_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n715_), .A2(new_n625_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(new_n557_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G57gat), .B1(new_n722_), .B2(new_n636_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n719_), .A2(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n721_), .B2(new_n652_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT48), .Z(new_n727_));
  NAND3_X1  g526(.A1(new_n717_), .A2(new_n725_), .A3(new_n652_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1333gat));
  INV_X1    g528(.A(G71gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n721_), .B2(new_n663_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT49), .Z(new_n732_));
  NAND3_X1  g531(.A1(new_n717_), .A2(new_n730_), .A3(new_n663_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1334gat));
  INV_X1    g533(.A(G78gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n721_), .B2(new_n377_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT111), .Z(new_n737_));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n738_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n717_), .A2(new_n735_), .A3(new_n377_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n739_), .A2(new_n740_), .A3(new_n741_), .ZN(G1335gat));
  NAND2_X1  g541(.A1(new_n716_), .A2(new_n689_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G85gat), .B1(new_n744_), .B2(new_n459_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n715_), .A2(new_n611_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n682_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n636_), .A2(new_n229_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(G1336gat));
  NOR3_X1   g548(.A1(new_n743_), .A2(G92gat), .A3(new_n699_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n652_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(G92gat), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT112), .ZN(G1337gat));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n682_), .A2(new_n663_), .A3(new_n746_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(G99gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n744_), .A2(new_n663_), .A3(new_n235_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n754_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(new_n754_), .A3(new_n757_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n759_), .A2(KEYINPUT113), .A3(KEYINPUT51), .A4(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n762_));
  INV_X1    g561(.A(new_n760_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n758_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(new_n764_), .ZN(G1338gat));
  XNOR2_X1  g564(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n682_), .A2(new_n377_), .A3(new_n746_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G106gat), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT52), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n770_), .A3(G106gat), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n744_), .A2(new_n236_), .A3(new_n377_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n766_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n767_), .A2(new_n770_), .A3(G106gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n770_), .B1(new_n767_), .B2(G106gat), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n773_), .B(new_n766_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n774_), .A2(new_n778_), .ZN(G1339gat));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n573_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n582_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n579_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n781_), .A2(new_n780_), .A3(new_n582_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n589_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT56), .ZN(new_n787_));
  INV_X1    g586(.A(new_n589_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n579_), .A2(new_n583_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n220_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n216_), .A2(new_n218_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n225_), .B1(new_n213_), .B2(new_n220_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n222_), .A2(new_n225_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT119), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n796_), .B(new_n589_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n787_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT58), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n787_), .A2(new_n795_), .A3(KEYINPUT58), .A4(new_n797_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n624_), .A3(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n566_), .B1(new_n265_), .B2(new_n564_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n581_), .A2(new_n567_), .B1(new_n803_), .B2(new_n576_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n578_), .B1(new_n804_), .B2(new_n575_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n579_), .B1(new_n805_), .B2(new_n780_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n785_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n788_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n796_), .B1(new_n808_), .B2(KEYINPUT118), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n786_), .A2(new_n810_), .A3(KEYINPUT56), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n789_), .A2(new_n226_), .ZN(new_n812_));
  XOR2_X1   g611(.A(new_n812_), .B(KEYINPUT117), .Z(new_n813_));
  NAND3_X1  g612(.A1(new_n809_), .A2(new_n811_), .A3(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n793_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n298_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n802_), .B1(new_n816_), .B2(KEYINPUT57), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n818_), .B(new_n298_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n625_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  XOR2_X1   g619(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n821_));
  NOR2_X1   g620(.A1(new_n630_), .A2(new_n226_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n626_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n626_), .B2(new_n822_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n820_), .A2(new_n825_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n652_), .A2(new_n377_), .A3(new_n432_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n459_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(G113gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n226_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n828_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n636_), .B1(new_n820_), .B2(new_n825_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(KEYINPUT59), .A3(new_n827_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n629_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n831_), .B1(new_n836_), .B2(new_n830_), .ZN(G1340gat));
  XOR2_X1   g636(.A(KEYINPUT120), .B(G120gat), .Z(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n596_), .B2(KEYINPUT60), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n829_), .B(new_n839_), .C1(KEYINPUT60), .C2(new_n838_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n596_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n838_), .ZN(G1341gat));
  INV_X1    g641(.A(G127gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n828_), .B2(new_n625_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT121), .B(new_n843_), .C1(new_n828_), .C2(new_n625_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n833_), .A2(new_n835_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n625_), .A2(new_n843_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n846_), .A2(new_n847_), .B1(new_n848_), .B2(new_n849_), .ZN(G1342gat));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n828_), .B2(new_n297_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT122), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n854_), .B(new_n851_), .C1(new_n828_), .C2(new_n297_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n624_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n851_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n853_), .A2(new_n855_), .B1(new_n848_), .B2(new_n857_), .ZN(G1343gat));
  NOR3_X1   g657(.A1(new_n652_), .A2(new_n378_), .A3(new_n663_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n834_), .A2(new_n226_), .A3(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g660(.A1(new_n834_), .A2(new_n630_), .A3(new_n859_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g662(.A1(new_n834_), .A2(new_n611_), .A3(new_n859_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT61), .B(G155gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT123), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n864_), .B(new_n866_), .ZN(G1346gat));
  AND2_X1   g666(.A1(new_n834_), .A2(new_n859_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G162gat), .B1(new_n868_), .B2(new_n298_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n624_), .A2(G162gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT124), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n868_), .B2(new_n871_), .ZN(G1347gat));
  AOI21_X1  g671(.A(new_n699_), .B1(new_n820_), .B2(new_n825_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT22), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n460_), .A2(new_n378_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n873_), .A2(new_n874_), .A3(new_n226_), .A4(new_n876_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n877_), .A2(KEYINPUT62), .A3(new_n403_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(KEYINPUT62), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n873_), .A2(new_n226_), .A3(new_n876_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n403_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n878_), .B1(new_n879_), .B2(new_n882_), .ZN(G1348gat));
  NAND2_X1  g682(.A1(new_n873_), .A2(new_n876_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n596_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n404_), .ZN(G1349gat));
  NAND3_X1  g685(.A1(new_n873_), .A2(new_n611_), .A3(new_n876_), .ZN(new_n887_));
  MUX2_X1   g686(.A(new_n398_), .B(G183gat), .S(new_n887_), .Z(G1350gat));
  OAI21_X1  g687(.A(G190gat), .B1(new_n884_), .B2(new_n856_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n298_), .A2(new_n399_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n884_), .B2(new_n890_), .ZN(G1351gat));
  NAND2_X1  g690(.A1(new_n536_), .A2(new_n432_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT125), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n873_), .A2(new_n226_), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(G197gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(KEYINPUT126), .B2(new_n895_), .ZN(new_n896_));
  XOR2_X1   g695(.A(KEYINPUT126), .B(G197gat), .Z(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n894_), .B2(new_n897_), .ZN(G1352gat));
  AND2_X1   g697(.A1(new_n873_), .A2(new_n893_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n630_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(G204gat), .ZN(new_n901_));
  INV_X1    g700(.A(G204gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n899_), .A2(new_n902_), .A3(new_n630_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1353gat));
  NAND3_X1  g703(.A1(new_n873_), .A2(new_n611_), .A3(new_n893_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  AND2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n905_), .B2(new_n906_), .ZN(G1354gat));
  AOI21_X1  g708(.A(G218gat), .B1(new_n899_), .B2(new_n298_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n624_), .A2(G218gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT127), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n899_), .B2(new_n912_), .ZN(G1355gat));
endmodule


