//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT10), .B(G99gat), .Z(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT64), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n206_), .A2(KEYINPUT64), .ZN(new_n210_));
  OR2_X1    g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n210_), .A2(new_n208_), .A3(new_n207_), .A4(new_n211_), .ZN(new_n212_));
  AND3_X1   g011(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n205_), .A2(new_n209_), .A3(new_n212_), .A4(new_n215_), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n211_), .A2(new_n208_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n219_), .A3(new_n204_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n215_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n221_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n225_));
  OAI211_X1 g024(.A(KEYINPUT8), .B(new_n217_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT6), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n220_), .A2(new_n229_), .A3(new_n230_), .A4(new_n222_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(new_n217_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n226_), .A2(KEYINPUT67), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT67), .B1(new_n226_), .B2(new_n234_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n216_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G43gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT70), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G43gat), .ZN(new_n241_));
  INV_X1    g040(.A(G50gat), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n239_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n242_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G29gat), .B(G36gat), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n245_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n240_), .A2(G43gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n238_), .A2(KEYINPUT70), .ZN(new_n249_));
  OAI21_X1  g048(.A(G50gat), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n239_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n247_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT71), .B1(new_n246_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n245_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n247_), .A3(new_n251_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT71), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n253_), .A2(KEYINPUT15), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT15), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n254_), .A2(new_n256_), .A3(new_n255_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n256_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n237_), .A2(new_n258_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G232gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT34), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n265_), .A2(KEYINPUT35), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n226_), .A2(new_n216_), .A3(new_n234_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n226_), .A2(KEYINPUT66), .A3(new_n216_), .A4(new_n234_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n254_), .A2(new_n255_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n265_), .A2(KEYINPUT35), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n275_), .B(KEYINPUT75), .Z(new_n276_));
  NAND4_X1  g075(.A1(new_n263_), .A2(new_n266_), .A3(new_n274_), .A4(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT76), .ZN(new_n278_));
  NOR3_X1   g077(.A1(new_n260_), .A2(new_n261_), .A3(new_n259_), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT15), .B1(new_n253_), .B2(new_n257_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n281_), .A2(new_n237_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT76), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(new_n266_), .A4(new_n276_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n278_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(new_n282_), .B2(new_n275_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n275_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n262_), .A2(new_n258_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n236_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n226_), .A2(KEYINPUT67), .A3(new_n234_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n289_), .B1(new_n216_), .B2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n272_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n294_));
  OAI211_X1 g093(.A(KEYINPUT72), .B(new_n288_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n287_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n285_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G190gat), .B(G218gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G134gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(G162gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n297_), .A2(KEYINPUT36), .A3(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(KEYINPUT36), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n278_), .A2(new_n284_), .B1(new_n287_), .B2(new_n295_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  AND4_X1   g104(.A1(new_n285_), .A2(new_n296_), .A3(new_n302_), .A4(new_n304_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n202_), .B(new_n301_), .C1(new_n305_), .C2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n285_), .A2(new_n296_), .A3(new_n304_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n302_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n285_), .A2(new_n296_), .A3(new_n302_), .A4(new_n304_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n202_), .B1(new_n313_), .B2(new_n301_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT84), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n317_), .B(new_n318_), .C1(G141gat), .C2(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(G141gat), .ZN(new_n320_));
  INV_X1    g119(.A(G148gat), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n320_), .B(new_n321_), .C1(KEYINPUT84), .C2(KEYINPUT3), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n319_), .A2(new_n322_), .B1(KEYINPUT84), .B2(KEYINPUT3), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G141gat), .A2(G148gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT2), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n328_), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n332_), .A2(KEYINPUT1), .B1(new_n320_), .B2(new_n321_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n327_), .A2(new_n334_), .A3(new_n328_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n324_), .A3(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G127gat), .B(G134gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G113gat), .ZN(new_n338_));
  OR2_X1    g137(.A1(G127gat), .A2(G134gat), .ZN(new_n339_));
  INV_X1    g138(.A(G113gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G127gat), .A2(G134gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n338_), .A2(G120gat), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G120gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n342_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n340_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n344_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n331_), .A2(new_n336_), .A3(new_n343_), .A4(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n329_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n336_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n345_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n351_));
  AOI21_X1  g150(.A(G120gat), .B1(new_n338_), .B2(new_n342_), .ZN(new_n352_));
  OAI22_X1  g151(.A1(new_n349_), .A2(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n348_), .A2(new_n353_), .A3(KEYINPUT4), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n331_), .A2(new_n336_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n347_), .A2(new_n343_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n354_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT93), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT93), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n354_), .A2(new_n363_), .A3(new_n356_), .A4(new_n360_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n348_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT96), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n348_), .A2(new_n353_), .A3(KEYINPUT96), .A4(new_n355_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n362_), .A2(new_n364_), .A3(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT95), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G57gat), .B(G85gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n374_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n370_), .A2(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n362_), .A2(new_n369_), .A3(new_n377_), .A4(new_n364_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G228gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT21), .ZN(new_n384_));
  INV_X1    g183(.A(G204gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G197gat), .ZN(new_n386_));
  INV_X1    g185(.A(G197gat), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n387_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT85), .B1(new_n387_), .B2(G204gat), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n384_), .B(new_n386_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT86), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n387_), .A2(G204gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n387_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n384_), .A4(new_n386_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n384_), .B1(new_n392_), .B2(new_n386_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G211gat), .B(G218gat), .Z(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n391_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n396_), .A2(new_n386_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(KEYINPUT21), .A3(new_n400_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT87), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n383_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT29), .B1(new_n349_), .B2(new_n350_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(G233gat), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n409_), .B1(new_n407_), .B2(G233gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G78gat), .B(G106gat), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n413_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n402_), .A2(new_n404_), .ZN(new_n416_));
  OAI211_X1 g215(.A(G228gat), .B(G233gat), .C1(new_n416_), .C2(KEYINPUT87), .ZN(new_n417_));
  INV_X1    g216(.A(new_n409_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n415_), .B1(new_n419_), .B2(new_n410_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G22gat), .B(G50gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT28), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OR3_X1    g222(.A1(new_n357_), .A2(KEYINPUT29), .A3(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n423_), .B1(new_n357_), .B2(KEYINPUT29), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT88), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n414_), .A2(new_n420_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT88), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n424_), .A2(new_n429_), .A3(new_n425_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n413_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n419_), .A2(new_n410_), .A3(new_n415_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT80), .ZN(new_n435_));
  INV_X1    g234(.A(G169gat), .ZN(new_n436_));
  INV_X1    g235(.A(G176gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT24), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G183gat), .A2(G190gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT23), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT23), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(G183gat), .A3(G190gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n441_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT81), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n441_), .A2(KEYINPUT81), .A3(new_n446_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT26), .B(G190gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT79), .ZN(new_n453_));
  INV_X1    g252(.A(G183gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n453_), .B1(new_n454_), .B2(KEYINPUT25), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT25), .B(G183gat), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n452_), .B(new_n455_), .C1(new_n456_), .C2(new_n453_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n438_), .A2(new_n440_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n436_), .A2(new_n437_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(KEYINPUT24), .A3(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n451_), .A2(new_n457_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT82), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n445_), .A2(new_n463_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n444_), .A2(KEYINPUT82), .A3(G183gat), .A4(G190gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n443_), .A3(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(G183gat), .A2(G190gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT83), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n472_));
  AOI21_X1  g271(.A(G176gat), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(new_n459_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n466_), .A2(KEYINPUT83), .A3(new_n467_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n470_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n462_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G15gat), .B(G43gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT31), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n477_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G71gat), .B(G99gat), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n481_), .B1(new_n347_), .B2(new_n343_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n347_), .A2(new_n343_), .A3(new_n481_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n485_), .B(KEYINPUT30), .Z(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n483_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n487_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n480_), .B(new_n490_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n428_), .A2(new_n434_), .A3(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n488_), .A2(new_n489_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n480_), .B(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n427_), .A2(new_n430_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n414_), .B2(new_n420_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n432_), .A2(KEYINPUT88), .A3(new_n426_), .A4(new_n433_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n494_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n382_), .B1(new_n492_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n471_), .A2(new_n472_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n437_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(new_n460_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT90), .B1(new_n473_), .B2(new_n459_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n446_), .A2(new_n467_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n452_), .A2(new_n456_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n439_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n461_), .A2(new_n466_), .A3(new_n507_), .A4(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n405_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n416_), .A2(new_n462_), .A3(new_n476_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n405_), .A2(new_n510_), .A3(KEYINPUT91), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(KEYINPUT20), .A4(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G226gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT19), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n518_), .B(KEYINPUT89), .Z(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n462_), .A2(new_n476_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT20), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n405_), .A2(new_n510_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n518_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT18), .B(G64gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(G92gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G8gat), .B(G36gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  NAND3_X1  g330(.A1(new_n521_), .A2(new_n527_), .A3(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n516_), .A2(new_n520_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n525_), .A2(new_n526_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(KEYINPUT27), .B(new_n532_), .C1(new_n535_), .C2(new_n531_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n531_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n405_), .A2(KEYINPUT91), .A3(new_n510_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT91), .B1(new_n405_), .B2(new_n510_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n466_), .A2(KEYINPUT83), .A3(new_n467_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT83), .B1(new_n466_), .B2(new_n467_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n461_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n543_), .A2(new_n474_), .B1(new_n545_), .B2(new_n457_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n523_), .B1(new_n546_), .B2(new_n416_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n519_), .B1(new_n540_), .B2(new_n547_), .ZN(new_n548_));
  NOR4_X1   g347(.A1(new_n522_), .A2(new_n524_), .A3(new_n523_), .A4(new_n518_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n537_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT92), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n532_), .A3(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n548_), .A2(new_n549_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(KEYINPUT92), .A3(new_n531_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n536_), .B1(new_n555_), .B2(KEYINPUT27), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n499_), .A2(new_n556_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n354_), .A2(new_n355_), .A3(new_n360_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n348_), .A2(new_n353_), .ZN(new_n559_));
  AOI211_X1 g358(.A(new_n377_), .B(new_n558_), .C1(new_n356_), .C2(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n362_), .A2(new_n364_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT33), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(new_n377_), .A4(new_n369_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n380_), .A2(KEYINPUT33), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n560_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n555_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n555_), .A2(new_n565_), .A3(KEYINPUT97), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n531_), .A2(KEYINPUT32), .ZN(new_n570_));
  AOI22_X1  g369(.A1(new_n379_), .A2(new_n380_), .B1(new_n553_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT98), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n572_), .B1(new_n535_), .B2(new_n570_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n570_), .ZN(new_n574_));
  OAI211_X1 g373(.A(KEYINPUT98), .B(new_n574_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n571_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n568_), .A2(new_n569_), .A3(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n428_), .A2(new_n434_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(new_n491_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n557_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n316_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G57gat), .B(G64gat), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n583_), .A2(KEYINPUT11), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(KEYINPUT11), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586_));
  OR3_X1    g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(new_n586_), .A3(KEYINPUT11), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n582_), .B1(new_n271_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n589_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n237_), .A2(KEYINPUT12), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n271_), .A2(new_n589_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n590_), .A2(new_n592_), .A3(new_n593_), .A4(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n271_), .A2(new_n589_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n591_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n597_));
  OAI211_X1 g396(.A(G230gat), .B(G233gat), .C1(new_n596_), .C2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G120gat), .B(G148gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(new_n385_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT5), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n437_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n604_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n599_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT13), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(KEYINPUT69), .B2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G15gat), .B(G22gat), .ZN(new_n614_));
  INV_X1    g413(.A(G1gat), .ZN(new_n615_));
  INV_X1    g414(.A(G8gat), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT14), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G1gat), .B(G8gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n618_), .B(new_n619_), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n281_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G229gat), .A2(G233gat), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n273_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n620_), .B(new_n273_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(G229gat), .A3(G233gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G113gat), .B(G141gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(new_n436_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(new_n387_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n625_), .A2(new_n627_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n631_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n613_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT77), .Z(new_n639_));
  XNOR2_X1  g438(.A(new_n620_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(new_n591_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT17), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT16), .B(G183gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(G211gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G127gat), .B(G155gat), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n644_), .B(new_n645_), .Z(new_n646_));
  OAI21_X1  g445(.A(new_n641_), .B1(new_n642_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(KEYINPUT17), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n641_), .B2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT78), .Z(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n637_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n581_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n381_), .B(KEYINPUT99), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n615_), .A3(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT38), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n652_), .A2(KEYINPUT100), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n313_), .A2(new_n301_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n652_), .B2(KEYINPUT100), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n499_), .A2(new_n556_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n555_), .A2(new_n565_), .A3(KEYINPUT97), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT97), .B1(new_n555_), .B2(new_n565_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n571_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n579_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n660_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n657_), .A2(new_n659_), .A3(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(new_n381_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n656_), .B1(new_n615_), .B2(new_n668_), .ZN(G1324gat));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n556_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT101), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G8gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT39), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(new_n674_), .A3(G8gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n653_), .A2(new_n616_), .A3(new_n556_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n676_), .A2(KEYINPUT40), .A3(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1325gat));
  INV_X1    g481(.A(G15gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n667_), .B2(new_n491_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT41), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n653_), .A2(new_n683_), .A3(new_n491_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1326gat));
  INV_X1    g486(.A(G22gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n578_), .B(KEYINPUT102), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n667_), .B2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT42), .Z(new_n691_));
  NAND3_X1  g490(.A1(new_n653_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1327gat));
  INV_X1    g492(.A(new_n658_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n580_), .A2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n637_), .A2(new_n650_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT105), .Z(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n381_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n316_), .A2(new_n700_), .A3(new_n666_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n315_), .B1(new_n580_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n666_), .A2(KEYINPUT103), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT104), .B1(new_n705_), .B2(KEYINPUT43), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n707_));
  AOI211_X1 g506(.A(new_n707_), .B(new_n700_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n701_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n696_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n709_), .A2(KEYINPUT44), .A3(new_n696_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n712_), .A2(G29gat), .A3(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n699_), .B1(new_n714_), .B2(new_n654_), .ZN(G1328gat));
  INV_X1    g514(.A(new_n698_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n556_), .B(KEYINPUT106), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n716_), .A2(G36gat), .A3(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT45), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n712_), .A2(new_n556_), .A3(new_n713_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G36gat), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n720_), .A2(KEYINPUT46), .A3(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1329gat));
  NAND4_X1  g526(.A1(new_n712_), .A2(G43gat), .A3(new_n491_), .A4(new_n713_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n238_), .B1(new_n716_), .B2(new_n494_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g530(.A1(new_n712_), .A2(new_n578_), .A3(new_n713_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G50gat), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n689_), .A2(new_n242_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT107), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n698_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT108), .ZN(G1331gat));
  INV_X1    g537(.A(new_n613_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n581_), .A2(new_n635_), .A3(new_n739_), .A4(new_n650_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G57gat), .B1(new_n741_), .B2(new_n654_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n635_), .ZN(new_n743_));
  NOR4_X1   g542(.A1(new_n743_), .A2(new_n580_), .A3(new_n651_), .A4(new_n658_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(new_n381_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n742_), .B1(G57gat), .B2(new_n745_), .ZN(G1332gat));
  INV_X1    g545(.A(G64gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n744_), .B2(new_n717_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT48), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n741_), .A2(new_n747_), .A3(new_n717_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1333gat));
  INV_X1    g550(.A(G71gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n744_), .B2(new_n491_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT109), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT49), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n741_), .A2(new_n752_), .A3(new_n491_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT110), .Z(G1334gat));
  INV_X1    g557(.A(G78gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n744_), .B2(new_n689_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT50), .Z(new_n761_));
  NAND3_X1  g560(.A1(new_n741_), .A2(new_n759_), .A3(new_n689_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT111), .Z(G1335gat));
  NOR2_X1   g563(.A1(new_n743_), .A2(new_n650_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n695_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(G85gat), .B1(new_n767_), .B2(new_n654_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n709_), .A2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n765_), .B(KEYINPUT113), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT112), .B(new_n701_), .C1(new_n706_), .C2(new_n708_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT114), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n770_), .A2(new_n775_), .A3(new_n771_), .A4(new_n772_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n774_), .A2(new_n381_), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n768_), .B1(new_n777_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g577(.A(G92gat), .B1(new_n767_), .B2(new_n556_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n774_), .A2(G92gat), .A3(new_n776_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(new_n717_), .ZN(G1337gat));
  NAND3_X1  g580(.A1(new_n774_), .A2(new_n491_), .A3(new_n776_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(G99gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n767_), .A2(new_n203_), .A3(new_n491_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT51), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n783_), .A2(new_n787_), .A3(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1338gat));
  NAND3_X1  g588(.A1(new_n709_), .A2(new_n578_), .A3(new_n771_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G106gat), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(KEYINPUT115), .A3(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n767_), .A2(new_n204_), .A3(new_n578_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(KEYINPUT115), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n792_), .A2(KEYINPUT115), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n790_), .A2(G106gat), .A3(new_n795_), .A4(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n793_), .A2(new_n794_), .A3(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g598(.A(new_n654_), .ZN(new_n800_));
  NOR4_X1   g599(.A1(new_n800_), .A2(new_n556_), .A3(new_n578_), .A4(new_n494_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n626_), .A2(new_n623_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n622_), .A2(new_n624_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n804_), .B2(new_n623_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n632_), .B1(new_n805_), .B2(new_n631_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n608_), .A2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n635_), .A2(new_n607_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n595_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT117), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n595_), .A2(new_n810_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n590_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(G230gat), .A3(G233gat), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n595_), .A2(new_n816_), .A3(new_n810_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n812_), .A2(new_n813_), .A3(new_n815_), .A4(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n606_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n809_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n819_), .A2(new_n820_), .A3(KEYINPUT56), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n807_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT119), .B1(new_n825_), .B2(new_n658_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828_));
  INV_X1    g627(.A(new_n824_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT118), .B1(new_n818_), .B2(new_n606_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n808_), .B1(new_n830_), .B2(KEYINPUT56), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n828_), .B(new_n694_), .C1(new_n832_), .C2(new_n807_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n826_), .A2(new_n827_), .A3(new_n833_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n825_), .A2(new_n827_), .A3(new_n658_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n819_), .A2(KEYINPUT56), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n806_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n607_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n819_), .A2(KEYINPUT56), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n841_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n843_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .A4(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n316_), .A3(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n834_), .A2(new_n836_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT121), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n834_), .A2(new_n850_), .A3(new_n836_), .A4(new_n847_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(new_n651_), .A3(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n613_), .A2(new_n635_), .A3(new_n650_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT116), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n315_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT54), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n802_), .B1(new_n852_), .B2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(G113gat), .B1(new_n857_), .B2(new_n636_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n802_), .A2(KEYINPUT59), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n834_), .A2(new_n847_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n835_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n834_), .A2(KEYINPUT122), .A3(new_n847_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n650_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n856_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n859_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n857_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n635_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n858_), .B1(new_n869_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g669(.A(G120gat), .B1(new_n868_), .B2(new_n613_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n344_), .B1(new_n613_), .B2(KEYINPUT60), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n857_), .B(new_n872_), .C1(KEYINPUT60), .C2(new_n344_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(G1341gat));
  AOI21_X1  g673(.A(G127gat), .B1(new_n857_), .B2(new_n650_), .ZN(new_n875_));
  INV_X1    g674(.A(G127gat), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n868_), .A2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n877_), .B2(new_n650_), .ZN(G1342gat));
  NOR2_X1   g677(.A1(new_n694_), .A2(G134gat), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n857_), .A2(new_n879_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n866_), .B(new_n316_), .C1(new_n867_), .C2(new_n857_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(G134gat), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  AOI211_X1 g683(.A(KEYINPUT123), .B(new_n880_), .C1(new_n881_), .C2(G134gat), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1343gat));
  NAND2_X1  g685(.A1(new_n852_), .A2(new_n856_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n887_), .A2(new_n492_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n717_), .A2(new_n800_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n635_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT124), .B(G141gat), .Z(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1344gat));
  NOR2_X1   g692(.A1(new_n890_), .A2(new_n613_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(new_n321_), .ZN(G1345gat));
  NOR2_X1   g694(.A1(new_n890_), .A2(new_n651_), .ZN(new_n896_));
  XOR2_X1   g695(.A(KEYINPUT61), .B(G155gat), .Z(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1346gat));
  INV_X1    g697(.A(G162gat), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n890_), .A2(new_n899_), .A3(new_n315_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n888_), .A2(new_n658_), .A3(new_n889_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n899_), .B2(new_n901_), .ZN(G1347gat));
  OR2_X1    g701(.A1(new_n864_), .A2(new_n865_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n689_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n718_), .A2(new_n494_), .A3(new_n654_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(G169gat), .B1(new_n906_), .B2(new_n635_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n906_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n910_), .A2(new_n636_), .A3(new_n500_), .ZN(new_n911_));
  OAI211_X1 g710(.A(KEYINPUT62), .B(G169gat), .C1(new_n906_), .C2(new_n635_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n909_), .A2(new_n911_), .A3(new_n912_), .ZN(G1348gat));
  AOI21_X1  g712(.A(G176gat), .B1(new_n910_), .B2(new_n739_), .ZN(new_n914_));
  AND4_X1   g713(.A1(new_n498_), .A2(new_n887_), .A3(new_n800_), .A4(new_n717_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n613_), .A2(new_n437_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n915_), .B2(new_n916_), .ZN(G1349gat));
  NOR3_X1   g716(.A1(new_n906_), .A2(new_n651_), .A3(new_n456_), .ZN(new_n918_));
  AOI21_X1  g717(.A(G183gat), .B1(new_n915_), .B2(new_n650_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n906_), .B2(new_n315_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n658_), .A2(new_n452_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n906_), .B2(new_n922_), .ZN(G1351gat));
  AOI21_X1  g722(.A(new_n718_), .B1(new_n852_), .B2(new_n856_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n492_), .A2(new_n382_), .ZN(new_n925_));
  XOR2_X1   g724(.A(new_n925_), .B(KEYINPUT125), .Z(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n635_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT126), .B(G197gat), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1352gat));
  NOR2_X1   g729(.A1(new_n927_), .A2(new_n613_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(new_n385_), .ZN(G1353gat));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  AND2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  NOR4_X1   g733(.A1(new_n927_), .A2(new_n651_), .A3(new_n933_), .A4(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n927_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n650_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n935_), .B1(new_n937_), .B2(new_n933_), .ZN(G1354gat));
  XOR2_X1   g737(.A(KEYINPUT127), .B(G218gat), .Z(new_n939_));
  AND3_X1   g738(.A1(new_n936_), .A2(new_n316_), .A3(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n939_), .B1(new_n936_), .B2(new_n658_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1355gat));
endmodule


