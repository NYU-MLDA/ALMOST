//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203_));
  INV_X1    g002(.A(G50gat), .ZN(new_n204_));
  INV_X1    g003(.A(G29gat), .ZN(new_n205_));
  INV_X1    g004(.A(G36gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G43gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G29gat), .A2(G36gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n208_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n204_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT68), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n207_), .A2(new_n209_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(G43gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G50gat), .A3(new_n210_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n214_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n214_), .B1(new_n213_), .B2(new_n217_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n203_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G85gat), .ZN(new_n222_));
  INV_X1    g021(.A(G92gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT65), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT9), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT9), .ZN(new_n226_));
  OAI211_X1 g025(.A(KEYINPUT65), .B(new_n226_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n225_), .B(new_n227_), .C1(G85gat), .C2(G92gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT6), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT10), .B(G99gat), .Z(new_n233_));
  INV_X1    g032(.A(G106gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n228_), .A2(new_n231_), .A3(new_n232_), .A4(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT7), .ZN(new_n237_));
  INV_X1    g036(.A(G99gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(new_n234_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n239_), .A2(new_n231_), .A3(new_n232_), .A4(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G85gat), .B(G92gat), .Z(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(KEYINPUT8), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT8), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n245_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n236_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n211_), .A2(new_n204_), .A3(new_n212_), .ZN(new_n248_));
  AOI21_X1  g047(.A(G50gat), .B1(new_n216_), .B2(new_n210_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT68), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(KEYINPUT15), .A3(new_n218_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n221_), .A2(new_n247_), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n202_), .B1(new_n252_), .B2(KEYINPUT69), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G232gat), .A2(G233gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT34), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n243_), .B(KEYINPUT8), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n248_), .A2(new_n249_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n236_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n255_), .A2(KEYINPUT35), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n253_), .A2(new_n255_), .A3(new_n252_), .A4(new_n259_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT36), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G190gat), .B(G218gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(G134gat), .ZN(new_n267_));
  INV_X1    g066(.A(G162gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n264_), .A2(new_n265_), .A3(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(KEYINPUT36), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .A4(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT37), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n274_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n273_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(KEYINPUT66), .B(G71gat), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(G78gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT66), .B(G71gat), .ZN(new_n281_));
  INV_X1    g080(.A(G78gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G57gat), .B(G64gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT11), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n285_), .A2(KEYINPUT11), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n289_), .A2(new_n280_), .A3(new_n286_), .A4(new_n283_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G231gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G1gat), .B(G8gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT71), .ZN(new_n295_));
  INV_X1    g094(.A(G15gat), .ZN(new_n296_));
  INV_X1    g095(.A(G22gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G15gat), .A2(G22gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G1gat), .A2(G8gat), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n298_), .A2(new_n299_), .B1(KEYINPUT14), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n295_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n293_), .B(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G127gat), .B(G155gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT73), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT74), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G183gat), .B(G211gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n307_), .B(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT17), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n311_), .A2(new_n312_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n304_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(new_n314_), .B2(new_n304_), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(KEYINPUT75), .Z(new_n317_));
  NOR2_X1   g116(.A1(new_n278_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n291_), .B1(new_n257_), .B2(new_n236_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT12), .B1(new_n319_), .B2(KEYINPUT67), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G230gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT64), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n288_), .A2(new_n290_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n247_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT67), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT12), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n257_), .A2(new_n291_), .A3(new_n236_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n320_), .A2(new_n323_), .A3(new_n328_), .A4(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n325_), .A2(new_n329_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n330_), .B1(new_n323_), .B2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G120gat), .B(G148gat), .ZN(new_n333_));
  INV_X1    g132(.A(G204gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT5), .ZN(new_n336_));
  INV_X1    g135(.A(G176gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n332_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT13), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n318_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT76), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT85), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G141gat), .A2(G148gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT3), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n348_), .B1(KEYINPUT86), .B2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT86), .B(KEYINPUT3), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n350_), .B1(new_n351_), .B2(new_n348_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G141gat), .A2(G148gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT2), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n346_), .B(new_n347_), .C1(new_n352_), .C2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n348_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n344_), .B(KEYINPUT85), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n347_), .B(KEYINPUT1), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n357_), .B(new_n353_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT29), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT88), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(new_n334_), .A3(G197gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n364_), .B1(G197gat), .B2(new_n334_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(G197gat), .B2(new_n334_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT21), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G211gat), .B(G218gat), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OR3_X1    g168(.A1(new_n334_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n370_));
  INV_X1    g169(.A(G197gat), .ZN(new_n371_));
  OR3_X1    g170(.A1(new_n371_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT90), .B1(new_n334_), .B2(G197gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT89), .B1(new_n371_), .B2(G204gat), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n370_), .A2(new_n372_), .A3(new_n373_), .A4(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n367_), .B(new_n369_), .C1(new_n375_), .C2(KEYINPUT21), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(KEYINPUT21), .A3(new_n368_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n362_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(G228gat), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n379_), .B(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G78gat), .B(G106gat), .Z(new_n385_));
  XOR2_X1   g184(.A(new_n384_), .B(new_n385_), .Z(new_n386_));
  NOR2_X1   g185(.A1(new_n361_), .A2(KEYINPUT29), .ZN(new_n387_));
  XOR2_X1   g186(.A(G22gat), .B(G50gat), .Z(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT28), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n387_), .B(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n384_), .A2(new_n385_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n391_), .B2(KEYINPUT91), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n386_), .B(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G8gat), .B(G36gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n378_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT24), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT94), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT94), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT24), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G169gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n337_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G183gat), .A2(G190gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT23), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n417_), .A2(new_n418_), .A3(KEYINPUT93), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT93), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT26), .ZN(new_n421_));
  INV_X1    g220(.A(G190gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n420_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n416_), .B1(new_n419_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G169gat), .A2(G176gat), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n406_), .A2(new_n401_), .A3(new_n403_), .A4(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT95), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT93), .B1(new_n417_), .B2(new_n418_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n423_), .A2(new_n420_), .A3(new_n424_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n415_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT95), .ZN(new_n433_));
  INV_X1    g232(.A(new_n428_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n412_), .B1(new_n429_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n410_), .B1(G183gat), .B2(G190gat), .ZN(new_n437_));
  XOR2_X1   g236(.A(KEYINPUT80), .B(G176gat), .Z(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT22), .B(G169gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n437_), .A2(new_n427_), .A3(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n399_), .A2(new_n436_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G226gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT19), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT81), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n440_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n438_), .A2(KEYINPUT81), .A3(new_n439_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n448_), .A2(new_n437_), .A3(new_n427_), .A4(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n416_), .B1(new_n418_), .B2(new_n417_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n407_), .A2(new_n400_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n406_), .A2(KEYINPUT24), .A3(new_n427_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n451_), .A2(new_n410_), .A3(new_n452_), .A4(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n446_), .B1(new_n455_), .B2(new_n378_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n442_), .A2(new_n445_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n436_), .A2(new_n441_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n378_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n455_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n446_), .B1(new_n460_), .B2(new_n399_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n444_), .B(KEYINPUT92), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n398_), .B(new_n457_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n436_), .A2(KEYINPUT101), .A3(new_n441_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT101), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n426_), .A2(KEYINPUT95), .A3(new_n428_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n433_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n411_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n441_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n466_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n465_), .A2(new_n471_), .A3(new_n399_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n456_), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT102), .B1(new_n473_), .B2(new_n444_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT102), .ZN(new_n475_));
  AOI211_X1 g274(.A(new_n475_), .B(new_n445_), .C1(new_n472_), .C2(new_n456_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n459_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n474_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  OAI211_X1 g277(.A(KEYINPUT27), .B(new_n464_), .C1(new_n478_), .C2(new_n398_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n398_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n463_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n457_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n464_), .A2(new_n483_), .A3(KEYINPUT97), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT97), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n485_), .B(new_n480_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT103), .B(KEYINPUT27), .Z(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n479_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G225gat), .A2(G233gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G127gat), .B(G134gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G113gat), .B(G120gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(KEYINPUT82), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n491_), .B(new_n492_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n493_), .B1(new_n494_), .B2(KEYINPUT82), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n495_), .A2(new_n361_), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n496_), .A2(KEYINPUT4), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n356_), .A2(new_n494_), .A3(new_n360_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT4), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n490_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n496_), .A2(new_n498_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n490_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G1gat), .B(G29gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G57gat), .B(G85gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(KEYINPUT98), .B(KEYINPUT0), .Z(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  OR3_X1    g307(.A1(new_n500_), .A2(new_n503_), .A3(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n508_), .B1(new_n500_), .B2(new_n503_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n393_), .B1(new_n489_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n473_), .A2(new_n444_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n475_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n477_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n473_), .A2(KEYINPUT102), .A3(new_n444_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n398_), .A2(KEYINPUT32), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NOR3_X1   g320(.A1(new_n481_), .A2(new_n482_), .A3(new_n520_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT100), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n523_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n521_), .A2(new_n511_), .A3(new_n524_), .A4(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n484_), .A2(new_n486_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n501_), .A2(new_n490_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n497_), .A2(new_n499_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n528_), .B(new_n508_), .C1(new_n529_), .C2(new_n502_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT99), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT33), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n509_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n500_), .A2(new_n503_), .A3(new_n508_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT33), .B1(new_n534_), .B2(KEYINPUT99), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n527_), .A2(new_n530_), .A3(new_n533_), .A4(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n526_), .A2(new_n393_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n455_), .A2(KEYINPUT30), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n455_), .A2(KEYINPUT30), .ZN(new_n540_));
  OAI21_X1  g339(.A(G43gat), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n455_), .A2(KEYINPUT30), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n542_), .A2(new_n208_), .A3(new_n538_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G227gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(G15gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G71gat), .B(G99gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  AND3_X1   g346(.A1(new_n541_), .A2(new_n543_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n547_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT31), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n550_), .A2(KEYINPUT83), .B1(new_n551_), .B2(new_n495_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n495_), .A2(new_n551_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT83), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT84), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n541_), .A2(new_n543_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n547_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n541_), .A2(new_n543_), .A3(new_n547_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT84), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n554_), .A3(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n552_), .A2(new_n553_), .A3(new_n556_), .A4(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n495_), .A2(new_n551_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n553_), .B(new_n565_), .C1(new_n561_), .C2(new_n554_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n562_), .B1(new_n561_), .B2(new_n554_), .ZN(new_n567_));
  AOI211_X1 g366(.A(KEYINPUT83), .B(KEYINPUT84), .C1(new_n559_), .C2(new_n560_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n537_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n513_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n393_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT27), .ZN(new_n575_));
  INV_X1    g374(.A(new_n464_), .ZN(new_n576_));
  AOI211_X1 g375(.A(new_n575_), .B(new_n576_), .C1(new_n518_), .C2(new_n480_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n488_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT104), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT104), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n479_), .A2(new_n580_), .A3(new_n488_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n574_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n511_), .B1(new_n564_), .B2(new_n569_), .ZN(new_n583_));
  AOI21_X1  g382(.A(KEYINPUT105), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n479_), .A2(new_n580_), .A3(new_n488_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n580_), .B1(new_n479_), .B2(new_n488_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n393_), .B(new_n583_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT105), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n573_), .B1(new_n584_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT106), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT77), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n302_), .A2(new_n258_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n302_), .A2(new_n258_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n592_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n595_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(KEYINPUT77), .A3(new_n593_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n596_), .A2(new_n598_), .A3(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n221_), .A2(new_n303_), .A3(new_n251_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n599_), .A3(new_n593_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT78), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT78), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n602_), .A2(new_n605_), .A3(new_n599_), .A4(new_n593_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n601_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G113gat), .B(G141gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(new_n405_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(new_n371_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n607_), .A2(KEYINPUT79), .A3(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n607_), .B2(KEYINPUT79), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n590_), .A2(new_n591_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n587_), .A2(new_n588_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n579_), .A2(new_n581_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n617_), .A2(KEYINPUT105), .A3(new_n393_), .A4(new_n583_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n572_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT106), .B1(new_n619_), .B2(new_n613_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n343_), .B1(new_n615_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(G1gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n622_), .A3(new_n511_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT38), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n624_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT109), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n270_), .A2(KEYINPUT108), .A3(new_n272_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT108), .B1(new_n270_), .B2(new_n272_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n590_), .A2(new_n627_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT108), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n273_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n270_), .A2(KEYINPUT108), .A3(new_n272_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT109), .B1(new_n619_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n340_), .A2(new_n613_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n317_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT107), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n637_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n642_), .A2(new_n511_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n625_), .B(new_n626_), .C1(new_n622_), .C2(new_n643_), .ZN(G1324gat));
  INV_X1    g443(.A(G8gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n617_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n621_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n637_), .A2(new_n646_), .A3(new_n641_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n648_), .A2(new_n649_), .A3(G8gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n648_), .B2(G8gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n647_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(G1325gat));
  INV_X1    g453(.A(new_n570_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n621_), .A2(new_n296_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n642_), .A2(new_n655_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT41), .B1(new_n657_), .B2(G15gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n656_), .B1(new_n658_), .B2(new_n659_), .ZN(G1326gat));
  NAND3_X1  g459(.A1(new_n621_), .A2(new_n297_), .A3(new_n574_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n642_), .A2(new_n574_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G22gat), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n663_), .A2(KEYINPUT42), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(KEYINPUT42), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(G1327gat));
  NAND2_X1  g465(.A1(KEYINPUT112), .A2(KEYINPUT44), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT43), .B1(new_n277_), .B2(KEYINPUT111), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n590_), .A2(new_n278_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n668_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n670_), .B1(new_n619_), .B2(new_n277_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  OR2_X1    g471(.A1(KEYINPUT112), .A2(KEYINPUT44), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n638_), .A2(new_n317_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT110), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AND4_X1   g475(.A1(new_n667_), .A2(new_n672_), .A3(new_n673_), .A4(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n675_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n667_), .B1(new_n678_), .B2(new_n673_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n512_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n340_), .B1(new_n615_), .B2(new_n620_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n639_), .A2(new_n630_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n205_), .A3(new_n511_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n681_), .A2(new_n685_), .ZN(G1328gat));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n682_), .A2(new_n206_), .A3(new_n646_), .A4(new_n683_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT45), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n668_), .B1(new_n590_), .B2(new_n278_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n619_), .A2(new_n277_), .A3(new_n670_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n676_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(KEYINPUT112), .A3(KEYINPUT44), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n678_), .A2(new_n667_), .A3(new_n673_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n206_), .B1(new_n696_), .B2(new_n646_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n687_), .B1(new_n690_), .B2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G36gat), .B1(new_n680_), .B2(new_n617_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n688_), .B(KEYINPUT45), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(KEYINPUT46), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(G1329gat));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n655_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G43gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n684_), .A2(new_n208_), .A3(new_n655_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n703_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n570_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n703_), .B(new_n706_), .C1(new_n708_), .C2(new_n208_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n707_), .A2(new_n710_), .ZN(G1330gat));
  OAI21_X1  g510(.A(G50gat), .B1(new_n680_), .B2(new_n393_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n684_), .A2(new_n204_), .A3(new_n574_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1331gat));
  NOR2_X1   g513(.A1(new_n341_), .A2(new_n614_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n619_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n318_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(G57gat), .B1(new_n719_), .B2(new_n511_), .ZN(new_n720_));
  AOI211_X1 g519(.A(new_n317_), .B(new_n716_), .C1(new_n631_), .C2(new_n636_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(new_n511_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n722_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g522(.A(G64gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(new_n724_), .A3(new_n646_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n721_), .A2(new_n646_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G64gat), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT48), .B(new_n724_), .C1(new_n721_), .C2(new_n646_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1333gat));
  OR3_X1    g529(.A1(new_n718_), .A2(G71gat), .A3(new_n570_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n637_), .A2(new_n655_), .A3(new_n639_), .A4(new_n715_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G71gat), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT113), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(new_n735_), .A3(G71gat), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n734_), .A2(KEYINPUT49), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT49), .B1(new_n734_), .B2(new_n736_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n731_), .B1(new_n737_), .B2(new_n738_), .ZN(G1334gat));
  NAND3_X1  g538(.A1(new_n719_), .A2(new_n282_), .A3(new_n574_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n721_), .A2(new_n574_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(G78gat), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT50), .B(new_n282_), .C1(new_n721_), .C2(new_n574_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1335gat));
  AND2_X1   g544(.A1(new_n717_), .A2(new_n683_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G85gat), .B1(new_n746_), .B2(new_n511_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT114), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n639_), .B(new_n716_), .C1(new_n669_), .C2(new_n671_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n749_), .A2(G85gat), .A3(new_n511_), .ZN(new_n750_));
  OR3_X1    g549(.A1(new_n748_), .A2(KEYINPUT115), .A3(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT115), .B1(new_n748_), .B2(new_n750_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1336gat));
  AOI21_X1  g552(.A(G92gat), .B1(new_n746_), .B2(new_n646_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n749_), .A2(G92gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(new_n646_), .ZN(G1337gat));
  NAND3_X1  g555(.A1(new_n746_), .A2(new_n233_), .A3(new_n655_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT116), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n749_), .A2(new_n655_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(G99gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT117), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(KEYINPUT51), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT51), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n758_), .A2(new_n764_), .A3(new_n760_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n746_), .A2(new_n234_), .A3(new_n574_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n672_), .A2(new_n574_), .A3(new_n317_), .A4(new_n715_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(G106gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G106gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g572(.A(G113gat), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n582_), .A2(new_n511_), .A3(new_n655_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n277_), .A2(new_n341_), .A3(new_n613_), .A4(new_n639_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT54), .Z(new_n777_));
  INV_X1    g576(.A(KEYINPUT56), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n330_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n330_), .B2(new_n779_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n320_), .A2(new_n329_), .A3(new_n328_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(new_n322_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n781_), .A2(new_n782_), .A3(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n778_), .B1(new_n785_), .B2(new_n338_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n787_));
  INV_X1    g586(.A(new_n338_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n330_), .A2(new_n779_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT55), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n330_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT56), .B(new_n788_), .C1(new_n792_), .C2(new_n784_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n786_), .A2(new_n787_), .A3(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT119), .B(new_n778_), .C1(new_n785_), .C2(new_n338_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n600_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n599_), .B1(new_n602_), .B2(new_n593_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n610_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n607_), .B2(new_n610_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n332_), .A2(new_n788_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n794_), .A2(new_n795_), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT120), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT58), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT58), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n802_), .A2(new_n803_), .A3(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n278_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n339_), .A2(new_n799_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n786_), .A2(new_n793_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n612_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n607_), .A2(KEYINPUT79), .A3(new_n610_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n800_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n810_), .B1(new_n811_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n809_), .B1(new_n815_), .B2(new_n635_), .ZN(new_n816_));
  OAI22_X1  g615(.A1(new_n611_), .A2(new_n612_), .B1(new_n332_), .B2(new_n788_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(new_n786_), .B2(new_n793_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n630_), .B(KEYINPUT57), .C1(new_n818_), .C2(new_n810_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n816_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n639_), .B1(new_n808_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n775_), .B1(new_n777_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n774_), .B1(new_n822_), .B2(new_n613_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT121), .ZN(new_n824_));
  INV_X1    g623(.A(new_n777_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n808_), .A2(new_n820_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT122), .B1(new_n826_), .B2(new_n317_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n828_), .B(new_n639_), .C1(new_n808_), .C2(new_n820_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n825_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n775_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n822_), .A2(KEYINPUT59), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n832_), .A2(KEYINPUT123), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT123), .B1(new_n832_), .B2(new_n833_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n613_), .A2(new_n774_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n824_), .B1(new_n836_), .B2(new_n837_), .ZN(G1340gat));
  INV_X1    g637(.A(new_n822_), .ZN(new_n839_));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n341_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT124), .B1(new_n840_), .B2(KEYINPUT60), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n839_), .B(new_n843_), .C1(new_n844_), .C2(new_n841_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n832_), .A2(new_n340_), .A3(new_n833_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n840_), .ZN(G1341gat));
  AOI21_X1  g646(.A(G127gat), .B1(new_n839_), .B2(new_n639_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(KEYINPUT125), .A2(G127gat), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n834_), .A2(new_n835_), .A3(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G127gat), .B1(new_n317_), .B2(KEYINPUT125), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n848_), .B1(new_n850_), .B2(new_n851_), .ZN(G1342gat));
  AOI21_X1  g651(.A(G134gat), .B1(new_n839_), .B2(new_n635_), .ZN(new_n853_));
  INV_X1    g652(.A(G134gat), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n834_), .A2(new_n835_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n855_), .B2(new_n278_), .ZN(G1343gat));
  OAI211_X1 g655(.A(new_n574_), .B(new_n570_), .C1(new_n777_), .C2(new_n821_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n646_), .A2(new_n512_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n614_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n340_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g663(.A1(new_n860_), .A2(new_n639_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT61), .B(G155gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  AOI21_X1  g666(.A(G162gat), .B1(new_n860_), .B2(new_n635_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n857_), .A2(new_n268_), .A3(new_n859_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n278_), .B2(new_n869_), .ZN(G1347gat));
  AND2_X1   g669(.A1(new_n830_), .A2(new_n393_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n617_), .A2(new_n511_), .A3(new_n570_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n614_), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G169gat), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n871_), .A2(new_n439_), .A3(new_n614_), .A4(new_n872_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n873_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n877_), .A3(new_n878_), .ZN(G1348gat));
  NAND3_X1  g678(.A1(new_n871_), .A2(new_n340_), .A3(new_n872_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n777_), .A2(new_n821_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n574_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n872_), .A2(G176gat), .A3(new_n340_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n880_), .A2(new_n438_), .B1(new_n882_), .B2(new_n883_), .ZN(G1349gat));
  NAND2_X1  g683(.A1(new_n872_), .A2(new_n639_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G183gat), .B1(new_n882_), .B2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n416_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n871_), .B2(new_n888_), .ZN(G1350gat));
  NAND2_X1  g688(.A1(new_n430_), .A2(new_n431_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n871_), .A2(new_n635_), .A3(new_n890_), .A4(new_n872_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n871_), .A2(new_n278_), .A3(new_n872_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n422_), .ZN(G1351gat));
  NOR3_X1   g692(.A1(new_n857_), .A2(new_n511_), .A3(new_n617_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n614_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n340_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT126), .B(G204gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1353gat));
  NAND2_X1  g698(.A1(new_n894_), .A2(new_n639_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  AND2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n900_), .B2(new_n901_), .ZN(G1354gat));
  INV_X1    g703(.A(KEYINPUT127), .ZN(new_n905_));
  INV_X1    g704(.A(new_n894_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n630_), .ZN(new_n907_));
  INV_X1    g706(.A(G218gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n894_), .A2(KEYINPUT127), .A3(new_n635_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n894_), .A2(G218gat), .A3(new_n278_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1355gat));
endmodule


