//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT10), .B(G99gat), .Z(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  AND3_X1   g004(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G85gat), .ZN(new_n210_));
  INV_X1    g009(.A(G92gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(KEYINPUT9), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(KEYINPUT9), .B2(new_n213_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n209_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G85gat), .B(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT64), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n212_), .A2(new_n219_), .A3(new_n213_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT7), .ZN(new_n222_));
  INV_X1    g021(.A(G99gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n204_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n208_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n225_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n221_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT8), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n208_), .A2(new_n226_), .A3(new_n224_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n221_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n216_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G57gat), .B(G64gat), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n238_));
  XOR2_X1   g037(.A(G71gat), .B(G78gat), .Z(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n238_), .A2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT68), .B1(new_n235_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT12), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G230gat), .A2(G233gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT12), .ZN(new_n246_));
  OAI211_X1 g045(.A(KEYINPUT68), .B(new_n246_), .C1(new_n235_), .C2(new_n242_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n235_), .A2(new_n242_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n244_), .A2(new_n245_), .A3(new_n247_), .A4(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n243_), .A2(KEYINPUT12), .B1(new_n242_), .B2(new_n235_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n252_), .A2(KEYINPUT69), .A3(new_n245_), .A4(new_n247_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n245_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n209_), .A2(new_n215_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n224_), .A2(new_n226_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT65), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(new_n208_), .A3(new_n227_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n232_), .B1(new_n259_), .B2(new_n221_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n221_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n256_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n263_));
  INV_X1    g062(.A(new_n242_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n248_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n263_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n267_));
  OAI211_X1 g066(.A(KEYINPUT67), .B(new_n255_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT66), .B1(new_n235_), .B2(new_n242_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(new_n248_), .A3(new_n265_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT67), .B1(new_n271_), .B2(new_n255_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G120gat), .B(G148gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(G204gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT5), .B(G176gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n275_), .B(new_n276_), .Z(new_n277_));
  NAND3_X1  g076(.A1(new_n254_), .A2(new_n273_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n277_), .B1(new_n254_), .B2(new_n273_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n202_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n254_), .A2(new_n273_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n277_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(KEYINPUT70), .A3(new_n278_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT13), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n281_), .A2(new_n285_), .A3(KEYINPUT13), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G29gat), .B(G36gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G43gat), .B(G50gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G15gat), .B(G22gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G1gat), .A2(G8gat), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n296_), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT74), .B1(new_n296_), .B2(KEYINPUT14), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n295_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(KEYINPUT75), .ZN(new_n300_));
  XOR2_X1   g099(.A(G1gat), .B(G8gat), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(KEYINPUT75), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n301_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n294_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n305_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(new_n303_), .A3(new_n293_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n308_), .A3(KEYINPUT79), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT79), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n310_), .B(new_n294_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n309_), .A2(G229gat), .A3(new_n311_), .A4(G233gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n304_), .A2(new_n305_), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n293_), .B(KEYINPUT15), .Z(new_n314_));
  OR2_X1    g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G229gat), .A2(G233gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(new_n316_), .A3(new_n308_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G169gat), .B(G197gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(G113gat), .B(G141gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT80), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n312_), .A2(new_n317_), .A3(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(new_n312_), .B2(new_n317_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n290_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(KEYINPUT82), .B(G176gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT22), .B(G169gat), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT23), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(G183gat), .A3(G190gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT23), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT83), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n335_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT81), .B(G183gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n342_), .A2(G190gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n332_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n337_), .A2(new_n334_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(G169gat), .B2(G176gat), .ZN(new_n348_));
  INV_X1    g147(.A(G169gat), .ZN(new_n349_));
  INV_X1    g148(.A(G176gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n346_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n353_), .B1(new_n342_), .B2(KEYINPUT25), .ZN(new_n354_));
  INV_X1    g153(.A(G190gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT26), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT26), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G190gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n345_), .B(new_n352_), .C1(new_n354_), .C2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n344_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT31), .B(G43gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G113gat), .B(G120gat), .Z(new_n366_));
  INV_X1    g165(.A(KEYINPUT84), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G113gat), .B(G120gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT84), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G127gat), .B(G134gat), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n368_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G71gat), .B(G99gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT30), .B(G15gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n374_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n365_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT85), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(G92gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT18), .B(G64gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G197gat), .B(G204gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT21), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G211gat), .B(G218gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n386_), .A2(new_n387_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n389_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n391_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n361_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT20), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n348_), .A2(new_n351_), .ZN(new_n400_));
  AND2_X1   g199(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n356_), .B(new_n358_), .C1(new_n401_), .C2(new_n353_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n346_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n405_));
  NOR2_X1   g204(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT82), .B(G176gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n328_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(G183gat), .A2(G190gat), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n337_), .B2(new_n334_), .ZN(new_n411_));
  OAI22_X1  g210(.A1(new_n404_), .A2(new_n341_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n395_), .B(new_n399_), .C1(new_n394_), .C2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT20), .B1(new_n361_), .B2(new_n394_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n412_), .A2(new_n394_), .A3(KEYINPUT94), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT94), .B1(new_n412_), .B2(new_n394_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n397_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n385_), .B(new_n413_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT27), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n344_), .A2(new_n360_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n394_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT20), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n392_), .A2(new_n393_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT92), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(new_n425_), .A3(new_n391_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n394_), .A2(KEYINPUT92), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n412_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n397_), .B1(new_n423_), .B2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n398_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n412_), .A2(new_n394_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT94), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n412_), .A2(new_n394_), .A3(KEYINPUT94), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n430_), .A2(new_n418_), .A3(new_n433_), .A4(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n385_), .B1(new_n429_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT99), .B1(new_n420_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT27), .ZN(new_n438_));
  INV_X1    g237(.A(new_n419_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n433_), .A2(new_n434_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n397_), .B1(new_n440_), .B2(new_n414_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n385_), .B1(new_n441_), .B2(new_n413_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n438_), .B1(new_n439_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n429_), .A2(new_n435_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n384_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT99), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(KEYINPUT27), .A4(new_n419_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n437_), .A2(new_n443_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT93), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n450_), .B1(G155gat), .B2(G162gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G155gat), .A2(G162gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n452_), .A2(KEYINPUT87), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT1), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(G155gat), .A2(G162gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(KEYINPUT88), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT1), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n452_), .A2(KEYINPUT87), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n450_), .A2(G155gat), .A3(G162gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n458_), .B1(new_n462_), .B2(new_n455_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n460_), .A2(new_n461_), .A3(new_n459_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n457_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(G141gat), .A2(G148gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G141gat), .A2(G148gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n466_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n455_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n466_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n476_));
  OAI22_X1  g275(.A1(KEYINPUT89), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .A4(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT2), .B1(new_n469_), .B2(new_n470_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n472_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT90), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n482_), .B(new_n472_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n465_), .A2(new_n471_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT29), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n426_), .A2(new_n427_), .ZN(new_n487_));
  OAI211_X1 g286(.A(G228gat), .B(G233gat), .C1(new_n486_), .C2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n465_), .A2(new_n471_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n481_), .A2(new_n483_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n484_), .A2(KEYINPUT91), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n485_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(G228gat), .ZN(new_n496_));
  INV_X1    g295(.A(G233gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n394_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n488_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G78gat), .B(G106gat), .Z(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n449_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT91), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT91), .B1(new_n489_), .B2(new_n490_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n485_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G22gat), .B(G50gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT28), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n506_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n498_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n511_), .B1(new_n505_), .B2(new_n485_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(new_n500_), .A3(new_n488_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n500_), .B1(new_n512_), .B2(new_n488_), .ZN(new_n515_));
  OAI22_X1  g314(.A1(new_n502_), .A2(new_n510_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n506_), .B(new_n508_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n499_), .A2(new_n501_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n517_), .A2(new_n449_), .A3(new_n513_), .A4(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n448_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT98), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G225gat), .A2(G233gat), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n374_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT95), .ZN(new_n524_));
  INV_X1    g323(.A(new_n374_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n524_), .B1(new_n491_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n484_), .A2(KEYINPUT95), .A3(new_n374_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT4), .B1(new_n523_), .B2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n525_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT4), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n522_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G1gat), .B(G29gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(new_n210_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT0), .B(G57gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  INV_X1    g336(.A(new_n522_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n523_), .A2(new_n528_), .A3(new_n538_), .ZN(new_n539_));
  NOR3_X1   g338(.A1(new_n533_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n537_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT95), .B1(new_n484_), .B2(new_n374_), .ZN(new_n542_));
  AND4_X1   g341(.A1(KEYINPUT95), .A2(new_n489_), .A3(new_n490_), .A4(new_n374_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n531_), .B1(new_n544_), .B2(new_n530_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n523_), .A2(KEYINPUT4), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n538_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n539_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n541_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n521_), .B1(new_n540_), .B2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n537_), .B1(new_n533_), .B2(new_n539_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n541_), .A3(new_n548_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(KEYINPUT98), .A3(new_n552_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n520_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n516_), .A2(new_n519_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT96), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(KEYINPUT33), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n557_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n547_), .A2(new_n541_), .A3(new_n548_), .A4(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n442_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n419_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n522_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n523_), .A2(new_n528_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n541_), .B1(new_n564_), .B2(new_n538_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n562_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n558_), .A2(new_n560_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n385_), .A2(KEYINPUT32), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n441_), .A2(new_n568_), .A3(new_n413_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n429_), .B2(new_n435_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT97), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n569_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n571_), .B2(new_n570_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n573_), .B1(new_n540_), .B2(new_n549_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n555_), .B1(new_n567_), .B2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n380_), .B1(new_n554_), .B2(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n550_), .A2(new_n553_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n516_), .A2(new_n519_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n448_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(KEYINPUT100), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT100), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(new_n555_), .B2(new_n448_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n577_), .A2(new_n580_), .A3(new_n379_), .A4(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n576_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(G231gat), .B(G233gat), .C1(new_n304_), .C2(new_n305_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n307_), .A2(new_n586_), .A3(new_n303_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n242_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n585_), .A2(new_n264_), .A3(new_n587_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G127gat), .B(G155gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(G211gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT16), .B(G183gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n594_), .A2(KEYINPUT17), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(KEYINPUT17), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n589_), .A2(new_n590_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT77), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n589_), .A2(new_n590_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n602_), .A2(KEYINPUT76), .A3(new_n595_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT76), .B1(new_n602_), .B2(new_n595_), .ZN(new_n604_));
  OAI22_X1  g403(.A1(new_n600_), .A2(new_n601_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT78), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OAI221_X1 g406(.A(KEYINPUT78), .B1(new_n603_), .B2(new_n604_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT34), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT35), .Z(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n314_), .A2(new_n262_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n235_), .A2(new_n294_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n613_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n614_), .A2(new_n615_), .A3(KEYINPUT35), .A4(new_n611_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n617_), .A2(KEYINPUT71), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(KEYINPUT71), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n616_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(G162gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT72), .B(G134gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(KEYINPUT36), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n624_), .B(KEYINPUT36), .Z(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(new_n620_), .B2(KEYINPUT73), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT73), .ZN(new_n629_));
  AOI211_X1 g428(.A(new_n629_), .B(new_n616_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT37), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n627_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n626_), .B(KEYINPUT37), .C1(new_n620_), .C2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n327_), .A2(new_n584_), .A3(new_n609_), .A4(new_n637_), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n638_), .A2(G1gat), .A3(new_n577_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT38), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT102), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n327_), .A2(new_n584_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n631_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(new_n605_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT101), .ZN(new_n647_));
  INV_X1    g446(.A(new_n577_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(G1gat), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n642_), .B(new_n650_), .C1(new_n640_), .C2(new_n639_), .ZN(G1324gat));
  OR3_X1    g450(.A1(new_n638_), .A2(G8gat), .A3(new_n579_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n327_), .A2(new_n584_), .A3(new_n448_), .A4(new_n645_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n654_), .B2(G8gat), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT103), .Z(new_n656_));
  NAND3_X1  g455(.A1(new_n654_), .A2(new_n653_), .A3(G8gat), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT104), .Z(new_n658_));
  OAI21_X1  g457(.A(new_n652_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1325gat));
  INV_X1    g460(.A(new_n380_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n647_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G15gat), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT41), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(KEYINPUT41), .ZN(new_n666_));
  OR3_X1    g465(.A1(new_n638_), .A2(G15gat), .A3(new_n380_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n665_), .A2(new_n666_), .A3(new_n667_), .ZN(G1326gat));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n647_), .A2(new_n555_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(G22gat), .ZN(new_n671_));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT42), .B(new_n672_), .C1(new_n647_), .C2(new_n555_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n555_), .A2(new_n672_), .ZN(new_n674_));
  OAI22_X1  g473(.A1(new_n671_), .A2(new_n673_), .B1(new_n638_), .B2(new_n674_), .ZN(G1327gat));
  NOR3_X1   g474(.A1(new_n290_), .A2(new_n609_), .A3(new_n326_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n584_), .B2(new_n636_), .ZN(new_n678_));
  AOI211_X1 g477(.A(KEYINPUT43), .B(new_n637_), .C1(new_n576_), .C2(new_n583_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n676_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT44), .B(new_n676_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n577_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n609_), .A2(new_n631_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n643_), .A2(new_n686_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n577_), .A2(G29gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n685_), .B1(new_n687_), .B2(new_n688_), .ZN(G1328gat));
  NAND3_X1  g488(.A1(new_n682_), .A2(new_n448_), .A3(new_n683_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT105), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n682_), .A2(new_n692_), .A3(new_n448_), .A4(new_n683_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(G36gat), .A3(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n579_), .A2(G36gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n643_), .A2(new_n686_), .A3(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT106), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n643_), .A2(new_n698_), .A3(new_n686_), .A4(new_n695_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n697_), .A2(KEYINPUT45), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT45), .B1(new_n697_), .B2(new_n699_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n694_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n694_), .A2(KEYINPUT46), .A3(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  NOR3_X1   g506(.A1(new_n687_), .A2(G43gat), .A3(new_n380_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n682_), .A2(new_n379_), .A3(new_n683_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(G43gat), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n710_), .B(new_n711_), .Z(G1330gat));
  OAI21_X1  g511(.A(G50gat), .B1(new_n684_), .B2(new_n578_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n578_), .A2(G50gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n687_), .B2(new_n714_), .ZN(G1331gat));
  AND3_X1   g514(.A1(new_n584_), .A2(new_n326_), .A3(new_n290_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n609_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n637_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT108), .ZN(new_n720_));
  OR3_X1    g519(.A1(new_n717_), .A2(KEYINPUT108), .A3(new_n636_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n648_), .A3(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(G57gat), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n722_), .A2(KEYINPUT109), .A3(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT109), .B1(new_n722_), .B2(new_n723_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n717_), .A2(new_n644_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n727_), .A2(new_n723_), .A3(new_n577_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n724_), .A2(new_n725_), .A3(new_n728_), .ZN(G1332gat));
  INV_X1    g528(.A(G64gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n726_), .B2(new_n448_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n731_), .A2(new_n732_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n448_), .A2(new_n730_), .ZN(new_n736_));
  OAI22_X1  g535(.A1(new_n734_), .A2(new_n735_), .B1(new_n719_), .B2(new_n736_), .ZN(G1333gat));
  OAI21_X1  g536(.A(G71gat), .B1(new_n727_), .B2(new_n380_), .ZN(new_n738_));
  XOR2_X1   g537(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n739_));
  OR2_X1    g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n739_), .ZN(new_n741_));
  OR3_X1    g540(.A1(new_n719_), .A2(G71gat), .A3(new_n380_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n740_), .A2(new_n741_), .A3(new_n742_), .ZN(G1334gat));
  INV_X1    g542(.A(G78gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n726_), .B2(new_n555_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n745_), .A2(new_n746_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n555_), .A2(new_n744_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT111), .ZN(new_n751_));
  OAI22_X1  g550(.A1(new_n748_), .A2(new_n749_), .B1(new_n719_), .B2(new_n751_), .ZN(G1335gat));
  NAND2_X1  g551(.A1(new_n716_), .A2(new_n686_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G85gat), .B1(new_n754_), .B2(new_n648_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n678_), .A2(new_n679_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n609_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n290_), .A2(new_n757_), .A3(new_n326_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n756_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n577_), .A2(new_n210_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n755_), .B1(new_n761_), .B2(new_n762_), .ZN(G1336gat));
  AOI21_X1  g562(.A(G92gat), .B1(new_n754_), .B2(new_n448_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n579_), .A2(new_n211_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n761_), .B2(new_n765_), .ZN(G1337gat));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n379_), .A2(new_n203_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n753_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n761_), .A2(new_n662_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(G99gat), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g571(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n756_), .A2(new_n555_), .A3(new_n760_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(G106gat), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n775_), .A2(new_n774_), .A3(G106gat), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n754_), .A2(new_n204_), .A3(new_n555_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n773_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n778_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n780_), .B(new_n773_), .C1(new_n782_), .C2(new_n776_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n781_), .A2(new_n784_), .ZN(G1339gat));
  XOR2_X1   g584(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n244_), .A2(new_n248_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n247_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n255_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n249_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n283_), .B1(new_n787_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT56), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT56), .B(new_n283_), .C1(new_n787_), .C2(new_n792_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n793_), .A2(KEYINPUT118), .A3(new_n794_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n316_), .B1(new_n315_), .B2(new_n308_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n309_), .A2(new_n311_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n316_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n312_), .A2(new_n317_), .ZN(new_n803_));
  MUX2_X1   g602(.A(new_n802_), .B(new_n803_), .S(new_n320_), .Z(new_n804_));
  AND2_X1   g603(.A1(new_n804_), .A2(new_n278_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n798_), .A2(new_n799_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n798_), .A2(KEYINPUT58), .A3(new_n805_), .A4(new_n799_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n636_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n795_), .A2(new_n797_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n279_), .B2(new_n326_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n278_), .A2(new_n325_), .A3(KEYINPUT115), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n279_), .A2(new_n280_), .A3(new_n202_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT70), .B1(new_n284_), .B2(new_n278_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n804_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n644_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT117), .B1(new_n819_), .B2(KEYINPUT57), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(KEYINPUT57), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n810_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n819_), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n605_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  AND4_X1   g623(.A1(new_n609_), .A2(new_n633_), .A3(new_n635_), .A4(new_n326_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(new_n289_), .A3(new_n288_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n824_), .A2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n648_), .A2(new_n379_), .A3(new_n582_), .A4(new_n580_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n832_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n830_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(G113gat), .B1(new_n838_), .B2(new_n325_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n830_), .B2(new_n836_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n835_), .A2(KEYINPUT59), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n813_), .A2(new_n814_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n846_), .A2(new_n811_), .B1(new_n286_), .B2(new_n804_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n845_), .B1(new_n847_), .B2(new_n644_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n815_), .A2(new_n818_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(KEYINPUT57), .A3(new_n631_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n810_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n757_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n828_), .B1(new_n852_), .B2(KEYINPUT120), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n854_), .A3(new_n757_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n844_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n840_), .B1(new_n842_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n853_), .A2(new_n855_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n843_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n850_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n848_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n823_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n810_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n828_), .B1(new_n864_), .B2(new_n605_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT59), .B1(new_n865_), .B2(new_n835_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n859_), .A2(new_n866_), .A3(KEYINPUT121), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n857_), .A2(new_n867_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n325_), .A2(G113gat), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n839_), .B1(new_n868_), .B2(new_n869_), .ZN(G1340gat));
  INV_X1    g669(.A(new_n290_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n842_), .A2(new_n856_), .A3(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(G120gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n871_), .B2(KEYINPUT60), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(KEYINPUT60), .B2(new_n873_), .ZN(new_n875_));
  OAI22_X1  g674(.A1(new_n872_), .A2(new_n873_), .B1(new_n837_), .B2(new_n875_), .ZN(G1341gat));
  AOI21_X1  g675(.A(G127gat), .B1(new_n838_), .B2(new_n609_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n605_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n878_), .A2(G127gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n868_), .B2(new_n879_), .ZN(G1342gat));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n881_));
  AOI211_X1 g680(.A(new_n631_), .B(new_n835_), .C1(new_n824_), .C2(new_n829_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(G134gat), .ZN(new_n883_));
  INV_X1    g682(.A(G134gat), .ZN(new_n884_));
  OAI211_X1 g683(.A(KEYINPUT122), .B(new_n884_), .C1(new_n837_), .C2(new_n631_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  XOR2_X1   g685(.A(KEYINPUT123), .B(G134gat), .Z(new_n887_));
  NOR2_X1   g686(.A1(new_n637_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n868_), .B2(new_n888_), .ZN(G1343gat));
  NOR2_X1   g688(.A1(new_n662_), .A2(new_n578_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n577_), .A2(new_n448_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n808_), .A2(new_n636_), .A3(new_n809_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n861_), .B2(new_n848_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n878_), .B1(new_n893_), .B2(new_n863_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n890_), .B(new_n891_), .C1(new_n894_), .C2(new_n828_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n325_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n290_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g699(.A(KEYINPUT124), .B1(new_n895_), .B2(new_n757_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n890_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n903_), .A2(new_n904_), .A3(new_n609_), .A4(new_n891_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT61), .B(G155gat), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n901_), .A2(new_n905_), .A3(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n901_), .B2(new_n905_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1346gat));
  INV_X1    g708(.A(G162gat), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n895_), .A2(new_n910_), .A3(new_n637_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n896_), .A2(new_n644_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n910_), .ZN(G1347gat));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n648_), .A2(new_n579_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n916_), .A2(new_n380_), .A3(new_n555_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n858_), .A2(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n326_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n914_), .B1(new_n919_), .B2(new_n349_), .ZN(new_n920_));
  OAI211_X1 g719(.A(KEYINPUT62), .B(G169gat), .C1(new_n918_), .C2(new_n326_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n331_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(G1348gat));
  INV_X1    g722(.A(new_n918_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n408_), .B1(new_n924_), .B2(new_n290_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n830_), .A2(new_n917_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n871_), .A2(new_n350_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n925_), .B1(new_n926_), .B2(new_n927_), .ZN(G1349gat));
  AOI21_X1  g727(.A(new_n342_), .B1(new_n926_), .B2(new_n609_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n605_), .A2(new_n353_), .A3(new_n401_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n924_), .B2(new_n930_), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n918_), .B2(new_n637_), .ZN(new_n932_));
  OR2_X1    g731(.A1(new_n631_), .A2(new_n359_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT125), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n932_), .B1(new_n918_), .B2(new_n934_), .ZN(G1351gat));
  NOR3_X1   g734(.A1(new_n865_), .A2(new_n902_), .A3(new_n916_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n325_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g737(.A1(new_n903_), .A2(new_n915_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n939_), .A2(new_n871_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(G204gat), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n940_), .B(new_n942_), .ZN(G1353gat));
  AOI211_X1 g742(.A(KEYINPUT63), .B(G211gat), .C1(new_n936_), .C2(new_n878_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(KEYINPUT63), .B(G211gat), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n939_), .A2(new_n605_), .A3(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n944_), .A2(new_n946_), .ZN(G1354gat));
  XOR2_X1   g746(.A(KEYINPUT127), .B(G218gat), .Z(new_n948_));
  NOR3_X1   g747(.A1(new_n939_), .A2(new_n637_), .A3(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n936_), .A2(new_n644_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n950_), .B2(new_n948_), .ZN(G1355gat));
endmodule


