//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n819_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_;
  AND2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  AOI22_X1  g001(.A1(new_n202_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G155gat), .B(G162gat), .ZN(new_n204_));
  OAI221_X1 g003(.A(new_n203_), .B1(G141gat), .B2(G148gat), .C1(KEYINPUT1), .C2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT79), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT2), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NOR3_X1   g009(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n211_));
  NOR3_X1   g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n205_), .B1(new_n212_), .B2(new_n204_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT80), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT77), .B(G127gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(G134gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G113gat), .B(G120gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n213_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(new_n214_), .B2(new_n218_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  MUX2_X1   g021(.A(new_n219_), .B(new_n222_), .S(KEYINPUT4), .Z(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G225gat), .A3(G233gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G225gat), .A2(G233gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT0), .B(G57gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(G85gat), .ZN(new_n229_));
  XOR2_X1   g028(.A(G1gat), .B(G29gat), .Z(new_n230_));
  XOR2_X1   g029(.A(new_n229_), .B(new_n230_), .Z(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n231_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n224_), .A2(new_n226_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT20), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G183gat), .A2(G190gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT23), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(G183gat), .B2(G190gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT22), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(KEYINPUT75), .ZN(new_n241_));
  OAI21_X1  g040(.A(G169gat), .B1(new_n241_), .B2(G176gat), .ZN(new_n242_));
  INV_X1    g041(.A(G169gat), .ZN(new_n243_));
  INV_X1    g042(.A(G176gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n239_), .B(new_n242_), .C1(new_n245_), .C2(new_n241_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT26), .B(G190gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT73), .B1(new_n248_), .B2(G183gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT25), .B(G183gat), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n247_), .B(new_n249_), .C1(new_n250_), .C2(KEYINPUT73), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT74), .Z(new_n252_));
  OAI21_X1  g051(.A(new_n238_), .B1(KEYINPUT24), .B2(new_n245_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n245_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT24), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n246_), .B1(new_n252_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT82), .ZN(new_n260_));
  INV_X1    g059(.A(G197gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(G204gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(G197gat), .B(G204gat), .Z(new_n263_));
  OAI211_X1 g062(.A(KEYINPUT21), .B(new_n262_), .C1(new_n263_), .C2(new_n260_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G211gat), .B(G218gat), .Z(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT83), .B(KEYINPUT21), .Z(new_n267_));
  OAI211_X1 g066(.A(new_n264_), .B(new_n266_), .C1(new_n263_), .C2(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n265_), .A2(KEYINPUT84), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(KEYINPUT84), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(KEYINPUT21), .A3(new_n263_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n268_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n236_), .B1(new_n259_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT89), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n253_), .A2(new_n274_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n256_), .B(KEYINPUT88), .ZN(new_n276_));
  OAI221_X1 g075(.A(new_n275_), .B1(new_n274_), .B2(new_n253_), .C1(new_n254_), .C2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(KEYINPUT22), .B(G169gat), .Z(new_n278_));
  OAI211_X1 g077(.A(new_n239_), .B(new_n255_), .C1(G176gat), .C2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT91), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n273_), .B1(new_n281_), .B2(new_n272_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G226gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT19), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n272_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n286_), .B(KEYINPUT20), .C1(new_n272_), .C2(new_n259_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT18), .B(G64gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(G92gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G8gat), .B(G36gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n290_), .B(new_n291_), .Z(new_n292_));
  AND2_X1   g091(.A1(new_n292_), .A2(KEYINPUT32), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n280_), .A2(new_n272_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(new_n284_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n273_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT90), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n287_), .A2(new_n284_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n296_), .A2(KEYINPUT90), .A3(new_n273_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n235_), .B(new_n294_), .C1(new_n302_), .C2(new_n293_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT33), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n234_), .A2(new_n304_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n299_), .A2(new_n292_), .A3(new_n300_), .A4(new_n301_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n292_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n302_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n234_), .A2(new_n304_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n305_), .A2(new_n306_), .A3(new_n308_), .A4(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n222_), .A2(new_n225_), .ZN(new_n311_));
  AOI211_X1 g110(.A(new_n233_), .B(new_n311_), .C1(new_n223_), .C2(new_n225_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n303_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n259_), .B(KEYINPUT30), .ZN(new_n314_));
  XOR2_X1   g113(.A(KEYINPUT78), .B(KEYINPUT31), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(KEYINPUT76), .B(G15gat), .Z(new_n317_));
  NAND2_X1  g116(.A1(G227gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G43gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n316_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G71gat), .B(G99gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n218_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n321_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n214_), .A2(KEYINPUT29), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT81), .B(KEYINPUT28), .Z(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G22gat), .B(G50gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(G228gat), .ZN(new_n331_));
  INV_X1    g130(.A(G233gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n213_), .A2(KEYINPUT29), .ZN(new_n333_));
  AOI211_X1 g132(.A(new_n331_), .B(new_n332_), .C1(new_n333_), .C2(new_n272_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT85), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n213_), .B(KEYINPUT80), .Z(new_n336_));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337_));
  OAI221_X1 g136(.A(new_n272_), .B1(new_n331_), .B2(new_n332_), .C1(new_n336_), .C2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G78gat), .B(G106gat), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n339_), .A2(new_n340_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n330_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT86), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT86), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n330_), .B(new_n345_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT87), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n342_), .A2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n349_), .A2(new_n330_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n341_), .B1(new_n348_), .B2(new_n342_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n313_), .A2(new_n325_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n347_), .A2(new_n324_), .A3(new_n352_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT27), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n359_), .B1(new_n288_), .B2(new_n307_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n306_), .A2(KEYINPUT93), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n306_), .A2(KEYINPUT93), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT94), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT94), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n360_), .A2(new_n362_), .A3(new_n365_), .A4(new_n361_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT27), .B1(new_n308_), .B2(new_n306_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT95), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT95), .ZN(new_n371_));
  AOI211_X1 g170(.A(new_n371_), .B(new_n368_), .C1(new_n364_), .C2(new_n366_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n358_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n353_), .A2(new_n325_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n367_), .A2(new_n369_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT92), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n235_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n356_), .B1(new_n377_), .B2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G29gat), .B(G36gat), .ZN(new_n382_));
  INV_X1    g181(.A(G43gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(G50gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G15gat), .B(G22gat), .ZN(new_n387_));
  INV_X1    g186(.A(G1gat), .ZN(new_n388_));
  INV_X1    g187(.A(G8gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT14), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G1gat), .B(G8gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n386_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n386_), .B(KEYINPUT15), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(new_n396_), .B2(new_n393_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G229gat), .A2(G233gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n386_), .B(new_n394_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(G229gat), .A3(G233gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G113gat), .B(G141gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(new_n243_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(new_n261_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n405_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n381_), .A2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(KEYINPUT10), .B(G99gat), .Z(new_n410_));
  INV_X1    g209(.A(G106gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(G85gat), .B(G92gat), .Z(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT9), .ZN(new_n414_));
  NAND2_X1  g213(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT9), .ZN(new_n416_));
  NOR2_X1   g215(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n417_));
  OAI21_X1  g216(.A(G85gat), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G99gat), .A2(G106gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT6), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n412_), .A2(new_n414_), .A3(new_n418_), .A4(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G99gat), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n411_), .A3(KEYINPUT67), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT67), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(G99gat), .B2(G106gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT7), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT68), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n423_), .A2(new_n425_), .A3(KEYINPUT68), .A4(new_n426_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT66), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n429_), .A2(new_n420_), .A3(new_n430_), .A4(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT8), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n413_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n437_), .B1(new_n436_), .B2(new_n413_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n421_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n396_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G232gat), .A2(G233gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT71), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT34), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT35), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n386_), .B(new_n421_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n441_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n444_), .A2(new_n445_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G190gat), .B(G218gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G134gat), .ZN(new_n452_));
  INV_X1    g251(.A(G162gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(KEYINPUT36), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(KEYINPUT36), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n450_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n448_), .A2(new_n449_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n448_), .A2(new_n449_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n456_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n459_), .A2(KEYINPUT72), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(KEYINPUT37), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n459_), .B(new_n462_), .C1(KEYINPUT72), .C2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G57gat), .B(G64gat), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n470_), .A2(KEYINPUT11), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(KEYINPUT11), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G71gat), .B(G78gat), .ZN(new_n473_));
  OR3_X1    g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n473_), .A3(KEYINPUT11), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(new_n394_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G231gat), .A2(G233gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT17), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT16), .B(G183gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(G211gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(G127gat), .B(G155gat), .Z(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  OR3_X1    g284(.A1(new_n480_), .A2(new_n481_), .A3(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(KEYINPUT17), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n480_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n469_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n476_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n440_), .A2(new_n491_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n421_), .B(new_n476_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(KEYINPUT12), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT12), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n440_), .A2(new_n495_), .A3(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G230gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT64), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT69), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT69), .ZN(new_n501_));
  INV_X1    g300(.A(new_n499_), .ZN(new_n502_));
  AOI211_X1 g301(.A(new_n501_), .B(new_n502_), .C1(new_n494_), .C2(new_n496_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n492_), .A2(new_n493_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n502_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(G120gat), .B(G148gat), .Z(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(G204gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT5), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(new_n244_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n504_), .A2(new_n506_), .A3(new_n511_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n515_), .A2(KEYINPUT13), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(KEYINPUT13), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n518_), .B(KEYINPUT70), .Z(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n409_), .A2(new_n490_), .A3(new_n520_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n521_), .A2(new_n388_), .A3(new_n379_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n522_), .A2(KEYINPUT38), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(KEYINPUT38), .ZN(new_n524_));
  INV_X1    g323(.A(new_n381_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n463_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(new_n489_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n408_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n525_), .A2(new_n527_), .A3(new_n518_), .A4(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(G1gat), .B1(new_n529_), .B2(new_n380_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n523_), .A2(new_n524_), .A3(new_n530_), .ZN(G1324gat));
  OR2_X1    g330(.A1(new_n370_), .A2(new_n372_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(G8gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n521_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(KEYINPUT96), .B(KEYINPUT39), .Z(new_n535_));
  OAI211_X1 g334(.A(G8gat), .B(new_n535_), .C1(new_n529_), .C2(new_n532_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n535_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n379_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n518_), .B(new_n528_), .C1(new_n538_), .C2(new_n356_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n527_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n532_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n537_), .B1(new_n541_), .B2(new_n389_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n534_), .A2(new_n536_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT97), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT97), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n534_), .A2(new_n536_), .A3(new_n542_), .A4(new_n545_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n544_), .A2(KEYINPUT40), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT40), .B1(new_n544_), .B2(new_n546_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(G1325gat));
  INV_X1    g348(.A(G15gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n521_), .A2(new_n550_), .A3(new_n324_), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT98), .Z(new_n552_));
  OAI21_X1  g351(.A(G15gat), .B1(new_n529_), .B2(new_n325_), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n553_), .B(KEYINPUT41), .Z(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(G1326gat));
  OAI21_X1  g354(.A(G22gat), .B1(new_n529_), .B2(new_n354_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT42), .ZN(new_n557_));
  INV_X1    g356(.A(G22gat), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n521_), .A2(new_n558_), .A3(new_n353_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(G1327gat));
  INV_X1    g359(.A(KEYINPUT100), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT43), .B1(new_n381_), .B2(new_n468_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT43), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n563_), .B(new_n469_), .C1(new_n538_), .C2(new_n356_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n518_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n489_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n408_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT99), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT44), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n565_), .A2(KEYINPUT44), .A3(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n561_), .B1(new_n575_), .B2(new_n380_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n569_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n572_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(KEYINPUT100), .A3(new_n379_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n576_), .A2(new_n579_), .A3(G29gat), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n525_), .A2(new_n526_), .A3(new_n568_), .ZN(new_n581_));
  OR3_X1    g380(.A1(new_n581_), .A2(G29gat), .A3(new_n380_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(G1328gat));
  INV_X1    g382(.A(KEYINPUT46), .ZN(new_n584_));
  INV_X1    g383(.A(G36gat), .ZN(new_n585_));
  INV_X1    g384(.A(new_n532_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n578_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n581_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT101), .B(KEYINPUT45), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n584_), .B1(new_n587_), .B2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G36gat), .B1(new_n575_), .B2(new_n532_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n590_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n589_), .B(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(KEYINPUT46), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n596_), .ZN(G1329gat));
  OAI21_X1  g396(.A(new_n383_), .B1(new_n581_), .B2(new_n325_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT102), .Z(new_n599_));
  INV_X1    g398(.A(KEYINPUT47), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n324_), .A2(G43gat), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n599_), .B(new_n600_), .C1(new_n575_), .C2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n575_), .A2(new_n601_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n598_), .B(KEYINPUT102), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT47), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(G1330gat));
  OAI21_X1  g405(.A(G50gat), .B1(new_n575_), .B2(new_n354_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n588_), .A2(new_n385_), .A3(new_n353_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1331gat));
  AOI21_X1  g408(.A(KEYINPUT103), .B1(new_n566_), .B2(new_n490_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n566_), .A2(KEYINPUT103), .A3(new_n490_), .ZN(new_n611_));
  NOR4_X1   g410(.A1(new_n381_), .A2(new_n528_), .A3(new_n610_), .A4(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(G57gat), .B1(new_n612_), .B2(new_n379_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n525_), .A2(new_n527_), .A3(new_n408_), .A4(new_n519_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(new_n380_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n613_), .B1(G57gat), .B2(new_n615_), .ZN(G1332gat));
  INV_X1    g415(.A(G64gat), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n612_), .A2(new_n617_), .A3(new_n586_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G64gat), .B1(new_n614_), .B2(new_n532_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n619_), .A2(KEYINPUT104), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(KEYINPUT104), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n620_), .A2(KEYINPUT48), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT48), .B1(new_n620_), .B2(new_n621_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n618_), .B1(new_n622_), .B2(new_n623_), .ZN(G1333gat));
  OAI21_X1  g423(.A(G71gat), .B1(new_n614_), .B2(new_n325_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT49), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n325_), .A2(G71gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT105), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n612_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(G1334gat));
  OAI21_X1  g429(.A(G78gat), .B1(new_n614_), .B2(new_n354_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT50), .ZN(new_n632_));
  INV_X1    g431(.A(G78gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n612_), .A2(new_n633_), .A3(new_n353_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(G1335gat));
  OAI211_X1 g434(.A(new_n526_), .B(new_n519_), .C1(new_n538_), .C2(new_n356_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n528_), .A2(new_n567_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(KEYINPUT106), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT106), .ZN(new_n640_));
  INV_X1    g439(.A(new_n638_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n640_), .B1(new_n636_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(G85gat), .B1(new_n643_), .B2(new_n379_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n565_), .A2(KEYINPUT107), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n518_), .A2(new_n641_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT108), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT107), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n562_), .A2(new_n649_), .A3(new_n564_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n645_), .A2(new_n648_), .A3(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n651_), .A2(new_n379_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n644_), .B1(new_n652_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g452(.A(G92gat), .B1(new_n643_), .B2(new_n586_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n417_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n532_), .B1(new_n655_), .B2(new_n415_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n654_), .B1(new_n651_), .B2(new_n656_), .ZN(G1337gat));
  NAND3_X1  g456(.A1(new_n645_), .A2(new_n648_), .A3(new_n650_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G99gat), .B1(new_n658_), .B2(new_n325_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n643_), .A2(new_n410_), .A3(new_n324_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT109), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n643_), .A2(KEYINPUT109), .A3(new_n410_), .A4(new_n324_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT51), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT51), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n659_), .A2(new_n662_), .A3(new_n666_), .A4(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1338gat));
  NAND3_X1  g467(.A1(new_n643_), .A2(new_n411_), .A3(new_n353_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n565_), .A2(new_n353_), .A3(new_n648_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT52), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(G106gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n670_), .B2(G106gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT53), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT53), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n676_), .B(new_n669_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1339gat));
  NAND3_X1  g477(.A1(new_n490_), .A2(new_n518_), .A3(new_n408_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT54), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n397_), .A2(G229gat), .A3(G233gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n400_), .A2(new_n398_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n405_), .A3(new_n683_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n406_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n514_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n494_), .A2(KEYINPUT110), .A3(new_n496_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT110), .B1(new_n494_), .B2(new_n496_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n502_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT111), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n497_), .A2(KEYINPUT55), .A3(new_n499_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n497_), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(new_n499_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT55), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n697_), .B1(new_n500_), .B2(new_n503_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT111), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n699_), .B(new_n502_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n691_), .A2(new_n696_), .A3(new_n698_), .A4(new_n700_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n701_), .A2(KEYINPUT56), .A3(new_n512_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT56), .B1(new_n701_), .B2(new_n512_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n687_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT58), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n469_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT114), .ZN(new_n708_));
  INV_X1    g507(.A(new_n703_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n701_), .A2(KEYINPUT56), .A3(new_n512_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n686_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT58), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT114), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n706_), .A2(new_n713_), .A3(new_n469_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n708_), .A2(new_n712_), .A3(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n514_), .B(new_n528_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n515_), .A2(KEYINPUT113), .A3(new_n685_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n515_), .A2(new_n685_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT113), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n716_), .A2(new_n717_), .A3(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(KEYINPUT57), .A3(new_n463_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT57), .B1(new_n721_), .B2(new_n463_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n715_), .A2(new_n722_), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n681_), .B1(new_n725_), .B2(new_n489_), .ZN(new_n726_));
  OR3_X1    g525(.A1(new_n373_), .A2(KEYINPUT115), .A3(new_n380_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT115), .B1(new_n373_), .B2(new_n380_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT59), .B1(new_n726_), .B2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n713_), .B1(new_n706_), .B2(new_n469_), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT114), .B(new_n468_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n712_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n731_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT117), .B1(new_n734_), .B2(new_n723_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT117), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n715_), .A2(new_n736_), .A3(new_n724_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n735_), .A2(new_n722_), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n681_), .B1(new_n738_), .B2(new_n489_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n729_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n730_), .B1(new_n739_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT118), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OAI211_X1 g544(.A(KEYINPUT118), .B(new_n730_), .C1(new_n739_), .C2(new_n742_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n528_), .A2(KEYINPUT119), .A3(G113gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n747_), .B1(KEYINPUT119), .B2(G113gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(new_n746_), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(G113gat), .ZN(new_n750_));
  INV_X1    g549(.A(new_n726_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n740_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n752_), .B2(new_n408_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n749_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT120), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT120), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n749_), .A2(new_n756_), .A3(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1340gat));
  INV_X1    g557(.A(new_n752_), .ZN(new_n759_));
  INV_X1    g558(.A(G120gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(new_n518_), .B2(KEYINPUT60), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n759_), .B(new_n761_), .C1(KEYINPUT60), .C2(new_n760_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n743_), .A2(new_n520_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n762_), .B1(new_n764_), .B2(new_n760_), .ZN(G1341gat));
  AOI21_X1  g564(.A(G127gat), .B1(new_n759_), .B2(new_n567_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n745_), .A2(new_n746_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n567_), .A2(G127gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(G1342gat));
  AOI21_X1  g568(.A(G134gat), .B1(new_n759_), .B2(new_n526_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT121), .B(G134gat), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n468_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n767_), .B2(new_n772_), .ZN(G1343gat));
  NOR2_X1   g572(.A1(new_n726_), .A2(new_n374_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n586_), .A2(new_n380_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT122), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT122), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n774_), .A2(new_n778_), .A3(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n528_), .ZN(new_n781_));
  XOR2_X1   g580(.A(KEYINPUT123), .B(G141gat), .Z(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(G1344gat));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n519_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g584(.A1(new_n780_), .A2(new_n567_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(KEYINPUT61), .B(G155gat), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n786_), .B(new_n787_), .ZN(G1346gat));
  AOI21_X1  g587(.A(G162gat), .B1(new_n780_), .B2(new_n526_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n453_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n469_), .B2(new_n790_), .ZN(G1347gat));
  NAND2_X1  g590(.A1(new_n586_), .A2(new_n380_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n739_), .A2(new_n357_), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n243_), .B1(new_n793_), .B2(new_n528_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n794_), .A2(KEYINPUT62), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(KEYINPUT62), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n793_), .A2(new_n528_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n795_), .B(new_n796_), .C1(new_n278_), .C2(new_n797_), .ZN(G1348gat));
  NOR2_X1   g597(.A1(new_n792_), .A2(new_n325_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n751_), .A2(new_n354_), .A3(new_n799_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n800_), .A2(new_n244_), .A3(new_n520_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT124), .ZN(new_n802_));
  AOI21_X1  g601(.A(G176gat), .B1(new_n793_), .B2(new_n566_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1349gat));
  INV_X1    g603(.A(new_n250_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n793_), .A2(new_n567_), .A3(new_n805_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n806_), .A2(KEYINPUT125), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(KEYINPUT125), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n800_), .A2(new_n489_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(G183gat), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n807_), .A2(new_n808_), .A3(new_n810_), .ZN(G1350gat));
  NAND2_X1  g610(.A1(new_n793_), .A2(new_n469_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G190gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n793_), .A2(new_n526_), .A3(new_n247_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1351gat));
  NOR3_X1   g614(.A1(new_n726_), .A2(new_n374_), .A3(new_n792_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n528_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n519_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g619(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n816_), .A2(new_n567_), .A3(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT126), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(KEYINPUT127), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(KEYINPUT127), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n825_), .B(new_n826_), .Z(G1354gat));
  AOI21_X1  g626(.A(G218gat), .B1(new_n816_), .B2(new_n526_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n816_), .A2(G218gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n469_), .B2(new_n829_), .ZN(G1355gat));
endmodule


