//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n905_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT6), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n205_));
  OR3_X1    g004(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G85gat), .B(G92gat), .Z(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT8), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT65), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n209_), .A2(KEYINPUT8), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(KEYINPUT8), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n208_), .A2(KEYINPUT9), .ZN(new_n219_));
  INV_X1    g018(.A(G85gat), .ZN(new_n220_));
  INV_X1    g019(.A(G92gat), .ZN(new_n221_));
  OR3_X1    g020(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT9), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n218_), .A2(new_n219_), .A3(new_n204_), .A4(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n211_), .A2(new_n215_), .A3(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G71gat), .B(G78gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(G57gat), .B(G64gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(KEYINPUT11), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(KEYINPUT11), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n229_), .A2(KEYINPUT12), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n224_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT66), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G230gat), .A2(G233gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n224_), .A2(new_n234_), .A3(new_n230_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n210_), .A2(new_n223_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT12), .B1(new_n236_), .B2(new_n229_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n229_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n232_), .A2(new_n233_), .A3(new_n235_), .A4(new_n239_), .ZN(new_n240_));
  OR3_X1    g039(.A1(new_n236_), .A2(KEYINPUT64), .A3(new_n229_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n233_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(KEYINPUT64), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n236_), .A2(new_n229_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n241_), .B(new_n242_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT68), .ZN(new_n247_));
  XOR2_X1   g046(.A(G120gat), .B(G148gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G176gat), .B(G204gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n240_), .A2(new_n245_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n240_), .A2(KEYINPUT69), .A3(new_n245_), .A4(new_n251_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n240_), .A2(new_n245_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n256_), .B1(new_n257_), .B2(new_n251_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT13), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n258_), .A2(new_n259_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G15gat), .B(G22gat), .ZN(new_n263_));
  INV_X1    g062(.A(G1gat), .ZN(new_n264_));
  INV_X1    g063(.A(G8gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT14), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G1gat), .B(G8gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G29gat), .B(G36gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G43gat), .B(G50gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n269_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G229gat), .A2(G233gat), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n272_), .B(KEYINPUT15), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n269_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n269_), .B(new_n273_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n275_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n276_), .A2(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G113gat), .B(G141gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(G169gat), .ZN(new_n283_));
  INV_X1    g082(.A(G197gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n281_), .B(new_n285_), .Z(new_n286_));
  NOR2_X1   g085(.A1(new_n262_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT100), .B(KEYINPUT27), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G226gat), .A2(G233gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT19), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n291_));
  INV_X1    g090(.A(G211gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(G218gat), .ZN(new_n293_));
  INV_X1    g092(.A(G218gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(G211gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n291_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(G211gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n292_), .A2(G218gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n298_), .A3(KEYINPUT90), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT21), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT89), .ZN(new_n302_));
  INV_X1    g101(.A(G204gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(G197gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n284_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n304_), .A2(new_n305_), .B1(G197gat), .B2(new_n303_), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n300_), .A2(new_n301_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT88), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n308_), .B1(new_n284_), .B2(G204gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n303_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n284_), .A2(G204gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT21), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n303_), .A2(G197gat), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n284_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT89), .B1(new_n284_), .B2(G204gat), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n301_), .B(new_n314_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n300_), .A2(new_n313_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT91), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n300_), .A2(new_n313_), .A3(KEYINPUT91), .A4(new_n317_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n307_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G183gat), .ZN(new_n325_));
  INV_X1    g124(.A(G190gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT81), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT81), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G169gat), .A3(G176gat), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n329_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT22), .B(G169gat), .ZN(new_n336_));
  INV_X1    g135(.A(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n325_), .A2(KEYINPUT25), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT25), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G183gat), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT26), .B(G190gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n342_), .A2(new_n343_), .B1(new_n330_), .B2(new_n345_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n347_));
  AND3_X1   g146(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n347_), .A2(new_n348_), .A3(new_n323_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n335_), .A2(new_n338_), .B1(new_n346_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT20), .B1(new_n322_), .B2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n345_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n343_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT26), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n355_), .B2(G190gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n349_), .B(new_n352_), .C1(new_n354_), .C2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT22), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT82), .B1(new_n359_), .B2(G169gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT82), .ZN(new_n361_));
  INV_X1    g160(.A(G169gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n362_), .A3(KEYINPUT22), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n363_), .A3(new_n337_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n359_), .A2(KEYINPUT83), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT83), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT22), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n362_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n329_), .B(new_n334_), .C1(new_n364_), .C2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n358_), .A2(new_n369_), .ZN(new_n370_));
  AOI211_X1 g169(.A(new_n307_), .B(new_n370_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n290_), .B1(new_n351_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT96), .ZN(new_n374_));
  XOR2_X1   g173(.A(G8gat), .B(G36gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n377_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT20), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n322_), .B2(new_n350_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n307_), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n301_), .A2(new_n306_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT91), .B1(new_n385_), .B2(new_n313_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n321_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n384_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n370_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n290_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n383_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n372_), .A2(new_n381_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n381_), .B1(new_n372_), .B2(new_n391_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n392_), .B1(new_n393_), .B2(KEYINPUT97), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT97), .ZN(new_n395_));
  AOI211_X1 g194(.A(new_n395_), .B(new_n381_), .C1(new_n372_), .C2(new_n391_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n288_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G155gat), .A2(G162gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n399_), .A2(new_n400_), .A3(KEYINPUT1), .ZN(new_n401_));
  OR2_X1    g200(.A1(G141gat), .A2(G148gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G141gat), .A2(G148gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT84), .B1(new_n401_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n400_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT1), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n398_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n404_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(G141gat), .A2(G148gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n409_), .A2(new_n412_), .A3(new_n413_), .A4(new_n403_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n406_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n399_), .A2(new_n400_), .ZN(new_n416_));
  NOR4_X1   g215(.A1(KEYINPUT85), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT3), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n411_), .B2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT86), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n424_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT2), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n404_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n423_), .A2(new_n425_), .A3(new_n427_), .A4(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n416_), .B1(new_n421_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n415_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT87), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n415_), .A2(new_n430_), .A3(KEYINPUT87), .ZN(new_n434_));
  XOR2_X1   g233(.A(G127gat), .B(G134gat), .Z(new_n435_));
  XOR2_X1   g234(.A(G113gat), .B(G120gat), .Z(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  NAND3_X1  g236(.A1(new_n433_), .A2(new_n434_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n437_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n415_), .A3(new_n430_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G225gat), .A2(G233gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n438_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n438_), .A2(KEYINPUT4), .A3(new_n440_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT4), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n433_), .A2(new_n444_), .A3(new_n434_), .A4(new_n437_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(G225gat), .A3(G233gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n442_), .B1(new_n443_), .B2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G1gat), .B(G29gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT0), .ZN(new_n449_));
  INV_X1    g248(.A(G57gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G85gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n447_), .A2(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n442_), .B(new_n452_), .C1(new_n443_), .C2(new_n446_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n351_), .A2(new_n371_), .A3(new_n290_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n390_), .B1(new_n383_), .B2(new_n389_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT99), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n381_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n379_), .A2(KEYINPUT99), .A3(new_n380_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OAI211_X1 g263(.A(KEYINPUT27), .B(new_n392_), .C1(new_n460_), .C2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n397_), .A2(new_n457_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT94), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n431_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT93), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n431_), .A2(KEYINPUT93), .A3(new_n468_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n388_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G228gat), .A2(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n322_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n433_), .A2(KEYINPUT29), .A3(new_n434_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n473_), .A2(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G78gat), .B(G106gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n467_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n433_), .A2(new_n434_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT29), .ZN(new_n483_));
  XOR2_X1   g282(.A(G22gat), .B(G50gat), .Z(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT28), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n485_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n473_), .A2(new_n475_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n476_), .A2(new_n477_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n480_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n478_), .A2(new_n480_), .ZN(new_n495_));
  OAI22_X1  g294(.A1(new_n481_), .A2(new_n490_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n492_), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT93), .B1(new_n431_), .B2(new_n468_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(new_n322_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n474_), .B1(new_n499_), .B2(new_n472_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n479_), .B1(new_n497_), .B2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n501_), .A2(new_n489_), .A3(new_n467_), .A4(new_n493_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT30), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n370_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n358_), .A2(KEYINPUT30), .A3(new_n369_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G71gat), .B(G99gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G227gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n504_), .A2(new_n505_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n439_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G15gat), .B(G43gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT31), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n510_), .A2(new_n439_), .A3(new_n512_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n514_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n516_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n496_), .A2(new_n502_), .A3(new_n520_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n518_), .A2(new_n519_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n502_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n493_), .A2(KEYINPUT94), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n524_), .A2(new_n489_), .B1(new_n501_), .B2(new_n493_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n522_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n466_), .B1(new_n521_), .B2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n520_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n381_), .A2(KEYINPUT32), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(new_n372_), .A3(new_n391_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n456_), .B(new_n530_), .C1(new_n529_), .C2(new_n460_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n394_), .A2(new_n396_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT98), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n455_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n438_), .A2(new_n440_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n441_), .B(new_n445_), .C1(new_n535_), .C2(new_n444_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n441_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(new_n452_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n534_), .A2(KEYINPUT33), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT33), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n455_), .A2(new_n533_), .A3(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n532_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n528_), .B1(new_n531_), .B2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n527_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n224_), .A2(new_n277_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT71), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  INV_X1    g350(.A(KEYINPUT35), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n553_), .A2(KEYINPUT74), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n210_), .A2(new_n223_), .A3(new_n272_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(KEYINPUT74), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n547_), .A2(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n551_), .A2(new_n552_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT72), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n554_), .A2(KEYINPUT73), .A3(new_n555_), .A4(new_n556_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n560_), .B(new_n561_), .C1(new_n547_), .C2(new_n557_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT75), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(new_n326_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(new_n294_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n563_), .A2(new_n564_), .A3(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n568_), .A2(KEYINPUT36), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n568_), .A2(KEYINPUT36), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT77), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n568_), .A2(KEYINPUT36), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT77), .B1(new_n577_), .B2(new_n572_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT37), .B1(new_n571_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n563_), .A2(new_n564_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n577_), .A2(new_n572_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT37), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n563_), .A2(new_n564_), .A3(new_n570_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n581_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n269_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(new_n229_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G127gat), .B(G155gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT17), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n591_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n591_), .A2(KEYINPUT17), .A3(new_n596_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT79), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n588_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n287_), .A2(new_n545_), .A3(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT101), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n456_), .A2(new_n264_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n202_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT101), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n603_), .B(new_n607_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n608_), .A2(KEYINPUT38), .A3(new_n264_), .A4(new_n456_), .ZN(new_n609_));
  NOR4_X1   g408(.A1(new_n260_), .A2(new_n261_), .A3(new_n286_), .A4(new_n600_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n584_), .A2(new_n586_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n544_), .A2(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G1gat), .B1(new_n615_), .B2(new_n457_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n606_), .A2(new_n609_), .A3(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT102), .ZN(G1324gat));
  AND2_X1   g417(.A1(new_n397_), .A2(new_n465_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n610_), .A2(new_n620_), .A3(new_n613_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n622_), .A3(G8gat), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n622_), .B1(new_n621_), .B2(G8gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT104), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n626_), .A2(KEYINPUT39), .ZN(new_n627_));
  INV_X1    g426(.A(new_n625_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n623_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(new_n630_), .A3(KEYINPUT39), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n608_), .A2(new_n265_), .A3(new_n620_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n627_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n627_), .A2(KEYINPUT40), .A3(new_n631_), .A4(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1325gat));
  INV_X1    g436(.A(G15gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n608_), .A2(new_n638_), .A3(new_n522_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n614_), .B2(new_n522_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT41), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(G1326gat));
  INV_X1    g441(.A(G22gat), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n523_), .A2(new_n525_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n614_), .B2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT42), .Z(new_n646_));
  NAND3_X1  g445(.A1(new_n608_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(G1327gat));
  INV_X1    g449(.A(new_n588_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n651_), .A2(new_n544_), .A3(KEYINPUT43), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT106), .B1(new_n527_), .B2(new_n543_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n526_), .A2(new_n521_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n397_), .A2(new_n457_), .A3(new_n465_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n534_), .A2(KEYINPUT33), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n538_), .A2(new_n536_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n541_), .A3(new_n659_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n393_), .A2(KEYINPUT97), .ZN(new_n661_));
  INV_X1    g460(.A(new_n396_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n662_), .A3(new_n392_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n531_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n528_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n657_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n654_), .A2(new_n588_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(new_n670_), .A3(KEYINPUT43), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n669_), .B2(KEYINPUT43), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n653_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n601_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n262_), .A2(new_n286_), .A3(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n673_), .A2(KEYINPUT44), .A3(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(G29gat), .A3(new_n456_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n669_), .A2(KEYINPUT43), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT107), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n669_), .A2(new_n670_), .A3(KEYINPUT43), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n652_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n675_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n678_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT108), .B(new_n678_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n677_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n544_), .A2(new_n611_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n675_), .A2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G29gat), .B1(new_n690_), .B2(new_n456_), .ZN(new_n691_));
  OR3_X1    g490(.A1(new_n688_), .A2(KEYINPUT109), .A3(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT109), .B1(new_n688_), .B2(new_n691_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1328gat));
  INV_X1    g493(.A(G36gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n690_), .A2(new_n695_), .A3(new_n620_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT45), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n676_), .A2(new_n620_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n699_), .B2(new_n695_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI221_X1 g501(.A(new_n697_), .B1(KEYINPUT110), .B2(KEYINPUT46), .C1(new_n699_), .C2(new_n695_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1329gat));
  NAND3_X1  g503(.A1(new_n676_), .A2(G43gat), .A3(new_n522_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n706_));
  XOR2_X1   g505(.A(KEYINPUT111), .B(G43gat), .Z(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n690_), .B2(new_n522_), .ZN(new_n708_));
  OR3_X1    g507(.A1(new_n706_), .A2(KEYINPUT47), .A3(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT47), .B1(new_n706_), .B2(new_n708_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n690_), .B2(new_n644_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n686_), .A2(new_n687_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n676_), .A2(G50gat), .A3(new_n644_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(G1331gat));
  NOR2_X1   g514(.A1(new_n260_), .A2(new_n261_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n286_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AND4_X1   g517(.A1(new_n545_), .A2(new_n718_), .A3(new_n651_), .A4(new_n674_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n457_), .B1(new_n719_), .B2(KEYINPUT112), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n720_), .B1(KEYINPUT112), .B2(new_n719_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n718_), .A2(new_n674_), .A3(new_n613_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n457_), .A2(new_n450_), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n721_), .A2(new_n450_), .B1(new_n722_), .B2(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n722_), .B2(new_n620_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT48), .Z(new_n727_));
  NAND3_X1  g526(.A1(new_n719_), .A2(new_n725_), .A3(new_n620_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1333gat));
  INV_X1    g528(.A(G71gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n722_), .B2(new_n522_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT49), .Z(new_n732_));
  NAND3_X1  g531(.A1(new_n719_), .A2(new_n730_), .A3(new_n522_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1334gat));
  INV_X1    g533(.A(G78gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n719_), .A2(new_n735_), .A3(new_n644_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n722_), .A2(new_n644_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G78gat), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n738_), .A2(KEYINPUT113), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(KEYINPUT113), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n739_), .A2(KEYINPUT50), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT50), .B1(new_n739_), .B2(new_n740_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n736_), .B1(new_n741_), .B2(new_n742_), .ZN(G1335gat));
  NAND3_X1  g542(.A1(new_n262_), .A2(new_n286_), .A3(new_n601_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n744_), .A2(new_n544_), .A3(new_n611_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G85gat), .B1(new_n745_), .B2(new_n456_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT114), .Z(new_n747_));
  NOR2_X1   g546(.A1(new_n682_), .A2(new_n744_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n457_), .A2(new_n220_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(G1336gat));
  NAND3_X1  g549(.A1(new_n745_), .A2(new_n221_), .A3(new_n620_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n682_), .A2(new_n619_), .A3(new_n744_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(new_n221_), .ZN(G1337gat));
  NAND3_X1  g552(.A1(new_n745_), .A2(new_n522_), .A3(new_n216_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n682_), .A2(new_n520_), .A3(new_n744_), .ZN(new_n755_));
  INV_X1    g554(.A(G99gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g557(.A(new_n744_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n673_), .A2(new_n644_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT116), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n673_), .A2(new_n762_), .A3(new_n644_), .A4(new_n759_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n761_), .A2(G106gat), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n761_), .A2(KEYINPUT52), .A3(G106gat), .A4(new_n763_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n745_), .A2(new_n217_), .A3(new_n644_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT115), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(new_n767_), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n766_), .A2(new_n772_), .A3(new_n769_), .A4(new_n767_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1339gat));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n588_), .A2(new_n717_), .A3(new_n601_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n716_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n716_), .B2(new_n776_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT58), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n281_), .A2(new_n285_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n285_), .B1(new_n279_), .B2(new_n275_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n278_), .A2(new_n274_), .A3(new_n280_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n231_), .A2(KEYINPUT66), .B1(new_n238_), .B2(new_n237_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n233_), .B1(new_n787_), .B2(new_n235_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n240_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n788_), .B1(new_n790_), .B2(KEYINPUT55), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n240_), .A2(new_n789_), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n251_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n786_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n240_), .A2(new_n789_), .A3(new_n792_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n792_), .B1(new_n240_), .B2(new_n789_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n788_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n800_), .A2(new_n251_), .A3(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n780_), .B1(new_n797_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n795_), .B1(new_n800_), .B2(new_n251_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n794_), .A2(new_n801_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(KEYINPUT58), .A4(new_n786_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(new_n588_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n794_), .B2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n800_), .C2(new_n251_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n286_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n258_), .A2(new_n781_), .A3(new_n784_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n612_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n808_), .B1(new_n816_), .B2(KEYINPUT57), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT121), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT121), .B(new_n808_), .C1(new_n816_), .C2(KEYINPUT57), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n821_), .B(new_n612_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n819_), .A2(new_n820_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n779_), .B1(new_n824_), .B2(new_n601_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n620_), .A2(new_n457_), .A3(new_n526_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n827_), .A2(KEYINPUT120), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(KEYINPUT120), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n828_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT122), .B1(new_n825_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n833_));
  INV_X1    g632(.A(new_n831_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n822_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n674_), .B1(new_n835_), .B2(new_n820_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n833_), .B(new_n834_), .C1(new_n836_), .C2(new_n779_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n779_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n600_), .B1(new_n817_), .B2(new_n822_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n826_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT59), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n832_), .A2(new_n717_), .A3(new_n837_), .A4(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(G113gat), .ZN(new_n844_));
  OR3_X1    g643(.A1(new_n841_), .A2(G113gat), .A3(new_n286_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1340gat));
  NAND4_X1  g645(.A1(new_n832_), .A2(new_n262_), .A3(new_n837_), .A4(new_n842_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G120gat), .ZN(new_n848_));
  INV_X1    g647(.A(new_n841_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT60), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n716_), .B2(G120gat), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n849_), .B(new_n851_), .C1(new_n850_), .C2(G120gat), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n848_), .A2(new_n852_), .ZN(G1341gat));
  INV_X1    g652(.A(new_n600_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n832_), .A2(new_n854_), .A3(new_n837_), .A4(new_n842_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G127gat), .ZN(new_n856_));
  OR3_X1    g655(.A1(new_n841_), .A2(G127gat), .A3(new_n601_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1342gat));
  AOI21_X1  g657(.A(G134gat), .B1(new_n849_), .B2(new_n612_), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n832_), .A2(new_n837_), .A3(new_n842_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT123), .B(G134gat), .Z(new_n861_));
  NOR2_X1   g660(.A1(new_n651_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n859_), .B1(new_n860_), .B2(new_n862_), .ZN(G1343gat));
  INV_X1    g662(.A(new_n840_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n521_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n620_), .A2(new_n457_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n717_), .A3(new_n866_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n262_), .A3(new_n866_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g669(.A1(new_n865_), .A2(new_n674_), .A3(new_n866_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  NAND2_X1  g672(.A1(new_n865_), .A2(new_n866_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G162gat), .B1(new_n874_), .B2(new_n651_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n611_), .A2(G162gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n874_), .B2(new_n876_), .ZN(G1347gat));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n619_), .A2(new_n456_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n522_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n644_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n878_), .B1(new_n825_), .B2(new_n882_), .ZN(new_n883_));
  OAI211_X1 g682(.A(KEYINPUT124), .B(new_n881_), .C1(new_n836_), .C2(new_n779_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n717_), .A2(new_n336_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT125), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n884_), .A3(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n717_), .B(new_n881_), .C1(new_n836_), .C2(new_n779_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n888_), .A2(new_n889_), .A3(G169gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n888_), .B2(G169gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n887_), .B1(new_n890_), .B2(new_n891_), .ZN(G1348gat));
  NAND3_X1  g691(.A1(new_n883_), .A2(new_n262_), .A3(new_n884_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n864_), .A2(new_n644_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n716_), .A2(new_n337_), .A3(new_n880_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n893_), .A2(new_n337_), .B1(new_n894_), .B2(new_n895_), .ZN(G1349gat));
  AND2_X1   g695(.A1(new_n883_), .A2(new_n884_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n600_), .A2(new_n342_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n894_), .A2(new_n522_), .A3(new_n674_), .A4(new_n879_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n897_), .A2(new_n898_), .B1(new_n325_), .B2(new_n899_), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n883_), .A2(new_n588_), .A3(new_n884_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G190gat), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n883_), .A2(new_n343_), .A3(new_n612_), .A4(new_n884_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1351gat));
  NAND3_X1  g703(.A1(new_n865_), .A2(new_n717_), .A3(new_n879_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g705(.A1(new_n865_), .A2(new_n262_), .A3(new_n879_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g707(.A1(new_n865_), .A2(new_n854_), .A3(new_n879_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n909_), .A2(new_n910_), .A3(new_n292_), .ZN(new_n911_));
  XOR2_X1   g710(.A(KEYINPUT63), .B(G211gat), .Z(new_n912_));
  NAND4_X1  g711(.A1(new_n865_), .A2(new_n854_), .A3(new_n879_), .A4(new_n912_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n911_), .A2(new_n913_), .ZN(G1354gat));
  AND2_X1   g713(.A1(new_n865_), .A2(new_n879_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT126), .B(G218gat), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n651_), .A2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n865_), .A2(new_n612_), .A3(new_n879_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n915_), .A2(new_n917_), .B1(new_n918_), .B2(new_n916_), .ZN(G1355gat));
endmodule


