//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n598_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n832_,
    new_n834_, new_n835_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G1gat), .A2(G8gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT14), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n202_), .A2(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(G1gat), .A2(G8gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(new_n203_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND4_X1  g007(.A1(new_n202_), .A2(new_n203_), .A3(new_n206_), .A4(new_n204_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G29gat), .B(G36gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT69), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n213_), .A2(KEYINPUT69), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n212_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n213_), .A2(KEYINPUT69), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(new_n214_), .A3(new_n211_), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n217_), .A2(KEYINPUT15), .A3(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT15), .B1(new_n217_), .B2(new_n219_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n210_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G229gat), .A2(G233gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT73), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR3_X1   g024(.A1(new_n215_), .A2(new_n216_), .A3(new_n212_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n211_), .B1(new_n218_), .B2(new_n214_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n210_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n225_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n219_), .A3(new_n217_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n210_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n223_), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n222_), .A2(new_n230_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G169gat), .B(G197gat), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n236_), .B(new_n237_), .Z(new_n238_));
  INV_X1    g037(.A(KEYINPUT75), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT74), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT74), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n235_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(new_n239_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n238_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n241_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT96), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT95), .B(KEYINPUT27), .Z(new_n249_));
  NOR2_X1   g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT24), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT23), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G169gat), .A2(G176gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT24), .ZN(new_n257_));
  INV_X1    g056(.A(G183gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT76), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT76), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT25), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n258_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT77), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G190gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(new_n259_), .B2(G183gat), .ZN(new_n267_));
  OAI221_X1 g066(.A(new_n255_), .B1(new_n250_), .B2(new_n257_), .C1(new_n265_), .C2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n254_), .B1(G183gat), .B2(G190gat), .ZN(new_n269_));
  INV_X1    g068(.A(G169gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(KEYINPUT78), .B2(KEYINPUT22), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT79), .B(G176gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(KEYINPUT78), .A3(KEYINPUT22), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n269_), .B(new_n256_), .C1(new_n271_), .C2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n268_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G204gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT84), .B1(new_n277_), .B2(G197gat), .ZN(new_n278_));
  INV_X1    g077(.A(G197gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n278_), .B1(new_n279_), .B2(G204gat), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n277_), .A2(KEYINPUT84), .A3(G197gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT21), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G211gat), .B(G218gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT85), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(G197gat), .B2(new_n277_), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n279_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n286_));
  OAI22_X1  g085(.A1(new_n285_), .A2(new_n286_), .B1(G197gat), .B2(new_n277_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n282_), .B(new_n283_), .C1(new_n287_), .C2(KEYINPUT21), .ZN(new_n288_));
  INV_X1    g087(.A(new_n283_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(KEYINPUT21), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT20), .B1(new_n276_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT88), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT22), .B(G169gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n272_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n256_), .B(KEYINPUT90), .Z(new_n297_));
  NAND3_X1  g096(.A1(new_n269_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n298_), .B(KEYINPUT91), .Z(new_n299_));
  AOI21_X1  g098(.A(new_n250_), .B1(new_n257_), .B2(KEYINPUT89), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(KEYINPUT89), .B2(new_n257_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT25), .B(G183gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n266_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n255_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n299_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n291_), .ZN(new_n306_));
  OAI211_X1 g105(.A(KEYINPUT88), .B(KEYINPUT20), .C1(new_n276_), .C2(new_n291_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n294_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G226gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT19), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT20), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(new_n276_), .B2(new_n291_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n310_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n313_), .B(new_n314_), .C1(new_n305_), .C2(new_n291_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G8gat), .B(G36gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT18), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G64gat), .B(G92gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n318_), .B(new_n319_), .Z(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n320_), .B1(new_n311_), .B2(new_n315_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n249_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n308_), .A2(new_n310_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n288_), .A2(new_n304_), .A3(new_n290_), .A4(new_n298_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n314_), .B1(new_n313_), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n321_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n328_), .B(KEYINPUT27), .C1(new_n321_), .C2(new_n316_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n324_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n334_), .B(KEYINPUT3), .Z(new_n335_));
  NAND2_X1  g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n336_), .B(KEYINPUT2), .Z(new_n337_));
  OAI211_X1 g136(.A(new_n331_), .B(new_n333_), .C1(new_n335_), .C2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n332_), .B1(KEYINPUT1), .B2(new_n331_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(KEYINPUT1), .B2(new_n331_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n334_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(new_n336_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT28), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G22gat), .B(G50gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n291_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G228gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n355_), .A2(KEYINPUT86), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n354_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n355_), .B2(KEYINPUT86), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n349_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  OR3_X1    g158(.A1(new_n352_), .A2(KEYINPUT87), .A3(new_n354_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT87), .B1(new_n352_), .B2(new_n354_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n360_), .A2(new_n348_), .A3(new_n361_), .A4(new_n357_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n248_), .B1(new_n330_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n363_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n365_), .A2(new_n324_), .A3(KEYINPUT96), .A4(new_n329_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G127gat), .B(G134gat), .Z(new_n368_));
  XOR2_X1   g167(.A(G113gat), .B(G120gat), .Z(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n343_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n338_), .A2(new_n342_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n370_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT93), .B(KEYINPUT4), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n372_), .A2(KEYINPUT4), .A3(new_n374_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n380_), .A2(KEYINPUT92), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(KEYINPUT92), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n379_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n377_), .B1(new_n383_), .B2(new_n376_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G1gat), .B(G29gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(G85gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT0), .B(G57gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  NAND2_X1  g187(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n388_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n390_), .B(new_n377_), .C1(new_n383_), .C2(new_n376_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT82), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G71gat), .B(G99gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(KEYINPUT80), .B(KEYINPUT30), .Z(new_n398_));
  XOR2_X1   g197(.A(new_n397_), .B(new_n398_), .Z(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(G15gat), .B(G43gat), .Z(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT81), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n276_), .B(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT31), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n403_), .A2(new_n404_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n400_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n407_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(new_n399_), .A3(new_n405_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT83), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n408_), .A2(new_n410_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n371_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n412_), .A2(new_n370_), .A3(new_n414_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n367_), .A2(new_n393_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n383_), .A2(new_n376_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n390_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT94), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT94), .ZN(new_n425_));
  AOI211_X1 g224(.A(new_n425_), .B(new_n422_), .C1(new_n383_), .C2(new_n376_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n322_), .A2(new_n323_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT33), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n389_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n384_), .A2(KEYINPUT33), .A3(new_n388_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n427_), .A2(new_n428_), .A3(new_n430_), .A4(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n320_), .A2(KEYINPUT32), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n433_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n392_), .B(new_n434_), .C1(new_n433_), .C2(new_n316_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n363_), .B1(new_n432_), .B2(new_n435_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n330_), .A2(new_n365_), .A3(new_n392_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n418_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n247_), .B1(new_n420_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G190gat), .B(G218gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G134gat), .B(G162gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n442_), .B(KEYINPUT36), .Z(new_n443_));
  OR2_X1    g242(.A1(new_n220_), .A2(new_n221_), .ZN(new_n444_));
  OR2_X1    g243(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n445_));
  OR2_X1    g244(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .A4(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G85gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(KEYINPUT9), .ZN(new_n451_));
  AND2_X1   g250(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G92gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G85gat), .A2(G92gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(KEYINPUT9), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G99gat), .A2(G106gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT6), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT6), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(G99gat), .A3(G106gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n449_), .A2(new_n454_), .A3(new_n458_), .A4(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(G99gat), .A2(G106gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT7), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n463_), .A2(new_n465_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT8), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n456_), .A2(new_n457_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n470_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n464_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n444_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT70), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT70), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n444_), .A2(new_n477_), .A3(new_n474_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G232gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT35), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n464_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n460_), .A2(new_n462_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n468_), .A2(new_n465_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n471_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT8), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n486_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n492_), .A2(new_n228_), .B1(new_n483_), .B2(new_n482_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n479_), .A2(new_n485_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n485_), .B1(new_n479_), .B2(new_n493_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n443_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n479_), .A2(new_n493_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n484_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n442_), .A2(KEYINPUT36), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(new_n494_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT37), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n497_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(new_n497_), .B2(new_n501_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G57gat), .B(G64gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G71gat), .B(G78gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(KEYINPUT11), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(KEYINPUT11), .ZN(new_n509_));
  INV_X1    g308(.A(new_n507_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n506_), .A2(KEYINPUT11), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n508_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT12), .B1(new_n474_), .B2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n513_), .B(new_n464_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT67), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G230gat), .A2(G233gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n474_), .A2(KEYINPUT12), .A3(new_n514_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .A4(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT12), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(new_n492_), .B2(new_n513_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n524_), .A2(new_n521_), .A3(new_n520_), .A4(new_n516_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT67), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n492_), .A2(new_n513_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n520_), .B1(new_n528_), .B2(KEYINPUT66), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n517_), .A2(KEYINPUT66), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n529_), .B1(new_n530_), .B2(new_n528_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G120gat), .B(G148gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT5), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G176gat), .B(G204gat), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n534_), .B(new_n535_), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n536_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n527_), .A2(new_n531_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT13), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(KEYINPUT13), .A3(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G231gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n210_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(new_n513_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT72), .B(KEYINPUT17), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G127gat), .B(G155gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT16), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G183gat), .B(G211gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n553_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n547_), .ZN(new_n556_));
  XOR2_X1   g355(.A(KEYINPUT71), .B(KEYINPUT17), .Z(new_n557_));
  AOI22_X1  g356(.A1(new_n554_), .A2(new_n555_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n505_), .A2(new_n544_), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n439_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n439_), .A2(KEYINPUT97), .A3(new_n559_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n393_), .A2(G1gat), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(KEYINPUT98), .A3(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n562_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT98), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n566_), .A2(KEYINPUT38), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n497_), .A2(new_n501_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n420_), .B2(new_n438_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n558_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n544_), .A2(new_n247_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(G1gat), .B1(new_n576_), .B2(new_n393_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT38), .B1(new_n566_), .B2(new_n569_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n578_), .A2(KEYINPUT99), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(KEYINPUT99), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n570_), .B(new_n577_), .C1(new_n579_), .C2(new_n580_), .ZN(G1324gat));
  INV_X1    g380(.A(G8gat), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n564_), .A2(new_n582_), .A3(new_n330_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n330_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n576_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n585_), .A2(G8gat), .A3(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n586_), .B1(new_n585_), .B2(G8gat), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n583_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n589_), .B(new_n590_), .Z(G1325gat));
  OAI21_X1  g390(.A(G15gat), .B1(new_n576_), .B2(new_n418_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT41), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n560_), .A2(G15gat), .A3(new_n418_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(G1326gat));
  OAI21_X1  g394(.A(G22gat), .B1(new_n576_), .B2(new_n365_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT42), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n365_), .A2(G22gat), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n597_), .B1(new_n560_), .B2(new_n598_), .ZN(G1327gat));
  NOR3_X1   g398(.A1(new_n544_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n439_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(G29gat), .B1(new_n602_), .B2(new_n392_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT43), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(KEYINPUT102), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n432_), .A2(new_n435_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n365_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n437_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n419_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n416_), .A2(new_n393_), .A3(new_n417_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n505_), .B(new_n606_), .C1(new_n610_), .C2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n504_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n497_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n420_), .B2(new_n438_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n613_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n544_), .A2(new_n247_), .A3(new_n574_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n619_), .A2(KEYINPUT44), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT44), .B1(new_n619_), .B2(new_n620_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n392_), .A2(G29gat), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n603_), .B1(new_n623_), .B2(new_n624_), .ZN(G1328gat));
  NAND2_X1  g424(.A1(new_n619_), .A2(new_n620_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT44), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n619_), .A2(KEYINPUT44), .A3(new_n620_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n330_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G36gat), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n584_), .A2(G36gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n602_), .A2(KEYINPUT45), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT45), .ZN(new_n634_));
  INV_X1    g433(.A(new_n632_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n601_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n631_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT46), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n637_), .B1(new_n630_), .B2(G36gat), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT46), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n642_), .A2(KEYINPUT103), .A3(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n641_), .A2(new_n644_), .ZN(G1329gat));
  NAND3_X1  g444(.A1(new_n623_), .A2(G43gat), .A3(new_n419_), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT104), .B(G43gat), .Z(new_n647_));
  OAI21_X1  g446(.A(new_n647_), .B1(new_n601_), .B2(new_n418_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(G1330gat));
  AOI21_X1  g450(.A(G50gat), .B1(new_n602_), .B2(new_n363_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n363_), .A2(G50gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n623_), .B2(new_n653_), .ZN(G1331gat));
  OAI21_X1  g453(.A(new_n247_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT106), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n656_), .A2(new_n544_), .A3(new_n616_), .A4(new_n574_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT107), .ZN(new_n658_));
  INV_X1    g457(.A(G57gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n659_), .A3(new_n392_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n558_), .A2(new_n246_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n573_), .A2(new_n544_), .A3(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G57gat), .B1(new_n662_), .B2(new_n393_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n663_), .ZN(G1332gat));
  INV_X1    g463(.A(G64gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n658_), .A2(new_n665_), .A3(new_n330_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G64gat), .B1(new_n662_), .B2(new_n584_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT48), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1333gat));
  INV_X1    g468(.A(G71gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n658_), .A2(new_n670_), .A3(new_n419_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G71gat), .B1(new_n662_), .B2(new_n418_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT49), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(G1334gat));
  INV_X1    g473(.A(G78gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n658_), .A2(new_n675_), .A3(new_n363_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G78gat), .B1(new_n662_), .B2(new_n365_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT50), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1335gat));
  INV_X1    g478(.A(new_n544_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n680_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n656_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n450_), .A3(new_n392_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n680_), .A2(new_n246_), .A3(new_n574_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n619_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G85gat), .B1(new_n685_), .B2(new_n393_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(G1336gat));
  NOR2_X1   g486(.A1(new_n452_), .A2(new_n453_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n685_), .A2(new_n584_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n682_), .A2(new_n330_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(new_n455_), .ZN(G1337gat));
  AND3_X1   g490(.A1(new_n419_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n656_), .A2(new_n681_), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n696_), .A2(KEYINPUT51), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n619_), .A2(new_n419_), .A3(new_n684_), .ZN(new_n698_));
  AOI22_X1  g497(.A1(new_n698_), .A2(G99gat), .B1(new_n696_), .B2(KEYINPUT51), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n695_), .A2(new_n697_), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n697_), .B1(new_n695_), .B2(new_n699_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1338gat));
  NAND4_X1  g501(.A1(new_n682_), .A2(new_n363_), .A3(new_n446_), .A4(new_n448_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT52), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n619_), .A2(new_n363_), .A3(new_n684_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(G106gat), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n705_), .A2(new_n704_), .A3(G106gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g508(.A1(new_n367_), .A2(new_n392_), .A3(new_n419_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n712_));
  AND2_X1   g511(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT55), .B1(new_n522_), .B2(new_n526_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n520_), .A2(KEYINPUT111), .ZN(new_n716_));
  AND4_X1   g515(.A1(new_n521_), .A2(new_n524_), .A3(new_n516_), .A4(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n716_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT55), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n520_), .A2(new_n719_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n524_), .A2(new_n521_), .A3(new_n516_), .A4(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n717_), .B1(new_n718_), .B2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT56), .B(new_n536_), .C1(new_n715_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT116), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n536_), .B1(new_n715_), .B2(new_n722_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT56), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n726_), .A2(new_n724_), .A3(new_n727_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n233_), .A2(new_n224_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n245_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n222_), .A2(new_n231_), .A3(new_n225_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n225_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT113), .B1(new_n736_), .B2(new_n238_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n734_), .A2(new_n735_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n235_), .A2(new_n238_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(KEYINPUT114), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT114), .B1(new_n738_), .B2(new_n739_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n539_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n539_), .B(KEYINPUT115), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n714_), .B1(new_n731_), .B2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(KEYINPUT118), .B1(new_n747_), .B2(new_n616_), .ZN(new_n748_));
  AOI22_X1  g547(.A1(new_n729_), .A2(new_n730_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT58), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT118), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n505_), .B(new_n751_), .C1(new_n749_), .C2(new_n714_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n750_), .A3(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n728_), .A2(new_n754_), .A3(new_n723_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n726_), .A2(KEYINPUT112), .A3(new_n727_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n246_), .A2(new_n539_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n540_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT57), .B1(new_n760_), .B2(new_n571_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT57), .ZN(new_n762_));
  AOI211_X1 g561(.A(new_n762_), .B(new_n572_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n574_), .B1(new_n753_), .B2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n542_), .A2(new_n543_), .A3(new_n661_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT110), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n542_), .A2(new_n768_), .A3(new_n543_), .A4(new_n661_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n616_), .A2(new_n767_), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT54), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n616_), .A2(new_n767_), .A3(new_n772_), .A4(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  OAI221_X1 g574(.A(new_n711_), .B1(new_n712_), .B2(new_n713_), .C1(new_n765_), .C2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n753_), .A2(new_n764_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n558_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(KEYINPUT119), .A3(new_n774_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT119), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n765_), .B2(new_n775_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n783_), .A2(new_n710_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT59), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n776_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G113gat), .B1(new_n786_), .B2(new_n247_), .ZN(new_n787_));
  INV_X1    g586(.A(G113gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n784_), .A2(new_n788_), .A3(new_n246_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1340gat));
  OAI21_X1  g589(.A(G120gat), .B1(new_n786_), .B2(new_n680_), .ZN(new_n791_));
  INV_X1    g590(.A(G120gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(new_n680_), .B2(KEYINPUT60), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n784_), .B(new_n793_), .C1(KEYINPUT60), .C2(new_n792_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(new_n794_), .ZN(G1341gat));
  OAI21_X1  g594(.A(G127gat), .B1(new_n786_), .B2(new_n558_), .ZN(new_n796_));
  INV_X1    g595(.A(G127gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n784_), .A2(new_n797_), .A3(new_n574_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1342gat));
  AND2_X1   g598(.A1(new_n505_), .A2(G134gat), .ZN(new_n800_));
  XOR2_X1   g599(.A(new_n800_), .B(KEYINPUT121), .Z(new_n801_));
  OR2_X1    g600(.A1(new_n786_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(G134gat), .B1(new_n784_), .B2(new_n572_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1343gat));
  NAND3_X1  g604(.A1(new_n418_), .A2(new_n363_), .A3(new_n392_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n783_), .A2(new_n330_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n246_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n544_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g610(.A1(new_n807_), .A2(new_n574_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(KEYINPUT61), .B(G155gat), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n812_), .B(new_n813_), .ZN(G1346gat));
  INV_X1    g613(.A(G162gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n807_), .A2(new_n815_), .A3(new_n572_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n807_), .A2(new_n505_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n815_), .ZN(G1347gat));
  AOI21_X1  g617(.A(new_n363_), .B1(new_n778_), .B2(new_n774_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n611_), .A2(new_n584_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n821_), .A2(new_n247_), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n270_), .B(new_n822_), .C1(KEYINPUT122), .C2(KEYINPUT62), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(KEYINPUT122), .B2(KEYINPUT62), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT62), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n825_), .B(new_n826_), .C1(new_n822_), .C2(new_n270_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n822_), .A2(new_n295_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n824_), .A2(new_n827_), .A3(new_n828_), .ZN(G1348gat));
  NOR2_X1   g628(.A1(new_n783_), .A2(new_n363_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n820_), .A2(G176gat), .A3(new_n544_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n819_), .A2(new_n544_), .A3(new_n820_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n830_), .A2(new_n831_), .B1(new_n272_), .B2(new_n832_), .ZN(G1349gat));
  NAND3_X1  g632(.A1(new_n830_), .A2(new_n574_), .A3(new_n820_), .ZN(new_n834_));
  NOR4_X1   g633(.A1(new_n611_), .A2(new_n302_), .A3(new_n584_), .A4(new_n558_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n834_), .A2(new_n258_), .B1(new_n819_), .B2(new_n835_), .ZN(G1350gat));
  OAI21_X1  g635(.A(G190gat), .B1(new_n821_), .B2(new_n616_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n572_), .A2(new_n266_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n821_), .B2(new_n838_), .ZN(G1351gat));
  NOR2_X1   g638(.A1(new_n365_), .A2(new_n392_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n418_), .A2(new_n840_), .A3(new_n330_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n783_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n246_), .ZN(new_n843_));
  OR3_X1    g642(.A1(new_n843_), .A2(KEYINPUT123), .A3(new_n279_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT123), .B1(new_n843_), .B2(new_n279_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n279_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(G1352gat));
  INV_X1    g646(.A(new_n841_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT119), .B1(new_n778_), .B2(new_n774_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n765_), .A2(new_n780_), .A3(new_n775_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n544_), .B(new_n848_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n782_), .A2(KEYINPUT124), .A3(new_n544_), .A4(new_n848_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(G204gat), .A3(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT125), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n680_), .B(new_n841_), .C1(new_n779_), .C2(new_n781_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n277_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT126), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n853_), .A2(new_n856_), .A3(G204gat), .A4(new_n854_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1353gat));
  INV_X1    g663(.A(KEYINPUT63), .ZN(new_n865_));
  INV_X1    g664(.A(G211gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(KEYINPUT127), .ZN(new_n867_));
  NAND2_X1  g666(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n842_), .A2(new_n574_), .A3(new_n867_), .A4(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT127), .B1(new_n865_), .B2(new_n866_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1354gat));
  INV_X1    g670(.A(G218gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n842_), .A2(new_n872_), .A3(new_n572_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n783_), .A2(new_n616_), .A3(new_n841_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n872_), .ZN(G1355gat));
endmodule


