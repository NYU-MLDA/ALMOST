//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G71gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT89), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G169gat), .ZN(new_n209_));
  INV_X1    g008(.A(G176gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  OR3_X1    g010(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT23), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n213_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G190gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT86), .B1(new_n221_), .B2(KEYINPUT26), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n222_), .B(new_n223_), .C1(new_n224_), .C2(KEYINPUT86), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT87), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n225_), .A2(KEYINPUT87), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n220_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G169gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n218_), .A2(KEYINPUT88), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n217_), .A2(KEYINPUT88), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n230_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n206_), .B1(new_n228_), .B2(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n227_), .A2(new_n226_), .ZN(new_n238_));
  OAI211_X1 g037(.A(KEYINPUT89), .B(new_n235_), .C1(new_n238_), .C2(new_n220_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G15gat), .B(G43gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT90), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT30), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n240_), .A2(new_n244_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n205_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n247_), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n249_), .A2(new_n245_), .A3(new_n204_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G127gat), .B(G134gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G113gat), .B(G120gat), .Z(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT92), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G113gat), .B(G120gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n255_), .B(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT31), .Z(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT91), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(G99gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n251_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G225gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT102), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n253_), .A2(new_n254_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n257_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT101), .ZN(new_n269_));
  XOR2_X1   g068(.A(G155gat), .B(G162gat), .Z(new_n270_));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n273_));
  INV_X1    g072(.A(G141gat), .ZN(new_n274_));
  INV_X1    g073(.A(G148gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n274_), .A2(new_n275_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n272_), .A2(new_n273_), .A3(new_n276_), .A4(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n274_), .A2(new_n275_), .A3(KEYINPUT93), .ZN(new_n280_));
  AOI22_X1  g079(.A1(KEYINPUT2), .A2(new_n277_), .B1(new_n280_), .B2(KEYINPUT3), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(KEYINPUT3), .B2(new_n280_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(KEYINPUT94), .Z(new_n284_));
  OAI21_X1  g083(.A(new_n270_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n269_), .A2(new_n279_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n279_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n258_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n266_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT4), .B1(new_n287_), .B2(new_n258_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n265_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n265_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n286_), .A2(new_n292_), .A3(new_n288_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G1gat), .B(G29gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(G85gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT0), .B(G57gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n295_), .B(new_n296_), .Z(new_n297_));
  NAND3_X1  g096(.A1(new_n291_), .A2(new_n293_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n297_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n261_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n263_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G8gat), .B(G36gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(G64gat), .B(G92gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G197gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(G204gat), .ZN(new_n311_));
  INV_X1    g110(.A(G204gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G197gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT21), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G211gat), .B(G218gat), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n315_), .B1(KEYINPUT98), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n317_), .B1(KEYINPUT98), .B2(new_n316_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n314_), .A2(KEYINPUT97), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT97), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT21), .B1(new_n311_), .B2(new_n320_), .ZN(new_n321_));
  OAI221_X1 g120(.A(new_n316_), .B1(KEYINPUT21), .B2(new_n314_), .C1(new_n319_), .C2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT19), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n230_), .B1(new_n218_), .B2(new_n234_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n231_), .A2(new_n232_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n224_), .A2(new_n223_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n331_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n330_), .A2(KEYINPUT99), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT99), .B1(new_n330_), .B2(new_n332_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n329_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n328_), .B1(new_n335_), .B2(new_n323_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT20), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n325_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(new_n335_), .B2(new_n323_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n237_), .A2(new_n239_), .A3(new_n324_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n328_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n309_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n340_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n327_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n240_), .A2(new_n323_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n329_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n334_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n330_), .A2(KEYINPUT99), .A3(new_n332_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n346_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n327_), .B1(new_n349_), .B2(new_n324_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n345_), .A2(new_n350_), .A3(KEYINPUT20), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n344_), .A2(new_n351_), .A3(new_n308_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n342_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT27), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n339_), .A2(new_n340_), .A3(new_n328_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n330_), .A2(new_n332_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n324_), .A2(new_n329_), .A3(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n345_), .A2(KEYINPUT20), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n356_), .B1(new_n327_), .B2(new_n359_), .ZN(new_n360_));
  OAI211_X1 g159(.A(KEYINPUT27), .B(new_n352_), .C1(new_n360_), .C2(new_n308_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n285_), .A2(new_n279_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364_));
  XOR2_X1   g163(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n287_), .B2(KEYINPUT29), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G22gat), .B(G50gat), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n370_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n367_), .A2(new_n372_), .A3(new_n368_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT96), .B1(new_n318_), .B2(new_n322_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377_));
  INV_X1    g176(.A(G78gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(G106gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n381_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n383_), .B(new_n375_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n374_), .A2(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n371_), .A2(new_n373_), .A3(new_n382_), .A4(new_n384_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(new_n303_), .A2(new_n362_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n300_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n388_), .A2(new_n390_), .A3(new_n298_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(new_n355_), .A3(new_n361_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT104), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n298_), .B(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n297_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n286_), .A2(new_n288_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n397_), .B1(new_n398_), .B2(new_n292_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT103), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n292_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n402_));
  OAI211_X1 g201(.A(KEYINPUT103), .B(new_n397_), .C1(new_n398_), .C2(new_n292_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n342_), .A2(new_n352_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n308_), .A2(KEYINPUT32), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n344_), .A2(new_n351_), .A3(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n407_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n359_), .A2(new_n327_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n356_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n406_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  OAI22_X1  g210(.A1(new_n396_), .A2(new_n405_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n388_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n391_), .A2(new_n355_), .A3(new_n361_), .A4(KEYINPUT104), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n394_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n263_), .A2(new_n302_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n389_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G113gat), .B(G141gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G169gat), .B(G197gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT84), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(G29gat), .B(G36gat), .Z(new_n424_));
  XOR2_X1   g223(.A(G43gat), .B(G50gat), .Z(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G29gat), .B(G36gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G43gat), .B(G50gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n426_), .A2(KEYINPUT81), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT81), .B1(new_n426_), .B2(new_n429_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT79), .B(G1gat), .ZN(new_n433_));
  INV_X1    g232(.A(G8gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT14), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G15gat), .B(G22gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G1gat), .B(G8gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n435_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n432_), .A2(new_n442_), .A3(KEYINPUT82), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT82), .B1(new_n432_), .B2(new_n442_), .ZN(new_n445_));
  OAI22_X1  g244(.A1(new_n444_), .A2(new_n445_), .B1(new_n442_), .B2(new_n432_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G229gat), .A2(G233gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n426_), .A2(new_n429_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(new_n441_), .A4(new_n440_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n451_), .A2(new_n452_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT83), .B1(new_n456_), .B2(new_n442_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n432_), .A2(new_n442_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT82), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n443_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n462_), .A3(new_n447_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n423_), .B1(new_n449_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n449_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n422_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n421_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n464_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n418_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G85gat), .B(G92gat), .Z(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT10), .B(G99gat), .Z(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n380_), .ZN(new_n475_));
  INV_X1    g274(.A(G85gat), .ZN(new_n476_));
  INV_X1    g275(.A(G92gat), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT9), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G85gat), .B(G92gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT64), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT6), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(G99gat), .A3(G106gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n473_), .A2(new_n475_), .A3(new_n481_), .A4(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT8), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT66), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n489_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n494_));
  INV_X1    g293(.A(G99gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n380_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(KEYINPUT66), .A3(new_n490_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n486_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n488_), .B1(new_n498_), .B2(new_n472_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n479_), .A2(KEYINPUT8), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n483_), .A2(new_n485_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n496_), .A2(new_n490_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT65), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n491_), .A2(new_n492_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT65), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(new_n486_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n501_), .B1(new_n504_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n487_), .B1(new_n499_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n453_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G232gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT35), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n426_), .A2(new_n429_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n510_), .B(new_n515_), .C1(new_n516_), .C2(new_n509_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n513_), .A2(new_n514_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n518_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G190gat), .B(G218gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT74), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G134gat), .B(G162gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n526_), .B(KEYINPUT75), .Z(new_n527_));
  NAND3_X1  g326(.A1(new_n519_), .A2(new_n520_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n519_), .A2(new_n520_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n530_), .A2(KEYINPUT77), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n524_), .B(new_n525_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n530_), .B2(KEYINPUT77), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n529_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT78), .B(KEYINPUT37), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n532_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT76), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n528_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT37), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G231gat), .A2(G233gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n543_), .B(KEYINPUT80), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n442_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(G64gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(G57gat), .ZN(new_n547_));
  INV_X1    g346(.A(G57gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(G64gat), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n549_), .A3(KEYINPUT11), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT68), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G57gat), .B(G64gat), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT68), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(KEYINPUT11), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT67), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT11), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n548_), .A2(G64gat), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n546_), .A2(G57gat), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n203_), .A2(G78gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n378_), .A2(G71gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n556_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT11), .B1(new_n547_), .B2(new_n549_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G71gat), .B(G78gat), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n565_), .A2(KEYINPUT67), .A3(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n555_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT67), .B1(new_n565_), .B2(new_n566_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n563_), .B(new_n556_), .C1(new_n552_), .C2(KEYINPUT11), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n569_), .A2(new_n551_), .A3(new_n554_), .A4(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n545_), .B(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G127gat), .B(G155gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT16), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT69), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n579_), .A3(KEYINPUT17), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n573_), .A2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n580_), .B1(KEYINPUT17), .B2(new_n578_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n573_), .A2(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n542_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n568_), .A2(new_n579_), .A3(new_n571_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n588_), .A2(KEYINPUT12), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT70), .ZN(new_n590_));
  INV_X1    g389(.A(new_n571_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n569_), .A2(new_n570_), .B1(new_n551_), .B2(new_n554_), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT69), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n589_), .A2(new_n590_), .A3(new_n509_), .A4(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n593_), .A2(new_n509_), .A3(KEYINPUT12), .A4(new_n588_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT70), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT12), .B1(new_n509_), .B2(new_n572_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n509_), .A2(new_n572_), .ZN(new_n599_));
  AND2_X1   g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n594_), .A2(new_n596_), .A3(new_n598_), .A4(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT71), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n588_), .A2(KEYINPUT12), .ZN(new_n605_));
  INV_X1    g404(.A(new_n487_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n498_), .A2(new_n472_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT8), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n502_), .A2(new_n503_), .A3(KEYINPUT65), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n506_), .B1(new_n505_), .B2(new_n486_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n500_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n606_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n579_), .B1(new_n568_), .B2(new_n571_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n605_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n597_), .B1(new_n614_), .B2(new_n590_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n615_), .A2(KEYINPUT71), .A3(new_n596_), .A4(new_n601_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n599_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n509_), .A2(new_n572_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n600_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n604_), .A2(new_n616_), .A3(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT5), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n623_), .B(new_n624_), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n625_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n604_), .A2(new_n616_), .A3(new_n620_), .A4(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT13), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n626_), .A2(KEYINPUT13), .A3(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n587_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n471_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT105), .ZN(new_n636_));
  INV_X1    g435(.A(new_n301_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n471_), .A2(new_n638_), .A3(new_n634_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n636_), .A2(new_n637_), .A3(new_n433_), .A4(new_n639_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(KEYINPUT106), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(KEYINPUT106), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n418_), .A2(new_n534_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n633_), .A2(new_n470_), .A3(new_n585_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n648_), .B2(new_n301_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n641_), .A2(new_n642_), .A3(KEYINPUT38), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n645_), .A2(new_n649_), .A3(new_n650_), .ZN(G1324gat));
  INV_X1    g450(.A(new_n418_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n534_), .ZN(new_n653_));
  AND4_X1   g452(.A1(new_n362_), .A2(new_n652_), .A3(new_n653_), .A4(new_n647_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n434_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  INV_X1    g456(.A(new_n362_), .ZN(new_n658_));
  OAI21_X1  g457(.A(KEYINPUT107), .B1(new_n648_), .B2(new_n658_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n656_), .A2(new_n657_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n657_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n636_), .A2(new_n639_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n362_), .A2(new_n434_), .ZN(new_n663_));
  OAI22_X1  g462(.A1(new_n660_), .A2(new_n661_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OAI221_X1 g465(.A(KEYINPUT40), .B1(new_n662_), .B2(new_n663_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1325gat));
  OAI21_X1  g467(.A(G15gat), .B1(new_n648_), .B2(new_n417_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n670_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n417_), .A2(G15gat), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n671_), .B(new_n672_), .C1(new_n662_), .C2(new_n673_), .ZN(G1326gat));
  OAI21_X1  g473(.A(G22gat), .B1(new_n648_), .B2(new_n413_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT42), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n413_), .A2(G22gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n662_), .B2(new_n677_), .ZN(G1327gat));
  NOR3_X1   g477(.A1(new_n633_), .A2(new_n586_), .A3(new_n653_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n471_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G29gat), .B1(new_n681_), .B2(new_n637_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT43), .B1(new_n418_), .B2(new_n542_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n536_), .A2(new_n541_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n417_), .ZN(new_n686_));
  AOI22_X1  g485(.A1(new_n392_), .A2(new_n393_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n687_), .B2(new_n415_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n684_), .B(new_n685_), .C1(new_n688_), .C2(new_n389_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n683_), .A2(new_n689_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n633_), .A2(new_n470_), .A3(new_n586_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n690_), .A2(KEYINPUT44), .A3(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT44), .B1(new_n690_), .B2(new_n691_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n637_), .A2(G29gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n682_), .B1(new_n694_), .B2(new_n695_), .ZN(G1328gat));
  INV_X1    g495(.A(G36gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n362_), .A2(new_n697_), .ZN(new_n698_));
  OR3_X1    g497(.A1(new_n680_), .A2(KEYINPUT45), .A3(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT45), .B1(new_n680_), .B2(new_n698_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n692_), .A2(new_n693_), .A3(new_n658_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(new_n697_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n701_), .B(KEYINPUT46), .C1(new_n702_), .C2(new_n697_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  AOI21_X1  g506(.A(G43gat), .B1(new_n681_), .B2(new_n686_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n686_), .A2(G43gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n694_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(G1330gat));
  AOI21_X1  g511(.A(G50gat), .B1(new_n681_), .B2(new_n388_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n388_), .A2(G50gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n694_), .B2(new_n714_), .ZN(G1331gat));
  NOR2_X1   g514(.A1(new_n418_), .A2(new_n469_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n633_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n587_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n548_), .B1(new_n719_), .B2(new_n301_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n469_), .A2(new_n585_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n646_), .A2(new_n633_), .A3(new_n721_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n722_), .A2(new_n548_), .A3(new_n301_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n723_), .B2(KEYINPUT109), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(KEYINPUT109), .B2(new_n723_), .ZN(G1332gat));
  OAI21_X1  g524(.A(G64gat), .B1(new_n722_), .B2(new_n658_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT48), .ZN(new_n727_));
  INV_X1    g526(.A(new_n719_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(new_n546_), .A3(new_n362_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1333gat));
  OAI21_X1  g529(.A(G71gat), .B1(new_n722_), .B2(new_n417_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT49), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n728_), .A2(new_n203_), .A3(new_n686_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1334gat));
  OAI21_X1  g533(.A(G78gat), .B1(new_n722_), .B2(new_n413_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT50), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n728_), .A2(new_n378_), .A3(new_n388_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1335gat));
  NOR2_X1   g537(.A1(new_n653_), .A2(new_n586_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n716_), .A2(new_n633_), .A3(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n476_), .B1(new_n740_), .B2(new_n301_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT110), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n633_), .A2(new_n470_), .A3(new_n585_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n683_), .B2(new_n689_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n745_), .A2(new_n476_), .A3(new_n301_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n742_), .A2(new_n746_), .ZN(G1336gat));
  OAI21_X1  g546(.A(G92gat), .B1(new_n745_), .B2(new_n658_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n740_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(new_n477_), .A3(new_n362_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1337gat));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(KEYINPUT51), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n686_), .A2(new_n474_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n745_), .A2(new_n417_), .ZN(new_n756_));
  OAI221_X1 g555(.A(new_n754_), .B1(new_n740_), .B2(new_n755_), .C1(new_n756_), .C2(new_n495_), .ZN(new_n757_));
  OAI22_X1  g556(.A1(new_n756_), .A2(new_n495_), .B1(new_n740_), .B2(new_n755_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n752_), .B2(KEYINPUT51), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n757_), .B1(new_n759_), .B2(new_n754_), .ZN(G1338gat));
  OAI211_X1 g559(.A(KEYINPUT113), .B(G106gat), .C1(new_n745_), .C2(new_n413_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762_));
  AOI211_X1 g561(.A(new_n413_), .B(new_n743_), .C1(new_n683_), .C2(new_n689_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n380_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n761_), .A2(new_n764_), .A3(KEYINPUT52), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n762_), .B(new_n766_), .C1(new_n763_), .C2(new_n380_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n749_), .A2(new_n380_), .A3(new_n388_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT53), .B1(new_n765_), .B2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n761_), .A2(new_n764_), .A3(KEYINPUT52), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n767_), .A4(new_n768_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(new_n773_), .ZN(G1339gat));
  NOR4_X1   g573(.A1(new_n362_), .A2(new_n388_), .A3(new_n301_), .A4(new_n417_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n469_), .A2(new_n776_), .A3(new_n628_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n469_), .B2(new_n628_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n604_), .A2(new_n616_), .A3(new_n780_), .ZN(new_n781_));
  AND4_X1   g580(.A1(new_n596_), .A2(new_n594_), .A3(new_n598_), .A4(new_n601_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n594_), .A2(new_n596_), .A3(new_n617_), .A4(new_n598_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n782_), .A2(KEYINPUT55), .B1(new_n783_), .B2(new_n600_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT118), .B1(new_n786_), .B2(KEYINPUT117), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n625_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n627_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(KEYINPUT117), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n788_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n789_), .B2(KEYINPUT56), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n779_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n446_), .A2(new_n447_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT119), .B1(new_n795_), .B2(new_n468_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n458_), .A2(new_n462_), .A3(new_n448_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(KEYINPUT119), .A3(new_n468_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n449_), .A2(new_n463_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n798_), .A2(new_n799_), .B1(new_n421_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n629_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n794_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n534_), .A2(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n801_), .A2(new_n628_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n789_), .A2(KEYINPUT56), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n786_), .B(new_n627_), .C1(new_n781_), .C2(new_n784_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n806_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n542_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n806_), .B(KEYINPUT58), .C1(new_n807_), .C2(new_n808_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n803_), .A2(new_n805_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n802_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n789_), .A2(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT118), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n789_), .A2(new_n790_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n788_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n814_), .B1(new_n818_), .B2(new_n779_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n804_), .B1(new_n819_), .B2(new_n534_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n586_), .B1(new_n813_), .B2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n631_), .A2(new_n632_), .A3(new_n721_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT114), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n631_), .A2(new_n824_), .A3(new_n632_), .A4(new_n721_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n542_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n828_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n826_), .A2(new_n542_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n775_), .B1(new_n821_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(G113gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(new_n469_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n833_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n809_), .A2(new_n810_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n685_), .A3(new_n812_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n805_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n819_), .B2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT57), .B1(new_n803_), .B2(new_n653_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n585_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n830_), .B1(new_n826_), .B2(new_n542_), .ZN(new_n845_));
  AOI211_X1 g644(.A(new_n685_), .B(new_n828_), .C1(new_n823_), .C2(new_n825_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n844_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(KEYINPUT59), .A3(new_n775_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n470_), .B1(new_n838_), .B2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n836_), .B1(new_n850_), .B2(new_n835_), .ZN(G1340gat));
  NOR2_X1   g650(.A1(new_n717_), .A2(KEYINPUT60), .ZN(new_n852_));
  MUX2_X1   g651(.A(new_n852_), .B(KEYINPUT60), .S(G120gat), .Z(new_n853_));
  NAND2_X1  g652(.A1(new_n834_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n717_), .B1(new_n838_), .B2(new_n849_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G120gat), .B1(new_n855_), .B2(KEYINPUT120), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857_));
  AOI211_X1 g656(.A(new_n857_), .B(new_n717_), .C1(new_n838_), .C2(new_n849_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n854_), .B1(new_n856_), .B2(new_n858_), .ZN(G1341gat));
  INV_X1    g658(.A(G127gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n834_), .A2(new_n860_), .A3(new_n586_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n585_), .B1(new_n838_), .B2(new_n849_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n860_), .ZN(G1342gat));
  INV_X1    g662(.A(G134gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n834_), .A2(new_n864_), .A3(new_n534_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n542_), .B1(new_n838_), .B2(new_n849_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n864_), .ZN(G1343gat));
  NOR2_X1   g666(.A1(new_n821_), .A2(new_n832_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n658_), .A2(new_n388_), .A3(new_n637_), .A4(new_n417_), .ZN(new_n869_));
  XOR2_X1   g668(.A(new_n869_), .B(KEYINPUT121), .Z(new_n870_));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n469_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT122), .B(G141gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1344gat));
  NAND2_X1  g673(.A1(new_n871_), .A2(new_n633_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g675(.A1(new_n871_), .A2(new_n586_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G155gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  INV_X1    g678(.A(G162gat), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n868_), .A2(new_n880_), .A3(new_n542_), .A4(new_n870_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n871_), .A2(new_n534_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n880_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n882_), .A2(KEYINPUT123), .A3(new_n880_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n881_), .B1(new_n885_), .B2(new_n886_), .ZN(G1347gat));
  NOR2_X1   g686(.A1(new_n658_), .A2(new_n303_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(KEYINPUT124), .Z(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n388_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n848_), .A2(new_n469_), .A3(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT62), .B1(new_n891_), .B2(KEYINPUT22), .ZN(new_n892_));
  OAI21_X1  g691(.A(G169gat), .B1(new_n891_), .B2(KEYINPUT62), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n894_), .B1(new_n209_), .B2(new_n892_), .ZN(G1348gat));
  NAND2_X1  g694(.A1(new_n848_), .A2(new_n890_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n717_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n210_), .ZN(G1349gat));
  INV_X1    g697(.A(new_n896_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n223_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n900_), .A3(new_n586_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902_));
  INV_X1    g701(.A(G183gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n896_), .B2(new_n585_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n901_), .A2(new_n902_), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n902_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n896_), .B2(new_n542_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n534_), .A2(new_n224_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n896_), .B2(new_n909_), .ZN(G1351gat));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n362_), .A2(new_n417_), .A3(new_n391_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n911_), .B1(new_n848_), .B2(new_n913_), .ZN(new_n914_));
  AOI211_X1 g713(.A(KEYINPUT126), .B(new_n912_), .C1(new_n844_), .C2(new_n847_), .ZN(new_n915_));
  OAI211_X1 g714(.A(G197gat), .B(new_n469_), .C1(new_n914_), .C2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n469_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n310_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n913_), .B1(new_n821_), .B2(new_n832_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(KEYINPUT126), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n848_), .A2(new_n911_), .A3(new_n913_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n924_), .A2(KEYINPUT127), .A3(G197gat), .A4(new_n469_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n918_), .A2(new_n920_), .A3(new_n925_), .ZN(G1352gat));
  AOI21_X1  g725(.A(new_n717_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(new_n312_), .ZN(G1353gat));
  OR2_X1    g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  AND4_X1   g729(.A1(new_n586_), .A2(new_n924_), .A3(new_n929_), .A4(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n929_), .B1(new_n924_), .B2(new_n586_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1354gat));
  INV_X1    g732(.A(G218gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n924_), .A2(new_n934_), .A3(new_n534_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n542_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n936_), .B2(new_n934_), .ZN(G1355gat));
endmodule


