//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT87), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G197gat), .B(G204gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT21), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT85), .ZN(new_n209_));
  INV_X1    g008(.A(G197gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n209_), .B1(new_n210_), .B2(G204gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT86), .ZN(new_n212_));
  INV_X1    g011(.A(G204gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n212_), .B1(new_n213_), .B2(G197gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n210_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n211_), .A2(new_n214_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT21), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n205_), .B(new_n218_), .C1(KEYINPUT21), .C2(new_n206_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n208_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT23), .ZN(new_n222_));
  OR3_X1    g021(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT93), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n227_), .A2(new_n228_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n222_), .A2(KEYINPUT93), .A3(new_n223_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n226_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n222_), .B1(G183gat), .B2(G190gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n231_), .B(KEYINPUT77), .Z(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT22), .B(G169gat), .Z(new_n237_));
  OAI211_X1 g036(.A(new_n235_), .B(new_n236_), .C1(G176gat), .C2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n202_), .B1(new_n220_), .B2(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n224_), .A2(KEYINPUT78), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(new_n230_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n224_), .A2(KEYINPUT78), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT76), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G190gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n245_), .B(KEYINPUT26), .Z(new_n246_));
  OR2_X1    g045(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT75), .B(G183gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .A4(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n248_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n222_), .B1(new_n253_), .B2(G190gat), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT79), .B(KEYINPUT22), .Z(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT80), .A3(G169gat), .ZN(new_n256_));
  INV_X1    g055(.A(G176gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(G169gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT22), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n255_), .A2(G169gat), .B1(KEYINPUT80), .B2(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n236_), .B(new_n254_), .C1(new_n258_), .C2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n252_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n240_), .B1(new_n220_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G226gat), .A2(G233gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT19), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n208_), .A2(new_n219_), .A3(new_n234_), .A4(new_n238_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n268_), .A2(KEYINPUT94), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n202_), .B1(new_n268_), .B2(KEYINPUT94), .ZN(new_n270_));
  INV_X1    g069(.A(new_n266_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n263_), .A2(new_n220_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .A4(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G8gat), .B(G36gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT96), .ZN(new_n275_));
  XOR2_X1   g074(.A(G64gat), .B(G92gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n267_), .A2(new_n273_), .A3(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n264_), .A2(new_n266_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n268_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT101), .B1(new_n283_), .B2(new_n202_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT101), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n268_), .A2(new_n285_), .A3(KEYINPUT20), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n286_), .A3(new_n272_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n282_), .B1(new_n266_), .B2(new_n287_), .ZN(new_n288_));
  OAI211_X1 g087(.A(KEYINPUT27), .B(new_n281_), .C1(new_n288_), .C2(new_n280_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT27), .ZN(new_n290_));
  INV_X1    g089(.A(new_n281_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n280_), .B1(new_n267_), .B2(new_n273_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G78gat), .B(G106gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT88), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT89), .ZN(new_n297_));
  OR2_X1    g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT3), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT84), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n298_), .A2(new_n300_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n301_), .A2(new_n304_), .A3(new_n305_), .A4(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n307_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT82), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n313_), .B1(G155gat), .B2(G162gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n312_), .B1(new_n314_), .B2(new_n309_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n308_), .A2(KEYINPUT1), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n310_), .A2(new_n316_), .A3(KEYINPUT82), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(G155gat), .A3(G162gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n298_), .A2(new_n302_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n319_), .A2(KEYINPUT83), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT83), .B1(new_n319_), .B2(new_n320_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n311_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT29), .ZN(new_n324_));
  INV_X1    g123(.A(G228gat), .ZN(new_n325_));
  INV_X1    g124(.A(G233gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(new_n328_), .A3(new_n220_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n324_), .B2(new_n220_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n297_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n307_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n319_), .A2(new_n320_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT83), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n319_), .A2(KEYINPUT83), .A3(new_n320_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n333_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n220_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n327_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n297_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n329_), .A3(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n332_), .A2(new_n343_), .A3(KEYINPUT90), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n343_), .A2(KEYINPUT90), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G22gat), .B(G50gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT28), .B1(new_n323_), .B2(KEYINPUT29), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n323_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n347_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n350_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(new_n348_), .A3(new_n346_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n344_), .A2(new_n345_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT91), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n356_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n341_), .A2(KEYINPUT91), .A3(new_n329_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(new_n358_), .A3(new_n296_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n343_), .A2(new_n353_), .A3(new_n351_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT92), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n359_), .A2(new_n360_), .A3(KEYINPUT92), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n294_), .B(new_n355_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G127gat), .B(G134gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G113gat), .B(G120gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT31), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n263_), .B(KEYINPUT30), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT81), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G227gat), .A2(G233gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G15gat), .ZN(new_n371_));
  INV_X1    g170(.A(G43gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G71gat), .B(G99gat), .Z(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n369_), .A2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n376_), .B1(new_n368_), .B2(KEYINPUT81), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n367_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n367_), .ZN(new_n381_));
  AOI211_X1 g180(.A(new_n378_), .B(new_n381_), .C1(new_n369_), .C2(new_n376_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G85gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT0), .B(G57gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  INV_X1    g186(.A(new_n366_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n323_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n311_), .B(new_n366_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT98), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT98), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n389_), .A2(new_n394_), .A3(new_n390_), .A4(new_n391_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT97), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(new_n389_), .B2(KEYINPUT4), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n389_), .A2(KEYINPUT4), .A3(new_n391_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n390_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n323_), .A2(KEYINPUT97), .A3(new_n401_), .A4(new_n388_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .A4(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n387_), .B1(new_n396_), .B2(new_n403_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n403_), .A2(new_n387_), .A3(new_n395_), .A4(new_n393_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT102), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n387_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n403_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n393_), .A2(new_n395_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT102), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n405_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n383_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n363_), .A2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n355_), .B1(new_n362_), .B2(new_n361_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(new_n414_), .A3(new_n294_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n267_), .A2(new_n273_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n279_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n281_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n405_), .A2(KEYINPUT33), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n396_), .A2(new_n423_), .A3(new_n387_), .A4(new_n403_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n398_), .A2(new_n399_), .A3(new_n390_), .A4(new_n402_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n389_), .A2(new_n400_), .A3(new_n391_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n408_), .A3(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT99), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n280_), .A2(KEYINPUT100), .A3(KEYINPUT32), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT100), .B1(new_n280_), .B2(KEYINPUT32), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n419_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n411_), .A2(new_n405_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT32), .ZN(new_n435_));
  OR3_X1    g234(.A1(new_n288_), .A2(new_n435_), .A3(new_n279_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n425_), .A2(new_n429_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n418_), .B1(new_n417_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n383_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n416_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT13), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT68), .ZN(new_n442_));
  AND2_X1   g241(.A1(G85gat), .A2(G92gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(G85gat), .A2(G92gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT9), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n445_), .A2(G85gat), .A3(G92gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n446_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(G99gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT10), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT10), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(G99gat), .ZN(new_n457_));
  AOI211_X1 g256(.A(KEYINPUT64), .B(G106gat), .C1(new_n455_), .C2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT64), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n457_), .ZN(new_n460_));
  INV_X1    g259(.A(G106gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n453_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT7), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(new_n454_), .A3(new_n461_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n465_), .A2(new_n449_), .A3(new_n451_), .A4(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n443_), .A2(new_n444_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT8), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(KEYINPUT65), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(KEYINPUT65), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT65), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT8), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n467_), .A2(new_n468_), .A3(new_n472_), .A4(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n463_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(G71gat), .A2(G78gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G71gat), .A2(G78gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(G57gat), .A2(G64gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(G57gat), .A2(G64gat), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n481_), .A2(new_n482_), .A3(KEYINPUT11), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT11), .ZN(new_n484_));
  INV_X1    g283(.A(G57gat), .ZN(new_n485_));
  INV_X1    g284(.A(G64gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G57gat), .A2(G64gat), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n484_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n480_), .B1(new_n483_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT11), .B1(new_n481_), .B2(new_n482_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n479_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n476_), .A2(KEYINPUT12), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT66), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n490_), .A2(new_n495_), .A3(new_n492_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n487_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n479_), .B1(new_n491_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n487_), .A2(new_n488_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n499_), .A2(KEYINPUT11), .B1(new_n477_), .B2(new_n478_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT66), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n496_), .A2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT12), .B1(new_n476_), .B2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n494_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT67), .ZN(new_n505_));
  AOI211_X1 g304(.A(new_n473_), .B(KEYINPUT8), .C1(new_n467_), .C2(new_n468_), .ZN(new_n506_));
  AND4_X1   g305(.A1(new_n468_), .A2(new_n467_), .A3(new_n472_), .A4(new_n474_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n508_), .A2(new_n463_), .A3(new_n501_), .A4(new_n496_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G230gat), .A2(G233gat), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n505_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n505_), .B(new_n510_), .C1(new_n476_), .C2(new_n502_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n504_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n476_), .A2(new_n502_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n509_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n510_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT5), .B(G176gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(G204gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G120gat), .B(G148gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  OAI21_X1  g322(.A(new_n442_), .B1(new_n519_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n523_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n514_), .A2(KEYINPUT68), .A3(new_n518_), .A4(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n519_), .A2(new_n523_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n441_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(new_n441_), .A3(new_n528_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT73), .B(G15gat), .ZN(new_n533_));
  INV_X1    g332(.A(G22gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(G1gat), .ZN(new_n536_));
  INV_X1    g335(.A(G8gat), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT14), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G1gat), .B(G8gat), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n540_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G29gat), .B(G36gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n541_), .A2(new_n542_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT15), .ZN(new_n550_));
  INV_X1    g349(.A(new_n544_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n551_), .A2(new_n545_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n545_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n550_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(KEYINPUT15), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n549_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n547_), .A2(new_n548_), .A3(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n549_), .B(new_n546_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n558_), .B1(new_n559_), .B2(new_n548_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT74), .B(G169gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(G197gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G113gat), .B(G141gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n565_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n558_), .B(new_n564_), .C1(new_n559_), .C2(new_n548_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n532_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n440_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n556_), .A2(new_n476_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT34), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT35), .Z(new_n574_));
  NAND4_X1  g373(.A1(new_n463_), .A2(new_n471_), .A3(new_n546_), .A4(new_n475_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n571_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(KEYINPUT35), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n577_), .B1(new_n571_), .B2(new_n575_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT70), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n576_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n571_), .A2(KEYINPUT70), .A3(new_n574_), .A4(new_n575_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G134gat), .B(G162gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(G218gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT69), .B(G190gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT36), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n582_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n586_), .A2(KEYINPUT36), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n580_), .A2(new_n581_), .A3(new_n589_), .ZN(new_n590_));
  AND4_X1   g389(.A1(KEYINPUT71), .A2(new_n590_), .A3(KEYINPUT72), .A4(KEYINPUT37), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(KEYINPUT71), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n588_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(KEYINPUT72), .B(new_n590_), .C1(new_n582_), .C2(new_n587_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT37), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(G231gat), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(new_n326_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n543_), .A2(new_n599_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n549_), .A2(new_n598_), .A3(new_n326_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(new_n493_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(G211gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT16), .B(G183gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(KEYINPUT17), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n490_), .B(new_n492_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n603_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n607_), .B(KEYINPUT17), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n602_), .A2(new_n502_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n501_), .B(new_n496_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n597_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n570_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n414_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n536_), .A3(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT38), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n588_), .A2(new_n590_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n616_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n570_), .A2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G1gat), .B1(new_n625_), .B2(new_n414_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n621_), .A2(new_n626_), .ZN(G1324gat));
  INV_X1    g426(.A(new_n294_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n618_), .A2(new_n537_), .A3(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n570_), .A2(new_n628_), .A3(new_n624_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(new_n631_), .A3(G8gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n631_), .B1(new_n630_), .B2(G8gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n629_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g435(.A(G15gat), .B1(new_n625_), .B2(new_n439_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT41), .Z(new_n638_));
  INV_X1    g437(.A(G15gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n618_), .A2(new_n639_), .A3(new_n383_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(G1326gat));
  INV_X1    g440(.A(new_n417_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G22gat), .B1(new_n625_), .B2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n618_), .A2(new_n534_), .A3(new_n417_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1327gat));
  NAND2_X1  g446(.A1(new_n438_), .A2(new_n439_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n416_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n615_), .A2(new_n622_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n650_), .A2(new_n568_), .A3(new_n532_), .A4(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n619_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n597_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT43), .B1(new_n440_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n425_), .A2(new_n429_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n434_), .A2(new_n436_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n642_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n383_), .B1(new_n660_), .B2(new_n418_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n657_), .B(new_n597_), .C1(new_n661_), .C2(new_n416_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n656_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n532_), .A2(new_n568_), .A3(new_n616_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT44), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  AOI211_X1 g466(.A(new_n667_), .B(new_n664_), .C1(new_n656_), .C2(new_n662_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(G29gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n654_), .B1(new_n670_), .B2(new_n619_), .ZN(G1328gat));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  INV_X1    g471(.A(G36gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n669_), .B2(new_n628_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT45), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n652_), .A2(G36gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(new_n628_), .ZN(new_n677_));
  NOR4_X1   g476(.A1(new_n652_), .A2(KEYINPUT45), .A3(G36gat), .A4(new_n294_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n672_), .B1(new_n674_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n679_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n666_), .A2(new_n668_), .A3(new_n294_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n681_), .B(KEYINPUT46), .C1(new_n673_), .C2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1329gat));
  INV_X1    g483(.A(new_n666_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n663_), .A2(KEYINPUT44), .A3(new_n665_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n685_), .A2(G43gat), .A3(new_n383_), .A4(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n372_), .B1(new_n652_), .B2(new_n439_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT47), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT47), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n687_), .A2(new_n691_), .A3(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1330gat));
  AOI21_X1  g492(.A(G50gat), .B1(new_n653_), .B2(new_n417_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n417_), .A2(G50gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n669_), .B2(new_n695_), .ZN(G1331gat));
  OR3_X1    g495(.A1(new_n440_), .A2(KEYINPUT104), .A3(new_n568_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT104), .B1(new_n440_), .B2(new_n568_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n527_), .A2(new_n441_), .A3(new_n528_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(new_n529_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n619_), .A3(new_n617_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n568_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n701_), .A2(new_n624_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n650_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT105), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n650_), .A2(new_n708_), .A3(new_n704_), .A4(new_n705_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n707_), .A2(G57gat), .A3(new_n709_), .ZN(new_n710_));
  AOI22_X1  g509(.A1(new_n703_), .A2(new_n485_), .B1(new_n619_), .B2(new_n710_), .ZN(G1332gat));
  NAND2_X1  g510(.A1(new_n702_), .A2(new_n617_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n628_), .A2(new_n486_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n707_), .A2(new_n709_), .A3(new_n628_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT106), .B(KEYINPUT48), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(G64gat), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n714_), .B2(G64gat), .ZN(new_n717_));
  OAI22_X1  g516(.A1(new_n712_), .A2(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(G1333gat));
  OR2_X1    g517(.A1(new_n439_), .A2(G71gat), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT49), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n707_), .A2(new_n709_), .A3(new_n383_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(G71gat), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n721_), .A2(new_n720_), .A3(G71gat), .ZN(new_n723_));
  OAI22_X1  g522(.A1(new_n712_), .A2(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1334gat));
  NOR2_X1   g523(.A1(new_n642_), .A2(G78gat), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n699_), .A2(new_n701_), .A3(new_n617_), .A4(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n707_), .A2(new_n709_), .A3(new_n417_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(G78gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G78gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT107), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n733_), .B(new_n726_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1335gat));
  NAND4_X1  g534(.A1(new_n697_), .A2(new_n701_), .A3(new_n651_), .A4(new_n698_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G85gat), .B1(new_n737_), .B2(new_n619_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n532_), .A2(new_n568_), .A3(new_n615_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n656_), .B2(new_n662_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT108), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n619_), .A2(G85gat), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT109), .Z(new_n744_));
  AOI21_X1  g543(.A(new_n738_), .B1(new_n742_), .B2(new_n744_), .ZN(G1336gat));
  AOI21_X1  g544(.A(G92gat), .B1(new_n737_), .B2(new_n628_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n742_), .A2(new_n628_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(G92gat), .ZN(G1337gat));
  NAND2_X1  g547(.A1(new_n383_), .A2(new_n460_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n736_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n741_), .A2(new_n383_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(G99gat), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n754_), .A2(KEYINPUT51), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(KEYINPUT51), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n750_), .A2(new_n754_), .A3(KEYINPUT51), .A4(new_n752_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1338gat));
  NAND3_X1  g558(.A1(new_n737_), .A2(new_n461_), .A3(new_n417_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n741_), .A2(new_n417_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(G106gat), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT52), .B(new_n461_), .C1(new_n741_), .C2(new_n417_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n760_), .B(new_n766_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1339gat));
  NOR3_X1   g569(.A1(new_n363_), .A2(new_n439_), .A3(new_n414_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT12), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n515_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n476_), .A2(KEYINPUT12), .A3(new_n493_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n509_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT114), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n774_), .A2(new_n778_), .A3(new_n509_), .A4(new_n775_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n777_), .A2(new_n517_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n514_), .A2(new_n781_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n504_), .B(KEYINPUT55), .C1(new_n511_), .C2(new_n513_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n780_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(KEYINPUT56), .A3(new_n523_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT56), .B1(new_n784_), .B2(new_n523_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n568_), .B(new_n527_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n543_), .A2(new_n546_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n549_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n548_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n547_), .A2(new_n557_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n791_), .B(new_n565_), .C1(new_n548_), .C2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n567_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n788_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT57), .B1(new_n797_), .B2(new_n622_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n799_));
  AOI211_X1 g598(.A(new_n799_), .B(new_n623_), .C1(new_n788_), .C2(new_n796_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n786_), .A2(new_n787_), .A3(KEYINPUT115), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n784_), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n523_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n793_), .A2(new_n567_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n804_), .A3(new_n527_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT116), .B1(new_n802_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n803_), .A2(new_n804_), .A3(new_n527_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n784_), .A2(new_n523_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n813_), .A3(new_n785_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n809_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(KEYINPUT116), .A3(KEYINPUT58), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n655_), .B1(new_n808_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n801_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT58), .B1(new_n815_), .B2(KEYINPUT116), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n821_), .B(new_n807_), .C1(new_n809_), .C2(new_n814_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n597_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(KEYINPUT117), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n616_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n593_), .A2(new_n615_), .A3(new_n596_), .A4(new_n704_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT112), .B1(new_n701_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n701_), .A2(new_n826_), .A3(KEYINPUT112), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n830_), .A2(new_n831_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n835_));
  INV_X1    g634(.A(new_n826_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n532_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT113), .B1(new_n837_), .B2(KEYINPUT54), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n832_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n834_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n772_), .B1(new_n825_), .B2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(G113gat), .B1(new_n842_), .B2(new_n568_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n704_), .B1(new_n812_), .B2(new_n785_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n795_), .B1(new_n844_), .B2(new_n527_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n799_), .B1(new_n845_), .B2(new_n623_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n797_), .A2(KEYINPUT57), .A3(new_n622_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n616_), .B1(new_n817_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT119), .B(new_n616_), .C1(new_n817_), .C2(new_n848_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n841_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n772_), .A2(KEYINPUT118), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n772_), .A2(KEYINPUT118), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT59), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n842_), .A2(KEYINPUT59), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n704_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n843_), .B1(new_n860_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g660(.A(G120gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n532_), .B2(KEYINPUT60), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n842_), .B(new_n863_), .C1(KEYINPUT60), .C2(new_n862_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n532_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n862_), .ZN(G1341gat));
  AOI21_X1  g665(.A(G127gat), .B1(new_n842_), .B2(new_n615_), .ZN(new_n867_));
  INV_X1    g666(.A(G127gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n869_), .B2(new_n615_), .ZN(G1342gat));
  AOI21_X1  g669(.A(G134gat), .B1(new_n842_), .B2(new_n623_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n655_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g672(.A1(new_n642_), .A2(new_n628_), .A3(new_n414_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n848_), .B1(KEYINPUT117), .B2(new_n823_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n817_), .A2(new_n818_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n615_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n833_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n838_), .A2(new_n832_), .A3(new_n839_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n439_), .B(new_n874_), .C1(new_n877_), .C2(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n704_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT120), .B(G141gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1344gat));
  NOR2_X1   g683(.A1(new_n881_), .A2(new_n532_), .ZN(new_n885_));
  XOR2_X1   g684(.A(new_n885_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g685(.A1(new_n881_), .A2(new_n616_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT61), .B(G155gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  OAI21_X1  g688(.A(G162gat), .B1(new_n881_), .B2(new_n655_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n383_), .B1(new_n825_), .B2(new_n841_), .ZN(new_n892_));
  INV_X1    g691(.A(G162gat), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n892_), .A2(new_n893_), .A3(new_n623_), .A4(new_n874_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n890_), .A2(new_n891_), .A3(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n891_), .B1(new_n890_), .B2(new_n894_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n415_), .A2(new_n294_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n853_), .A2(new_n568_), .A3(new_n642_), .A4(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G169gat), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n899_), .A2(G169gat), .A3(new_n901_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n903_), .B(new_n904_), .C1(new_n237_), .C2(new_n899_), .ZN(G1348gat));
  AND2_X1   g704(.A1(new_n853_), .A2(new_n642_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n906_), .A2(new_n701_), .A3(new_n898_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n417_), .B1(new_n825_), .B2(new_n841_), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n908_), .A2(G176gat), .A3(new_n701_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n907_), .A2(new_n257_), .B1(new_n898_), .B2(new_n909_), .ZN(G1349gat));
  NAND3_X1  g709(.A1(new_n908_), .A2(new_n615_), .A3(new_n898_), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n415_), .A2(new_n227_), .A3(new_n294_), .A4(new_n616_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n911_), .A2(new_n248_), .B1(new_n906_), .B2(new_n912_), .ZN(G1350gat));
  NAND3_X1  g712(.A1(new_n906_), .A2(new_n597_), .A3(new_n898_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(G190gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n623_), .A2(new_n228_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT123), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n906_), .A2(new_n898_), .A3(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n915_), .A2(new_n918_), .ZN(G1351gat));
  NOR3_X1   g718(.A1(new_n642_), .A2(new_n619_), .A3(new_n294_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n892_), .A2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n704_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(new_n210_), .ZN(G1352gat));
  NOR2_X1   g722(.A1(new_n921_), .A2(new_n532_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT124), .B(G204gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n924_), .B(new_n925_), .ZN(G1353gat));
  NAND3_X1  g725(.A1(new_n892_), .A2(new_n615_), .A3(new_n920_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT63), .ZN(new_n929_));
  INV_X1    g728(.A(G211gat), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n928_), .A2(KEYINPUT125), .A3(new_n929_), .A4(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n929_), .A2(new_n930_), .A3(KEYINPUT125), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n933_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n929_), .A2(new_n930_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n932_), .B(new_n934_), .C1(new_n927_), .C2(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n931_), .A2(new_n936_), .ZN(G1354gat));
  XNOR2_X1  g736(.A(KEYINPUT126), .B(G218gat), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n921_), .A2(new_n655_), .A3(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n921_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n623_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n942_), .B2(new_n939_), .ZN(G1355gat));
endmodule


