//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  OR3_X1    g001(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n204_));
  AOI22_X1  g003(.A1(new_n203_), .A2(new_n204_), .B1(G155gat), .B2(G162gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n206_));
  NOR3_X1   g005(.A1(new_n206_), .A2(G141gat), .A3(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(G141gat), .ZN(new_n208_));
  INV_X1    g007(.A(G148gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT3), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  OAI22_X1  g011(.A1(new_n207_), .A2(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT83), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT83), .A2(G141gat), .A3(G148gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT2), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n205_), .B1(new_n213_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n216_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n208_), .A2(new_n209_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n204_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G155gat), .ZN(new_n224_));
  INV_X1    g023(.A(G162gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT1), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(G155gat), .A3(G162gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n219_), .B(new_n220_), .C1(new_n223_), .C2(new_n229_), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n218_), .A2(KEYINPUT85), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT85), .B1(new_n218_), .B2(new_n230_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(KEYINPUT29), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G22gat), .B(G50gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n234_), .B(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G78gat), .B(G106gat), .Z(new_n239_));
  NAND2_X1  g038(.A1(new_n233_), .A2(KEYINPUT29), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G228gat), .A2(G233gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT87), .ZN(new_n242_));
  XOR2_X1   g041(.A(G197gat), .B(G204gat), .Z(new_n243_));
  XNOR2_X1  g042(.A(G211gat), .B(G218gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT88), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n243_), .A2(KEYINPUT21), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n244_), .B1(new_n243_), .B2(KEYINPUT21), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n240_), .A2(new_n242_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n242_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n218_), .A2(new_n230_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT29), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n251_), .B1(new_n254_), .B2(new_n248_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n239_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT89), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n238_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n250_), .A2(new_n239_), .A3(new_n255_), .ZN(new_n259_));
  OR3_X1    g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n256_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n256_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT20), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT22), .B(G169gat), .ZN(new_n265_));
  INV_X1    g064(.A(G176gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT79), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n265_), .A2(KEYINPUT79), .A3(new_n266_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT80), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G183gat), .A2(G190gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n274_), .B(KEYINPUT23), .Z(new_n275_));
  NOR2_X1   g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT80), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n269_), .A2(new_n278_), .A3(new_n270_), .A4(new_n271_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n273_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT25), .B(G183gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(G190gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT78), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n287_), .A2(new_n270_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n275_), .B1(KEYINPUT24), .B2(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n285_), .B(new_n289_), .C1(KEYINPUT24), .C2(new_n287_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n280_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n264_), .B1(new_n291_), .B2(new_n248_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G226gat), .A2(G233gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n293_), .B(KEYINPUT90), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT19), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT91), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n282_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n281_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(new_n287_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n275_), .B1(new_n299_), .B2(new_n288_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n298_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT93), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n277_), .A2(new_n267_), .A3(new_n270_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n298_), .A2(KEYINPUT93), .A3(new_n301_), .A4(new_n300_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n249_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n292_), .A2(new_n295_), .A3(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n302_), .A2(new_n248_), .A3(new_n305_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT20), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT98), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n280_), .A2(new_n290_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n249_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(KEYINPUT98), .A3(KEYINPUT20), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n313_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n309_), .B1(new_n295_), .B2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G8gat), .B(G36gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT18), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(G64gat), .ZN(new_n321_));
  INV_X1    g120(.A(G92gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n295_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n308_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT20), .B1(new_n314_), .B2(new_n249_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n326_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n295_), .A2(KEYINPUT20), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n315_), .B(new_n331_), .C1(new_n249_), .C2(new_n307_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(new_n332_), .A3(new_n323_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n325_), .A2(KEYINPUT27), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n295_), .B1(new_n292_), .B2(new_n308_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n332_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n324_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n333_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT101), .B(KEYINPUT27), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G127gat), .B(G134gat), .ZN(new_n342_));
  INV_X1    g141(.A(G113gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G120gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n342_), .B(G113gat), .ZN(new_n346_));
  INV_X1    g145(.A(G120gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n314_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT30), .B(G71gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G15gat), .B(G43gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(G99gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT31), .ZN(new_n356_));
  XOR2_X1   g155(.A(KEYINPUT81), .B(KEYINPUT82), .Z(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  XNOR2_X1  g159(.A(new_n353_), .B(new_n360_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n263_), .A2(new_n341_), .A3(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n349_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT94), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n350_), .A2(new_n252_), .ZN(new_n366_));
  OAI211_X1 g165(.A(KEYINPUT94), .B(new_n349_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT4), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(KEYINPUT95), .Z(new_n371_));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n363_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n369_), .A2(new_n371_), .A3(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G1gat), .B(G29gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G85gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT0), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G57gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n371_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n368_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n374_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT99), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n374_), .A2(new_n380_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n378_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT99), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n374_), .A2(new_n386_), .A3(new_n378_), .A4(new_n380_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n382_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n362_), .A2(new_n389_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n341_), .A2(new_n262_), .A3(new_n388_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n323_), .A2(KEYINPUT32), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n335_), .A2(new_n336_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n393_), .B1(new_n318_), .B2(new_n392_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n388_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT100), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n338_), .B1(new_n385_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT33), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT96), .B1(new_n385_), .B2(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n368_), .A2(new_n379_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n369_), .A2(new_n373_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n402_), .B(new_n378_), .C1(new_n403_), .C2(new_n371_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT96), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n383_), .A2(new_n405_), .A3(KEYINPUT33), .A4(new_n384_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n399_), .A2(new_n401_), .A3(new_n404_), .A4(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n388_), .A2(new_n394_), .A3(KEYINPUT100), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n397_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n391_), .B1(new_n409_), .B2(new_n262_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n361_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n390_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G230gat), .A2(G233gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT64), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G71gat), .B(G78gat), .Z(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G57gat), .B(G64gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT11), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n418_), .A2(KEYINPUT11), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n416_), .A2(KEYINPUT11), .A3(new_n418_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(G85gat), .A2(G92gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G85gat), .A2(G92gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(KEYINPUT68), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT68), .ZN(new_n428_));
  INV_X1    g227(.A(new_n426_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n428_), .B1(new_n429_), .B2(new_n424_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT69), .ZN(new_n432_));
  AND3_X1   g231(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n432_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G99gat), .A2(G106gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(KEYINPUT69), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT67), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G99gat), .A2(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT66), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n443_), .A2(new_n444_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n431_), .B1(new_n441_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n433_), .A2(new_n434_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n447_), .A2(new_n445_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT7), .B1(new_n442_), .B2(KEYINPUT67), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT8), .B1(new_n427_), .B2(new_n430_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n449_), .A2(KEYINPUT8), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(KEYINPUT10), .B(G99gat), .Z(new_n456_));
  INV_X1    g255(.A(KEYINPUT65), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT10), .B(G99gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT65), .ZN(new_n460_));
  AOI21_X1  g259(.A(G106gat), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT9), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n429_), .A2(new_n424_), .A3(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n450_), .B1(KEYINPUT9), .B2(new_n426_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n461_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n423_), .B1(new_n455_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n463_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n464_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n459_), .B(new_n457_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n467_), .B(new_n468_), .C1(new_n469_), .C2(G106gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n423_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT8), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n435_), .B(new_n440_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n472_), .B1(new_n473_), .B2(new_n431_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n453_), .A2(new_n454_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n470_), .B(new_n471_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n466_), .A2(KEYINPUT12), .A3(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n470_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT12), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(new_n423_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n415_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n414_), .B1(new_n466_), .B2(new_n476_), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G120gat), .B(G148gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT5), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(new_n266_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(G204gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  OR3_X1    g287(.A1(new_n481_), .A2(new_n482_), .A3(new_n487_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(KEYINPUT70), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT70), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n483_), .A2(new_n491_), .A3(new_n487_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT13), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n490_), .A2(KEYINPUT13), .A3(new_n492_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G50gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G29gat), .B(G36gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT72), .ZN(new_n501_));
  INV_X1    g300(.A(G43gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT72), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G29gat), .A2(G36gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n501_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n502_), .B1(new_n501_), .B2(new_n507_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n499_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n507_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n505_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n512_));
  OAI21_X1  g311(.A(G43gat), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n501_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(G50gat), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n510_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G15gat), .B(G22gat), .ZN(new_n517_));
  INV_X1    g316(.A(G8gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G1gat), .B(G8gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n516_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT77), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n510_), .A2(new_n515_), .A3(new_n522_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n510_), .A2(new_n515_), .A3(KEYINPUT77), .A4(new_n522_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT15), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n508_), .A2(new_n509_), .A3(new_n499_), .ZN(new_n533_));
  AOI21_X1  g332(.A(G50gat), .B1(new_n513_), .B2(new_n514_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n510_), .A2(new_n515_), .A3(KEYINPUT15), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n522_), .A3(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(new_n529_), .A3(new_n524_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n531_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G113gat), .B(G141gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(G169gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n541_), .B(G197gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n539_), .B(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n498_), .A2(new_n544_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n412_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n535_), .A2(new_n536_), .A3(new_n478_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT73), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT71), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT34), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n548_), .A2(KEYINPUT35), .A3(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n516_), .B(new_n470_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n547_), .A2(new_n553_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n556_), .A2(KEYINPUT35), .A3(new_n551_), .A4(new_n548_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n551_), .A2(KEYINPUT35), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n555_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT75), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT74), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(G134gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n225_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT36), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n555_), .A2(new_n557_), .A3(KEYINPUT75), .A4(new_n558_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n561_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n559_), .A2(new_n569_), .A3(new_n565_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G127gat), .B(G155gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT16), .ZN(new_n573_));
  INV_X1    g372(.A(G183gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(G211gat), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n576_), .A2(new_n577_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n522_), .B(new_n423_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT76), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n580_), .B(new_n582_), .ZN(new_n583_));
  OR3_X1    g382(.A1(new_n578_), .A2(new_n579_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n579_), .A2(new_n583_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n571_), .A2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n546_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n202_), .B1(new_n588_), .B2(new_n388_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT102), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n555_), .A2(new_n557_), .A3(new_n566_), .A4(new_n558_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n570_), .A2(KEYINPUT37), .A3(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n571_), .B2(KEYINPUT37), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n586_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n546_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(new_n202_), .A3(new_n388_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT38), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n590_), .A2(new_n597_), .ZN(G1324gat));
  XNOR2_X1  g397(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT40), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n588_), .A2(new_n341_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(G8gat), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT39), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT39), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(new_n604_), .A3(G8gat), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n595_), .A2(new_n518_), .A3(new_n341_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n600_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n604_), .B1(new_n601_), .B2(G8gat), .ZN(new_n609_));
  AOI211_X1 g408(.A(KEYINPUT39), .B(new_n518_), .C1(new_n588_), .C2(new_n341_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n607_), .B(new_n600_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n608_), .A2(new_n612_), .ZN(G1325gat));
  INV_X1    g412(.A(G15gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n588_), .B2(new_n411_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT41), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n595_), .A2(new_n614_), .A3(new_n411_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1326gat));
  INV_X1    g417(.A(G22gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n262_), .B(KEYINPUT105), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n619_), .B1(new_n588_), .B2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT42), .Z(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n619_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT106), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n595_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(G1327gat));
  INV_X1    g426(.A(G29gat), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n568_), .A2(new_n570_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n586_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n546_), .A2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n632_), .B2(new_n389_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n545_), .A2(new_n586_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n412_), .A2(new_n636_), .A3(new_n593_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n636_), .B1(new_n412_), .B2(new_n593_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(G29gat), .A3(new_n388_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n412_), .A2(new_n593_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT43), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n637_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(KEYINPUT44), .A3(new_n635_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n633_), .B1(new_n643_), .B2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT107), .ZN(G1328gat));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n341_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n634_), .B1(new_n645_), .B2(new_n637_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(KEYINPUT44), .ZN(new_n653_));
  OAI21_X1  g452(.A(G36gat), .B1(new_n651_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT108), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT46), .ZN(new_n656_));
  INV_X1    g455(.A(new_n632_), .ZN(new_n657_));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n657_), .A2(KEYINPUT45), .A3(new_n658_), .A4(new_n341_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT45), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n546_), .A2(new_n658_), .A3(new_n631_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n341_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n660_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n659_), .A2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n654_), .A2(new_n655_), .A3(new_n656_), .A4(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n655_), .A2(new_n656_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n662_), .B1(new_n652_), .B2(KEYINPUT44), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n658_), .B1(new_n668_), .B2(new_n642_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n659_), .A2(new_n663_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n666_), .B(new_n667_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n665_), .A2(new_n671_), .ZN(G1329gat));
  OAI21_X1  g471(.A(new_n502_), .B1(new_n632_), .B2(new_n361_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT109), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n642_), .A2(new_n647_), .A3(G43gat), .A4(new_n411_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT47), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT47), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n674_), .A2(new_n678_), .A3(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1330gat));
  AOI21_X1  g479(.A(G50gat), .B1(new_n657_), .B2(new_n621_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n648_), .A2(new_n653_), .A3(new_n499_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(new_n263_), .ZN(G1331gat));
  NOR2_X1   g482(.A1(new_n497_), .A2(new_n543_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n412_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n594_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G57gat), .B1(new_n687_), .B2(new_n388_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n685_), .A2(new_n587_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n388_), .A2(G57gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(G1332gat));
  INV_X1    g490(.A(G64gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n689_), .B2(new_n341_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT48), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n687_), .A2(new_n692_), .A3(new_n341_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1333gat));
  INV_X1    g495(.A(G71gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n689_), .B2(new_n411_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT49), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n687_), .A2(new_n697_), .A3(new_n411_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1334gat));
  NAND2_X1  g500(.A1(new_n689_), .A2(new_n621_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G78gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n620_), .A2(G78gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n686_), .B2(new_n706_), .ZN(G1335gat));
  NAND2_X1  g506(.A1(new_n685_), .A2(new_n631_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G85gat), .B1(new_n709_), .B2(new_n388_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n586_), .B(new_n684_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n388_), .A2(G85gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n710_), .B1(new_n712_), .B2(new_n713_), .ZN(G1336gat));
  AOI21_X1  g513(.A(G92gat), .B1(new_n709_), .B2(new_n341_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n662_), .A2(new_n322_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n712_), .B2(new_n716_), .ZN(G1337gat));
  OR3_X1    g516(.A1(new_n708_), .A2(new_n469_), .A3(new_n361_), .ZN(new_n718_));
  OAI211_X1 g517(.A(KEYINPUT111), .B(G99gat), .C1(new_n711_), .C2(new_n361_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n646_), .A2(new_n411_), .A3(new_n586_), .A4(new_n684_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT111), .B1(new_n721_), .B2(G99gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT51), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT51), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n725_), .B(new_n718_), .C1(new_n720_), .C2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1338gat));
  OR3_X1    g526(.A1(new_n708_), .A2(G106gat), .A3(new_n262_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n729_), .B(G106gat), .C1(new_n711_), .C2(new_n262_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n646_), .A2(new_n263_), .A3(new_n586_), .A4(new_n684_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n729_), .B1(new_n732_), .B2(G106gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n728_), .B1(new_n731_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT53), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT53), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n736_), .B(new_n728_), .C1(new_n731_), .C2(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1339gat));
  INV_X1    g537(.A(KEYINPUT117), .ZN(new_n739_));
  INV_X1    g538(.A(new_n489_), .ZN(new_n740_));
  OAI21_X1  g539(.A(KEYINPUT55), .B1(new_n481_), .B2(KEYINPUT115), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT115), .B1(new_n481_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n477_), .A2(new_n480_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT114), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n477_), .A2(new_n747_), .A3(new_n480_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n746_), .A2(new_n415_), .A3(new_n748_), .ZN(new_n749_));
  OAI211_X1 g548(.A(KEYINPUT115), .B(KEYINPUT55), .C1(new_n481_), .C2(new_n742_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n744_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n487_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT56), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n487_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n740_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n539_), .A2(new_n542_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n542_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT116), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n537_), .A2(new_n530_), .A3(new_n524_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT58), .B1(new_n756_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n592_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT37), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n629_), .B2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n739_), .B1(new_n763_), .B2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n756_), .A2(KEYINPUT58), .A3(new_n762_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n755_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT56), .B1(new_n751_), .B2(new_n487_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n489_), .B(new_n762_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT58), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(KEYINPUT117), .A3(new_n593_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n767_), .A2(new_n768_), .A3(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT112), .B1(new_n544_), .B2(new_n740_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n543_), .A2(new_n489_), .A3(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n776_), .B(new_n778_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n762_), .A2(new_n492_), .A3(new_n490_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT57), .B1(new_n781_), .B2(new_n629_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n783_));
  AOI211_X1 g582(.A(new_n783_), .B(new_n571_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n775_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n586_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n498_), .A2(new_n543_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n594_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n594_), .B2(new_n788_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n787_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(new_n388_), .A3(new_n362_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n795_), .A2(KEYINPUT59), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n544_), .A2(new_n343_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n798_), .A2(new_n799_), .A3(new_n800_), .A4(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(G113gat), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n801_), .A2(KEYINPUT118), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n796_), .B(new_n543_), .C1(new_n797_), .C2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1340gat));
  NAND2_X1  g605(.A1(new_n798_), .A2(new_n800_), .ZN(new_n807_));
  OAI21_X1  g606(.A(G120gat), .B1(new_n807_), .B2(new_n497_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n347_), .B1(new_n497_), .B2(KEYINPUT60), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n347_), .A2(KEYINPUT60), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(KEYINPUT119), .B2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n796_), .B(new_n811_), .C1(KEYINPUT119), .C2(new_n809_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n808_), .A2(new_n812_), .ZN(G1341gat));
  AOI21_X1  g612(.A(G127gat), .B1(new_n796_), .B2(new_n630_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n807_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n630_), .A2(G127gat), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n814_), .B1(new_n815_), .B2(new_n816_), .ZN(G1342gat));
  AOI21_X1  g616(.A(G134gat), .B1(new_n796_), .B2(new_n571_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n593_), .A2(G134gat), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n815_), .B2(new_n819_), .ZN(G1343gat));
  NOR2_X1   g619(.A1(new_n411_), .A2(new_n262_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n794_), .A2(new_n388_), .A3(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n822_), .A2(new_n341_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n543_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n498_), .ZN(new_n826_));
  XOR2_X1   g625(.A(KEYINPUT120), .B(G148gat), .Z(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1345gat));
  NAND2_X1  g627(.A1(new_n823_), .A2(new_n630_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT121), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n829_), .B(new_n831_), .ZN(G1346gat));
  OR2_X1    g631(.A1(new_n822_), .A2(new_n341_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n833_), .A2(new_n225_), .A3(new_n766_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT122), .B(new_n225_), .C1(new_n833_), .C2(new_n629_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n822_), .A2(new_n341_), .A3(new_n629_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(G162gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n834_), .B1(new_n835_), .B2(new_n838_), .ZN(G1347gat));
  INV_X1    g638(.A(KEYINPUT62), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n662_), .A2(new_n388_), .A3(new_n361_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n794_), .A2(new_n620_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n543_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n840_), .B1(new_n844_), .B2(G169gat), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n840_), .B(G169gat), .C1(new_n842_), .C2(new_n544_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n543_), .A2(new_n265_), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(KEYINPUT123), .Z(new_n849_));
  OAI22_X1  g648(.A1(new_n845_), .A2(new_n847_), .B1(new_n842_), .B2(new_n849_), .ZN(G1348gat));
  NAND3_X1  g649(.A1(new_n794_), .A2(new_n262_), .A3(new_n841_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n851_), .A2(new_n266_), .A3(new_n497_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n843_), .A2(new_n498_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n266_), .B2(new_n853_), .ZN(G1349gat));
  NOR3_X1   g653(.A1(new_n842_), .A2(new_n281_), .A3(new_n586_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n851_), .A2(new_n586_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT124), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n857_), .B2(new_n574_), .ZN(G1350gat));
  NAND3_X1  g657(.A1(new_n843_), .A2(new_n297_), .A3(new_n571_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G190gat), .B1(new_n842_), .B2(new_n766_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1351gat));
  AOI21_X1  g660(.A(new_n792_), .B1(new_n786_), .B2(new_n586_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n662_), .A2(new_n388_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n821_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT125), .B1(new_n862_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT125), .ZN(new_n866_));
  INV_X1    g665(.A(new_n864_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n630_), .B1(new_n775_), .B2(new_n785_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n866_), .B(new_n867_), .C1(new_n868_), .C2(new_n792_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n865_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n543_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n498_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n874_));
  XOR2_X1   g673(.A(new_n873_), .B(new_n874_), .Z(G1353gat));
  NOR2_X1   g674(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n870_), .B2(new_n630_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT63), .B(G211gat), .Z(new_n878_));
  AOI211_X1 g677(.A(new_n586_), .B(new_n878_), .C1(new_n865_), .C2(new_n869_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT127), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n878_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n870_), .A2(new_n630_), .A3(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT127), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n586_), .B1(new_n865_), .B2(new_n869_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n882_), .B(new_n883_), .C1(new_n884_), .C2(new_n876_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n880_), .A2(new_n885_), .ZN(G1354gat));
  AOI21_X1  g685(.A(G218gat), .B1(new_n870_), .B2(new_n571_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n766_), .B1(new_n865_), .B2(new_n869_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(G218gat), .ZN(G1355gat));
endmodule


