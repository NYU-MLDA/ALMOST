//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n955_, new_n956_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_;
  XOR2_X1   g000(.A(G71gat), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT30), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206_));
  INV_X1    g005(.A(G15gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n205_), .B(new_n208_), .Z(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  INV_X1    g010(.A(G183gat), .ZN(new_n212_));
  INV_X1    g011(.A(G190gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n211_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n213_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT22), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G169gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT83), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT82), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(new_n218_), .B2(G169gat), .ZN(new_n223_));
  INV_X1    g022(.A(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(KEYINPUT82), .A3(KEYINPUT22), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n210_), .B(new_n217_), .C1(new_n221_), .C2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT26), .B(G190gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT25), .B1(new_n212_), .B2(KEYINPUT81), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n212_), .A2(KEYINPUT25), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n229_), .B(new_n230_), .C1(new_n231_), .C2(KEYINPUT81), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n225_), .A2(new_n224_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(KEYINPUT24), .A3(new_n210_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(KEYINPUT24), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n214_), .A2(new_n215_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n232_), .A2(new_n234_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n228_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n209_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n205_), .B(new_n208_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n228_), .A2(new_n237_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT86), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT31), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G113gat), .B(G120gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT84), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G134gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G127gat), .ZN(new_n251_));
  INV_X1    g050(.A(G127gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G134gat), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n251_), .A2(new_n253_), .A3(new_n248_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n246_), .B1(new_n249_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n253_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT84), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n247_), .A2(new_n248_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n246_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT85), .B1(new_n255_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT85), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n249_), .A2(new_n254_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n262_), .B1(new_n263_), .B2(new_n259_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT31), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n239_), .A2(new_n242_), .A3(new_n243_), .A4(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n245_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n265_), .B1(new_n245_), .B2(new_n267_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n255_), .A2(new_n260_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n262_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT3), .ZN(new_n273_));
  INV_X1    g072(.A(G141gat), .ZN(new_n274_));
  INV_X1    g073(.A(G148gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n276_), .A2(new_n279_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G141gat), .B(G148gat), .Z(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(KEYINPUT1), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n283_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n284_), .A2(KEYINPUT1), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n287_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n263_), .A2(new_n259_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT85), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n272_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT97), .ZN(new_n296_));
  INV_X1    g095(.A(new_n292_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n297_), .B2(new_n271_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT98), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n272_), .A2(new_n294_), .A3(new_n296_), .A4(new_n292_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n299_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n295_), .A2(KEYINPUT4), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n261_), .A2(new_n264_), .A3(new_n297_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n297_), .A2(new_n271_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT97), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n303_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n305_), .B1(new_n309_), .B2(KEYINPUT4), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n304_), .B1(new_n310_), .B2(new_n302_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G1gat), .B(G29gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(G85gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT0), .B(G57gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n313_), .B(new_n314_), .Z(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT4), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n301_), .B1(new_n318_), .B2(new_n305_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n315_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n304_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n270_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT20), .ZN(new_n325_));
  OR2_X1    g124(.A1(G197gat), .A2(G204gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G197gat), .A2(G204gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G211gat), .B(G218gat), .Z(new_n329_));
  NAND4_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(KEYINPUT89), .A4(KEYINPUT21), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT89), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n326_), .A2(KEYINPUT21), .A3(new_n327_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G211gat), .B(G218gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n332_), .A2(new_n333_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n326_), .A2(new_n327_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT21), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n335_), .A2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n325_), .B1(new_n238_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT93), .ZN(new_n343_));
  XOR2_X1   g142(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n344_));
  NAND2_X1  g143(.A1(G226gat), .A2(G233gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n217_), .A2(KEYINPUT92), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n217_), .A2(KEYINPUT92), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT22), .B(G169gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n224_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n347_), .A2(new_n210_), .A3(new_n348_), .A4(new_n350_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n334_), .A2(new_n330_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT25), .B(G183gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n229_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n236_), .A2(new_n354_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n352_), .A3(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n342_), .A2(new_n343_), .A3(new_n346_), .A4(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n342_), .A2(new_n346_), .A3(new_n356_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT93), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n325_), .B1(new_n241_), .B2(new_n352_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n351_), .A2(new_n355_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n341_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n346_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n357_), .B1(new_n359_), .B2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G8gat), .B(G36gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n364_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT95), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n369_), .B(new_n357_), .C1(new_n359_), .C2(new_n363_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT27), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n359_), .A2(new_n363_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n376_), .A2(KEYINPUT95), .A3(new_n369_), .A4(new_n357_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n360_), .A2(new_n362_), .A3(new_n346_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n342_), .A2(new_n356_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n379_), .B1(new_n380_), .B2(new_n346_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n375_), .B1(new_n381_), .B2(new_n369_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n371_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n378_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G22gat), .B(G50gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n352_), .B1(KEYINPUT29), .B2(new_n292_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n390_), .A2(KEYINPUT90), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n388_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n390_), .A2(KEYINPUT90), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n292_), .A2(KEYINPUT29), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n341_), .A2(new_n394_), .B1(KEYINPUT90), .B2(new_n390_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n387_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n392_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT88), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n393_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n386_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n399_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n386_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n401_), .A2(KEYINPUT88), .A3(new_n402_), .A4(new_n397_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n292_), .A2(KEYINPUT29), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n404_), .B(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT100), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n385_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n404_), .B(new_n407_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT100), .B1(new_n412_), .B2(new_n384_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n324_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n315_), .B1(new_n310_), .B2(new_n302_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n302_), .B1(new_n309_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n416_), .B2(new_n309_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  AOI211_X1 g218(.A(KEYINPUT33), .B(new_n320_), .C1(new_n319_), .C2(new_n304_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n311_), .B2(new_n315_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n419_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n374_), .A2(KEYINPUT96), .A3(new_n377_), .ZN(new_n424_));
  AOI21_X1  g223(.A(KEYINPUT96), .B1(new_n374_), .B2(new_n377_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT32), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n364_), .B1(new_n427_), .B2(new_n369_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n381_), .A2(KEYINPUT32), .A3(new_n370_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n322_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n409_), .B1(new_n426_), .B2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n409_), .A2(new_n322_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n385_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n270_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n414_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G229gat), .A2(G233gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G29gat), .B(G36gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G43gat), .B(G50gat), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n440_), .A2(new_n441_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G1gat), .B(G8gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(G22gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(KEYINPUT72), .A2(G15gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(KEYINPUT72), .A2(G15gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n447_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT72), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n207_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(G22gat), .A3(new_n448_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT14), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(G1gat), .B2(G8gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n446_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n459_));
  AOI211_X1 g258(.A(new_n457_), .B(new_n445_), .C1(new_n451_), .C2(new_n454_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n444_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n449_), .A2(new_n450_), .A3(new_n447_), .ZN(new_n462_));
  AOI21_X1  g261(.A(G22gat), .B1(new_n453_), .B2(new_n448_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n458_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n445_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n455_), .A2(new_n446_), .A3(new_n458_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n440_), .B(new_n441_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n461_), .A2(new_n468_), .A3(KEYINPUT77), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT77), .B1(new_n461_), .B2(new_n468_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n439_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n444_), .A2(KEYINPUT15), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT15), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n467_), .A2(new_n473_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n472_), .B(new_n474_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n468_), .A3(new_n438_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G113gat), .B(G141gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT78), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G169gat), .B(G197gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n471_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT79), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT79), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n471_), .A2(new_n483_), .A3(new_n476_), .A4(new_n480_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n471_), .A2(new_n476_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n480_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT80), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT80), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n485_), .A2(new_n491_), .A3(new_n488_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n437_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G230gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT64), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT6), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT6), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(G99gat), .A3(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n503_));
  INV_X1    g302(.A(G106gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G85gat), .ZN(new_n507_));
  INV_X1    g306(.A(G92gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G85gat), .A2(G92gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(KEYINPUT9), .A3(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n510_), .A2(KEYINPUT9), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n502_), .A2(new_n506_), .A3(new_n511_), .A4(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n509_), .A2(new_n510_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n499_), .A2(new_n501_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n518_));
  INV_X1    g317(.A(G99gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(new_n504_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n516_), .B1(new_n517_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT8), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n502_), .A2(new_n521_), .A3(new_n520_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT8), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n516_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n514_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G57gat), .B(G64gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G71gat), .B(G78gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(KEYINPUT11), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n532_));
  INV_X1    g331(.A(new_n530_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n531_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n528_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT12), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n528_), .A2(new_n536_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n521_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI211_X1 g342(.A(KEYINPUT8), .B(new_n515_), .C1(new_n543_), .C2(new_n502_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n526_), .B1(new_n525_), .B2(new_n516_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n544_), .A2(new_n545_), .A3(KEYINPUT65), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT65), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n547_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n513_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT12), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n536_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT66), .B1(new_n549_), .B2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT65), .B1(new_n544_), .B2(new_n545_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n524_), .A2(new_n547_), .A3(new_n527_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n514_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT66), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n551_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n497_), .B(new_n540_), .C1(new_n553_), .C2(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n539_), .A2(new_n537_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n559_), .B1(new_n497_), .B2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G120gat), .B(G148gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT5), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G176gat), .B(G204gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n565_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n569_), .A2(KEYINPUT13), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(KEYINPUT13), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT37), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT35), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT67), .B(KEYINPUT34), .Z(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n528_), .A2(new_n467_), .B1(new_n574_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n472_), .A2(new_n474_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n578_), .B1(new_n556_), .B2(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n577_), .A2(new_n574_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n578_), .B(new_n581_), .C1(new_n556_), .C2(new_n579_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT36), .Z(new_n589_));
  NAND2_X1  g388(.A1(new_n585_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT69), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n583_), .A2(new_n592_), .A3(new_n584_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT68), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n573_), .B1(new_n591_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT71), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n585_), .A2(KEYINPUT70), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT70), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n597_), .B1(new_n601_), .B2(new_n589_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n597_), .B(new_n589_), .C1(new_n598_), .C2(new_n600_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n595_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n596_), .B1(new_n605_), .B2(new_n573_), .ZN(new_n606_));
  XOR2_X1   g405(.A(G183gat), .B(G211gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT74), .ZN(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G127gat), .B(G155gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT76), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT17), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n465_), .A2(new_n466_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(new_n536_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n620_));
  OR3_X1    g419(.A1(new_n618_), .A2(new_n612_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n606_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n495_), .A2(new_n572_), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT101), .ZN(new_n625_));
  INV_X1    g424(.A(G1gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n626_), .A3(new_n322_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n437_), .A2(new_n605_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n572_), .A2(new_n493_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n631_), .A2(new_n622_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G1gat), .B1(new_n633_), .B2(new_n323_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n627_), .A2(new_n628_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n629_), .A2(new_n634_), .A3(new_n635_), .ZN(G1324gat));
  INV_X1    g435(.A(G8gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n625_), .A2(new_n637_), .A3(new_n384_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G8gat), .B1(new_n633_), .B2(new_n385_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT102), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n642_), .B(G8gat), .C1(new_n633_), .C2(new_n385_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n640_), .A2(new_n641_), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n641_), .B1(new_n640_), .B2(new_n643_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n638_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n638_), .B(new_n647_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1325gat));
  OAI21_X1  g450(.A(G15gat), .B1(new_n633_), .B2(new_n436_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT41), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n625_), .A2(new_n207_), .A3(new_n270_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1326gat));
  XNOR2_X1  g454(.A(new_n409_), .B(KEYINPUT104), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n625_), .A2(new_n447_), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G22gat), .B1(new_n633_), .B2(new_n656_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT42), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(G1327gat));
  NAND2_X1  g460(.A1(new_n605_), .A2(new_n573_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n596_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT43), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n667_), .B1(new_n437_), .B2(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n374_), .A2(new_n377_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT96), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n316_), .A2(KEYINPUT33), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n311_), .A2(new_n421_), .A3(new_n315_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n374_), .A2(KEYINPUT96), .A3(new_n377_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n671_), .A2(new_n674_), .A3(new_n675_), .A4(new_n419_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n412_), .B1(new_n676_), .B2(new_n430_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n409_), .A2(new_n384_), .A3(new_n322_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n436_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n413_), .A2(new_n411_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n324_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n606_), .A3(new_n666_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n668_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n572_), .A2(new_n493_), .A3(new_n622_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT44), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689_));
  AOI211_X1 g488(.A(new_n689_), .B(new_n686_), .C1(new_n668_), .C2(new_n684_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n322_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G29gat), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n570_), .A2(new_n571_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n605_), .A2(new_n622_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n495_), .A2(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n323_), .A2(G29gat), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT106), .Z(new_n699_));
  OAI21_X1  g498(.A(new_n693_), .B1(new_n697_), .B2(new_n699_), .ZN(G1328gat));
  NOR3_X1   g499(.A1(new_n697_), .A2(G36gat), .A3(new_n385_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n691_), .B2(new_n384_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n683_), .A2(new_n606_), .A3(new_n666_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n666_), .B1(new_n683_), .B2(new_n606_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n687_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n689_), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT44), .B(new_n687_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n709_), .A2(new_n704_), .A3(new_n384_), .A4(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G36gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n703_), .B1(new_n705_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(KEYINPUT46), .B(new_n703_), .C1(new_n705_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  NOR3_X1   g516(.A1(new_n688_), .A2(new_n690_), .A3(new_n436_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n270_), .A2(new_n203_), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n718_), .A2(new_n203_), .B1(new_n697_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1330gat));
  OR3_X1    g521(.A1(new_n697_), .A2(G50gat), .A3(new_n656_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n709_), .A2(KEYINPUT109), .A3(new_n412_), .A4(new_n710_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(G50gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n709_), .A2(new_n412_), .A3(new_n710_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT110), .B1(new_n725_), .B2(new_n728_), .ZN(new_n729_));
  AND4_X1   g528(.A1(KEYINPUT110), .A2(new_n728_), .A3(G50gat), .A4(new_n724_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n723_), .B1(new_n729_), .B2(new_n730_), .ZN(G1331gat));
  NAND2_X1  g530(.A1(new_n694_), .A2(new_n494_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n732_), .A2(new_n622_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n630_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G57gat), .B1(new_n734_), .B2(new_n323_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n437_), .A2(new_n493_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n694_), .A3(new_n623_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n323_), .A2(G57gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n737_), .B2(new_n738_), .ZN(G1332gat));
  OAI21_X1  g538(.A(G64gat), .B1(new_n734_), .B2(new_n385_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT48), .ZN(new_n741_));
  OR3_X1    g540(.A1(new_n737_), .A2(G64gat), .A3(new_n385_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(G1333gat));
  OAI21_X1  g544(.A(G71gat), .B1(new_n734_), .B2(new_n436_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT49), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n436_), .A2(G71gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n737_), .B2(new_n748_), .ZN(G1334gat));
  OAI21_X1  g548(.A(G78gat), .B1(new_n734_), .B2(new_n656_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT50), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n656_), .A2(G78gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n737_), .B2(new_n752_), .ZN(G1335gat));
  NOR4_X1   g552(.A1(new_n437_), .A2(new_n493_), .A3(new_n572_), .A4(new_n695_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n507_), .A3(new_n322_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n756_));
  INV_X1    g555(.A(new_n622_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n732_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n685_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n685_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n323_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n755_), .B1(new_n762_), .B2(new_n507_), .ZN(G1336gat));
  NAND3_X1  g562(.A1(new_n754_), .A2(new_n508_), .A3(new_n384_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n385_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n508_), .ZN(G1337gat));
  INV_X1    g565(.A(new_n761_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n270_), .B1(new_n767_), .B2(new_n759_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(G99gat), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n270_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT113), .B1(new_n754_), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n769_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1338gat));
  NAND3_X1  g574(.A1(new_n754_), .A2(new_n504_), .A3(new_n412_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n685_), .A2(new_n412_), .A3(new_n758_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(G106gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n777_), .B2(G106gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g581(.A1(new_n623_), .A2(new_n572_), .A3(new_n494_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT77), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n459_), .A2(new_n460_), .A3(new_n444_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n467_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n787_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n461_), .A2(new_n468_), .A3(KEYINPUT77), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n439_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n475_), .A2(new_n468_), .A3(new_n439_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n487_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT117), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n438_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n788_), .A2(new_n438_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n480_), .B1(new_n797_), .B2(new_n475_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  AOI221_X4 g599(.A(KEYINPUT118), .B1(new_n795_), .B2(new_n800_), .C1(new_n482_), .C2(new_n484_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n795_), .A2(new_n800_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n485_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n566_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n549_), .A2(KEYINPUT66), .A3(new_n552_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n557_), .B1(new_n556_), .B2(new_n551_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n806_), .A2(new_n807_), .B1(new_n539_), .B2(new_n538_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT115), .B1(new_n808_), .B2(new_n497_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n540_), .B1(new_n553_), .B2(new_n558_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  INV_X1    g610(.A(new_n497_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n809_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n559_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n808_), .A2(KEYINPUT55), .A3(new_n497_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n565_), .B1(new_n814_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n809_), .A2(new_n816_), .A3(new_n813_), .A4(new_n817_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(KEYINPUT56), .A3(new_n565_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n805_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n786_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n561_), .A2(new_n565_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n804_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n485_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n827_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n823_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT56), .B1(new_n822_), .B2(new_n565_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n830_), .B(new_n825_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n606_), .B1(new_n826_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n824_), .A2(KEYINPUT58), .ZN(new_n838_));
  OAI211_X1 g637(.A(KEYINPUT121), .B(new_n606_), .C1(new_n826_), .C2(new_n834_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n494_), .A2(new_n827_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n832_), .A2(KEYINPUT116), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n823_), .B1(new_n832_), .B2(KEYINPUT116), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n841_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n569_), .B1(new_n829_), .B2(new_n828_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n605_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT57), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n848_), .B2(KEYINPUT57), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n832_), .A2(KEYINPUT116), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n842_), .A3(new_n823_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n846_), .B1(new_n854_), .B2(new_n841_), .ZN(new_n855_));
  OAI211_X1 g654(.A(KEYINPUT119), .B(new_n852_), .C1(new_n855_), .C2(new_n605_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n840_), .A2(new_n849_), .A3(new_n851_), .A4(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n785_), .B1(new_n857_), .B2(new_n622_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n680_), .A2(new_n322_), .A3(new_n270_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT59), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n852_), .B1(new_n855_), .B2(new_n605_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n839_), .A2(new_n838_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n830_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT120), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(new_n786_), .A3(new_n833_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT121), .B1(new_n865_), .B2(new_n606_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n849_), .B(new_n861_), .C1(new_n862_), .C2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n622_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n785_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n859_), .A2(KEYINPUT59), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n860_), .A2(new_n493_), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G113gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n849_), .B1(new_n862_), .B2(new_n866_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n851_), .A2(new_n856_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n622_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n869_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n859_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n494_), .A2(G113gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n874_), .B1(new_n880_), .B2(new_n881_), .ZN(G1340gat));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n572_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n860_), .B2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n883_), .A2(KEYINPUT60), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n887_));
  AOI21_X1  g686(.A(G120gat), .B1(new_n694_), .B2(new_n887_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n880_), .A2(new_n886_), .A3(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT122), .B1(new_n885_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n785_), .B1(new_n867_), .B2(new_n622_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n871_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n694_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G120gat), .B1(new_n892_), .B2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897_));
  OR4_X1    g696(.A1(new_n858_), .A2(new_n859_), .A3(new_n886_), .A4(new_n888_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n890_), .A2(new_n899_), .ZN(G1341gat));
  INV_X1    g699(.A(new_n880_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n901_), .A2(new_n252_), .A3(new_n757_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n860_), .A2(new_n757_), .A3(new_n872_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n902_), .B1(new_n904_), .B2(new_n252_), .ZN(G1342gat));
  NAND3_X1  g704(.A1(new_n901_), .A2(new_n250_), .A3(new_n605_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n860_), .A2(new_n606_), .A3(new_n872_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n908_), .B2(new_n250_), .ZN(G1343gat));
  NOR3_X1   g708(.A1(new_n270_), .A2(new_n409_), .A3(new_n323_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n878_), .A2(new_n385_), .A3(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n494_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n274_), .ZN(G1344gat));
  NOR2_X1   g712(.A1(new_n911_), .A2(new_n572_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n275_), .ZN(G1345gat));
  NOR2_X1   g714(.A1(new_n911_), .A2(new_n622_), .ZN(new_n916_));
  XOR2_X1   g715(.A(KEYINPUT61), .B(G155gat), .Z(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1346gat));
  OAI21_X1  g717(.A(G162gat), .B1(new_n911_), .B2(new_n664_), .ZN(new_n919_));
  OR3_X1    g718(.A1(new_n602_), .A2(new_n604_), .A3(G162gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n911_), .B2(new_n920_), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n324_), .A2(new_n385_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n656_), .ZN(new_n923_));
  OR3_X1    g722(.A1(new_n893_), .A2(KEYINPUT123), .A3(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT123), .B1(new_n893_), .B2(new_n923_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n926_), .A2(new_n349_), .A3(new_n493_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n893_), .A2(new_n923_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n493_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n928_), .B1(new_n930_), .B2(G169gat), .ZN(new_n931_));
  AOI211_X1 g730(.A(KEYINPUT62), .B(new_n225_), .C1(new_n929_), .C2(new_n493_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n927_), .B1(new_n931_), .B2(new_n932_), .ZN(G1348gat));
  NOR2_X1   g732(.A1(new_n858_), .A2(new_n412_), .ZN(new_n934_));
  AND4_X1   g733(.A1(G176gat), .A2(new_n934_), .A3(new_n694_), .A4(new_n922_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n926_), .A2(new_n694_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n936_), .B2(new_n224_), .ZN(G1349gat));
  NOR2_X1   g736(.A1(new_n622_), .A2(new_n353_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n934_), .A2(new_n757_), .A3(new_n922_), .ZN(new_n939_));
  AOI22_X1  g738(.A1(new_n926_), .A2(new_n938_), .B1(new_n939_), .B2(new_n212_), .ZN(G1350gat));
  INV_X1    g739(.A(new_n926_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n605_), .A2(new_n229_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(KEYINPUT124), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n664_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n944_));
  OAI22_X1  g743(.A1(new_n941_), .A2(new_n943_), .B1(new_n944_), .B2(new_n213_), .ZN(G1351gat));
  AND3_X1   g744(.A1(new_n433_), .A2(KEYINPUT125), .A3(new_n436_), .ZN(new_n946_));
  AOI21_X1  g745(.A(KEYINPUT125), .B1(new_n433_), .B2(new_n436_), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n946_), .A2(new_n947_), .A3(new_n385_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n878_), .A2(new_n493_), .A3(new_n948_), .ZN(new_n949_));
  INV_X1    g748(.A(G197gat), .ZN(new_n950_));
  OR3_X1    g749(.A1(new_n949_), .A2(KEYINPUT126), .A3(new_n950_), .ZN(new_n951_));
  OAI21_X1  g750(.A(KEYINPUT126), .B1(new_n949_), .B2(new_n950_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n949_), .A2(new_n950_), .ZN(new_n953_));
  AND3_X1   g752(.A1(new_n951_), .A2(new_n952_), .A3(new_n953_), .ZN(G1352gat));
  AND2_X1   g753(.A1(new_n878_), .A2(new_n948_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(new_n694_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g756(.A(new_n622_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n955_), .A2(new_n958_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n960_), .B(new_n961_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n959_), .A2(new_n962_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n960_), .A2(new_n961_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n955_), .A2(new_n958_), .A3(new_n964_), .ZN(new_n965_));
  AND2_X1   g764(.A1(new_n963_), .A2(new_n965_), .ZN(G1354gat));
  INV_X1    g765(.A(G218gat), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n955_), .A2(new_n967_), .A3(new_n605_), .ZN(new_n968_));
  AND2_X1   g767(.A1(new_n955_), .A2(new_n606_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n968_), .B1(new_n969_), .B2(new_n967_), .ZN(G1355gat));
endmodule


