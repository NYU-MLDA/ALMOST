//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G211gat), .A2(G218gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G211gat), .A2(G218gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  AND2_X1   g009(.A1(G211gat), .A2(G218gat), .ZN(new_n211_));
  NOR3_X1   g010(.A1(new_n211_), .A2(new_n206_), .A3(KEYINPUT83), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n205_), .B(new_n210_), .C1(new_n212_), .C2(new_n208_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n207_), .A2(new_n209_), .ZN(new_n214_));
  OAI211_X1 g013(.A(KEYINPUT21), .B(new_n204_), .C1(new_n214_), .C2(KEYINPUT83), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT84), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n213_), .A2(KEYINPUT84), .A3(new_n215_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT29), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT81), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT81), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(G155gat), .A3(G162gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT1), .ZN(new_n227_));
  OR2_X1    g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n223_), .A2(new_n225_), .A3(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G141gat), .A2(G148gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G141gat), .A2(G148gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT2), .B1(new_n233_), .B2(KEYINPUT82), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT82), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT2), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n232_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n237_), .A2(new_n239_), .A3(new_n242_), .A4(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(G155gat), .A2(G162gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n245_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n221_), .B1(new_n236_), .B2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n203_), .B1(new_n220_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT85), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n231_), .A2(new_n235_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n218_), .B(new_n219_), .C1(new_n252_), .C2(new_n221_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(KEYINPUT85), .A3(new_n203_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n216_), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n248_), .A2(new_n256_), .A3(new_n203_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n202_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n202_), .ZN(new_n260_));
  AOI211_X1 g059(.A(new_n257_), .B(new_n260_), .C1(new_n251_), .C2(new_n254_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT28), .B(G106gat), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n259_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n262_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n253_), .A2(KEYINPUT85), .A3(new_n203_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT85), .B1(new_n253_), .B2(new_n203_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n258_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n260_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n255_), .A2(new_n258_), .A3(new_n202_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n264_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n252_), .A2(new_n221_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT86), .B(G78gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n263_), .A2(new_n270_), .A3(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n262_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n268_), .A2(new_n269_), .A3(new_n264_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n273_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n236_), .A2(new_n247_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G127gat), .A2(G134gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G127gat), .A2(G134gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(G113gat), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(G127gat), .ZN(new_n284_));
  INV_X1    g083(.A(G134gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G113gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(new_n280_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n283_), .A2(new_n288_), .A3(G120gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(G120gat), .B1(new_n283_), .B2(new_n288_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n279_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n252_), .A2(new_n291_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT4), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT90), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT91), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n293_), .A2(KEYINPUT4), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT90), .A4(KEYINPUT4), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n297_), .A2(new_n300_), .A3(new_n301_), .A4(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n293_), .A2(new_n294_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n298_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT92), .B(KEYINPUT0), .Z(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G29gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G57gat), .B(G85gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n306_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT94), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n303_), .A2(new_n305_), .A3(new_n311_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT94), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n306_), .A2(new_n316_), .A3(new_n312_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT23), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G169gat), .ZN(new_n324_));
  INV_X1    g123(.A(G176gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n326_), .A2(KEYINPUT24), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(KEYINPUT24), .A3(new_n328_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n323_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n331_));
  AND2_X1   g130(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n332_));
  AND2_X1   g131(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n334_));
  OAI22_X1  g133(.A1(new_n331_), .A2(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n321_), .A2(new_n336_), .A3(new_n322_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n337_), .A2(new_n328_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT22), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(G169gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT22), .B(G169gat), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n325_), .B(new_n341_), .C1(new_n342_), .C2(new_n339_), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n330_), .A2(new_n335_), .B1(new_n338_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT88), .B1(new_n344_), .B2(new_n256_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT19), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n323_), .A2(new_n327_), .A3(new_n335_), .A4(new_n329_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n342_), .A2(new_n325_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n328_), .A2(KEYINPUT87), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n328_), .A2(KEYINPUT87), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n349_), .A2(new_n337_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n347_), .B1(new_n354_), .B2(new_n256_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n338_), .A2(new_n343_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n348_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT88), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(new_n358_), .A3(new_n216_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n345_), .A2(new_n355_), .A3(KEYINPUT20), .A4(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G8gat), .B(G36gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT18), .ZN(new_n362_));
  INV_X1    g161(.A(G64gat), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n363_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n364_), .A2(new_n365_), .A3(G92gat), .ZN(new_n366_));
  AOI21_X1  g165(.A(G92gat), .B1(new_n364_), .B2(new_n365_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n356_), .A2(new_n215_), .A3(new_n213_), .A4(new_n348_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n353_), .A2(new_n216_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n370_), .A3(KEYINPUT20), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n347_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n360_), .A2(new_n368_), .A3(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n345_), .A2(KEYINPUT20), .A3(new_n359_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n353_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n347_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n347_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n369_), .A2(new_n370_), .A3(KEYINPUT20), .A4(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT93), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n378_), .A2(new_n379_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n376_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n368_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n373_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT27), .ZN(new_n385_));
  XOR2_X1   g184(.A(KEYINPUT95), .B(KEYINPUT27), .Z(new_n386_));
  NAND2_X1  g185(.A1(new_n360_), .A2(new_n372_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n383_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n360_), .A2(new_n368_), .A3(new_n372_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n385_), .A2(new_n391_), .ZN(new_n392_));
  OAI22_X1  g191(.A1(new_n275_), .A2(new_n278_), .B1(new_n318_), .B2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n291_), .B(KEYINPUT31), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT80), .ZN(new_n395_));
  INV_X1    g194(.A(G99gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G15gat), .B(G71gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(new_n357_), .B(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n395_), .B(G99gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n399_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G227gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT30), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT79), .B(G43gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n406_), .B(new_n407_), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n404_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n368_), .A2(KEYINPUT32), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n382_), .A2(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n412_), .A2(new_n387_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n318_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n315_), .A2(KEYINPUT33), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n303_), .A2(new_n305_), .A3(new_n417_), .A4(new_n311_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n368_), .B1(new_n360_), .B2(new_n372_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT89), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n373_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT89), .B1(new_n388_), .B2(new_n389_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n297_), .A2(new_n298_), .A3(new_n301_), .A4(new_n302_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n304_), .A2(new_n300_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n312_), .A3(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n419_), .A2(new_n424_), .A3(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n274_), .B1(new_n263_), .B2(new_n270_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n276_), .A2(new_n273_), .A3(new_n277_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n393_), .B(new_n411_), .C1(new_n415_), .C2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT96), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n318_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n434_), .A2(new_n430_), .A3(new_n429_), .A4(new_n428_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n429_), .A2(new_n430_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n390_), .B1(new_n384_), .B2(KEYINPUT27), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n437_), .A2(new_n315_), .A3(new_n314_), .A4(new_n317_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n410_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT96), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n435_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n433_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n411_), .A2(new_n436_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n318_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n437_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G1gat), .B(G8gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT72), .ZN(new_n448_));
  OR2_X1    g247(.A1(G15gat), .A2(G22gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G15gat), .A2(G22gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G1gat), .A2(G8gat), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n449_), .A2(new_n450_), .B1(KEYINPUT14), .B2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n448_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G29gat), .B(G36gat), .ZN(new_n454_));
  INV_X1    g253(.A(G43gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G50gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n453_), .A2(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n459_), .B(KEYINPUT75), .Z(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(new_n453_), .B2(new_n458_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G229gat), .A2(G233gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n458_), .B(KEYINPUT15), .ZN(new_n465_));
  INV_X1    g264(.A(new_n453_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n460_), .A2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n464_), .B1(new_n463_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT77), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G113gat), .B(G141gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT76), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(new_n324_), .ZN(new_n473_));
  INV_X1    g272(.A(G197gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n469_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G57gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n363_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT11), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G57gat), .A2(G64gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  OR2_X1    g282(.A1(G71gat), .A2(G78gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G71gat), .A2(G78gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT66), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT66), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n483_), .A2(new_n488_), .A3(new_n484_), .A4(new_n485_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n480_), .A2(new_n482_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(new_n481_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n487_), .A2(new_n492_), .A3(new_n489_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(KEYINPUT12), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(G85gat), .A2(G92gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(G85gat), .A2(G92gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G99gat), .A2(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT6), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(G99gat), .A3(G106gat), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  INV_X1    g305(.A(G106gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n396_), .A3(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n500_), .B1(new_n505_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT8), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n502_), .A2(new_n504_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(new_n509_), .A3(new_n508_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n500_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n512_), .A2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n499_), .B1(new_n498_), .B2(KEYINPUT9), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT65), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n519_), .B1(new_n498_), .B2(KEYINPUT9), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G85gat), .A2(G92gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT9), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(KEYINPUT65), .A3(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n518_), .A2(new_n520_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n396_), .A2(KEYINPUT10), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT10), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(G99gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n528_), .A2(new_n507_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT68), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n523_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(G85gat), .B2(G92gat), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT65), .B1(new_n521_), .B2(new_n522_), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n532_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT10), .B(G99gat), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n513_), .B1(new_n537_), .B2(G106gat), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT68), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n517_), .A2(KEYINPUT69), .A3(new_n531_), .A4(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n524_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n530_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT69), .B1(new_n544_), .B2(new_n517_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n497_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n487_), .A2(new_n492_), .A3(new_n489_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n492_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n514_), .A2(new_n515_), .A3(new_n500_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n515_), .B1(new_n514_), .B2(new_n500_), .ZN(new_n551_));
  OAI22_X1  g350(.A1(new_n550_), .A2(new_n551_), .B1(new_n538_), .B2(new_n536_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT12), .B1(new_n549_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT64), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n556_), .B1(new_n549_), .B2(new_n552_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n546_), .A2(new_n554_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT67), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n560_), .B1(new_n549_), .B2(new_n552_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n494_), .A2(new_n495_), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n512_), .A2(new_n516_), .B1(new_n529_), .B2(new_n524_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(KEYINPUT67), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n549_), .A2(new_n552_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n559_), .B1(new_n567_), .B2(new_n556_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G120gat), .B(G148gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT5), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n325_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(G204gat), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n568_), .A2(new_n572_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT13), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n573_), .A2(KEYINPUT13), .A3(new_n574_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n478_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n446_), .A2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n465_), .B1(new_n545_), .B2(new_n541_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT71), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT70), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT34), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT35), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n458_), .A2(new_n563_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n582_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n586_), .A2(new_n587_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(G134gat), .ZN(new_n594_));
  INV_X1    g393(.A(G162gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT36), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n592_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n592_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n602_), .A2(KEYINPUT37), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(KEYINPUT37), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n562_), .B(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(new_n466_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G183gat), .B(G211gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT17), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n608_), .A2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT74), .Z(new_n617_));
  NOR2_X1   g416(.A1(new_n613_), .A2(new_n614_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n605_), .A2(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n581_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(G1gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n622_), .A3(new_n318_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT97), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT38), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n624_), .A2(new_n625_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT100), .ZN(new_n630_));
  INV_X1    g429(.A(new_n619_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n602_), .B(KEYINPUT99), .Z(new_n632_));
  NAND3_X1  g431(.A1(new_n581_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G1gat), .B1(new_n633_), .B2(new_n444_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(new_n630_), .A3(new_n634_), .ZN(G1324gat));
  OAI21_X1  g434(.A(G8gat), .B1(new_n633_), .B2(new_n437_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT39), .Z(new_n637_));
  INV_X1    g436(.A(new_n621_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(G8gat), .A3(new_n437_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g440(.A(G15gat), .B1(new_n633_), .B2(new_n411_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT101), .Z(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT41), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n411_), .A2(G15gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n638_), .B2(new_n645_), .ZN(G1326gat));
  INV_X1    g445(.A(new_n436_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G22gat), .B1(new_n633_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n647_), .A2(G22gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n650_), .B1(new_n638_), .B2(new_n651_), .ZN(G1327gat));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n603_), .A2(new_n604_), .ZN(new_n654_));
  AOI211_X1 g453(.A(KEYINPUT43), .B(new_n654_), .C1(new_n442_), .C2(new_n445_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n435_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n440_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n656_), .B(new_n445_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n605_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n656_), .B1(new_n442_), .B2(new_n445_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT43), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT104), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n664_), .B(KEYINPUT43), .C1(new_n660_), .C2(new_n661_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n655_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n619_), .A2(new_n580_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n653_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n653_), .B(KEYINPUT44), .C1(new_n666_), .C2(new_n667_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G29gat), .B1(new_n672_), .B2(new_n444_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n602_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n631_), .A2(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n581_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  OR3_X1    g476(.A1(new_n677_), .A2(G29gat), .A3(new_n444_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n673_), .A2(new_n678_), .ZN(G1328gat));
  INV_X1    g478(.A(G36gat), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n437_), .B(KEYINPUT106), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n676_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT45), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n437_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n684_), .B2(new_n680_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(KEYINPUT46), .B(new_n683_), .C1(new_n684_), .C2(new_n680_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1329gat));
  NOR3_X1   g488(.A1(new_n677_), .A2(G43gat), .A3(new_n411_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n411_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n692_), .B2(new_n455_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI211_X1 g494(.A(KEYINPUT47), .B(new_n691_), .C1(new_n692_), .C2(new_n455_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1330gat));
  OAI21_X1  g496(.A(G50gat), .B1(new_n672_), .B2(new_n647_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n676_), .A2(new_n457_), .A3(new_n436_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1331gat));
  INV_X1    g499(.A(new_n478_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n619_), .A2(new_n701_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n446_), .A2(new_n579_), .A3(new_n632_), .A4(new_n702_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n703_), .A2(new_n479_), .A3(new_n444_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n446_), .A2(new_n478_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT108), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n620_), .A2(new_n579_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT107), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n318_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n704_), .B1(new_n711_), .B2(new_n479_), .ZN(G1332gat));
  INV_X1    g511(.A(new_n681_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G64gat), .B1(new_n703_), .B2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT48), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n681_), .A2(new_n363_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n709_), .B2(new_n716_), .ZN(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n703_), .B2(new_n411_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n709_), .A2(G71gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(new_n411_), .ZN(G1334gat));
  OAI21_X1  g521(.A(G78gat), .B1(new_n703_), .B2(new_n647_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT50), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n647_), .A2(G78gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n709_), .B2(new_n725_), .ZN(G1335gat));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n666_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n619_), .A2(new_n478_), .A3(new_n579_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT112), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n666_), .A2(new_n727_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n728_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(G85gat), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n444_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n706_), .A2(new_n579_), .A3(new_n675_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n318_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n735_), .A2(new_n739_), .ZN(G1336gat));
  INV_X1    g539(.A(G92gat), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n733_), .A2(new_n741_), .A3(new_n713_), .ZN(new_n742_));
  AOI21_X1  g541(.A(G92gat), .B1(new_n738_), .B2(new_n392_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1337gat));
  OAI21_X1  g543(.A(G99gat), .B1(new_n733_), .B2(new_n411_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n738_), .A2(new_n528_), .A3(new_n410_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT51), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n745_), .A2(new_n749_), .A3(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1338gat));
  NAND3_X1  g550(.A1(new_n738_), .A2(new_n507_), .A3(new_n436_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n731_), .A2(new_n436_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G106gat), .B1(new_n666_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT114), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(G106gat), .C1(new_n666_), .C2(new_n753_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n755_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n756_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n754_), .A2(KEYINPUT114), .A3(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n752_), .A2(new_n759_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT53), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n752_), .A2(new_n759_), .A3(new_n764_), .A4(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1339gat));
  OAI21_X1  g565(.A(new_n573_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n539_), .B(new_n531_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT69), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n496_), .B1(new_n771_), .B2(new_n540_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n772_), .A2(new_n553_), .A3(new_n557_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n768_), .B1(new_n773_), .B2(KEYINPUT55), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n559_), .A2(KEYINPUT115), .A3(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n565_), .A2(new_n546_), .A3(new_n554_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n556_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n773_), .A2(KEYINPUT55), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n774_), .A2(new_n776_), .A3(new_n779_), .A4(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n778_), .A2(new_n777_), .B1(new_n773_), .B2(KEYINPUT55), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n784_), .A2(KEYINPUT116), .A3(new_n774_), .A4(new_n776_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n572_), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n787_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n767_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n475_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n469_), .A2(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n461_), .A2(new_n462_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n468_), .A2(new_n462_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n475_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n793_), .A2(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(new_n575_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n674_), .B1(new_n791_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  OR2_X1    g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n790_), .A2(KEYINPUT117), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n786_), .A2(new_n805_), .A3(new_n787_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n788_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n797_), .A2(new_n573_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n803_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n786_), .A2(new_n805_), .A3(new_n787_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n805_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n789_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n808_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(KEYINPUT58), .A3(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n809_), .A2(new_n605_), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n799_), .A2(new_n800_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n619_), .B1(new_n802_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n579_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n654_), .A2(new_n819_), .A3(new_n702_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT54), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n443_), .A2(new_n318_), .A3(new_n437_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(G113gat), .B1(new_n826_), .B2(new_n701_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n815_), .A2(new_n816_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n802_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n821_), .B1(new_n831_), .B2(new_n631_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n823_), .A2(KEYINPUT59), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n832_), .A2(new_n833_), .B1(new_n825_), .B2(KEYINPUT59), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n478_), .A2(new_n287_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n827_), .B1(new_n834_), .B2(new_n835_), .ZN(G1340gat));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT60), .B1(new_n579_), .B2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n825_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n834_), .A2(new_n840_), .A3(new_n579_), .ZN(new_n841_));
  OAI22_X1  g640(.A1(new_n841_), .A2(new_n837_), .B1(KEYINPUT60), .B2(new_n840_), .ZN(G1341gat));
  AOI21_X1  g641(.A(G127gat), .B1(new_n826_), .B2(new_n631_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n619_), .A2(new_n284_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n834_), .B2(new_n844_), .ZN(G1342gat));
  OAI21_X1  g644(.A(new_n285_), .B1(new_n825_), .B2(new_n632_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(KEYINPUT119), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n846_), .A2(KEYINPUT119), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT120), .B(G134gat), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n654_), .A2(new_n849_), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n847_), .B(new_n848_), .C1(new_n834_), .C2(new_n850_), .ZN(G1343gat));
  INV_X1    g650(.A(new_n822_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n852_), .A2(new_n647_), .A3(new_n410_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n318_), .A3(new_n713_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n478_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT121), .B(G141gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1344gat));
  NOR2_X1   g656(.A1(new_n854_), .A2(new_n819_), .ZN(new_n858_));
  INV_X1    g657(.A(G148gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1345gat));
  NOR2_X1   g659(.A1(new_n854_), .A2(new_n619_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT61), .B(G155gat), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n861_), .B(new_n863_), .ZN(G1346gat));
  NOR3_X1   g663(.A1(new_n854_), .A2(new_n595_), .A3(new_n654_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n854_), .A2(new_n632_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n595_), .ZN(G1347gat));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n820_), .B(KEYINPUT54), .Z(new_n869_));
  NAND2_X1  g668(.A1(new_n817_), .A2(KEYINPUT118), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n815_), .A2(new_n816_), .A3(new_n828_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(new_n801_), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n869_), .B1(new_n872_), .B2(new_n619_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n713_), .A2(new_n318_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n443_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n873_), .A2(new_n478_), .A3(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n324_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n868_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n878_), .ZN(new_n880_));
  OAI211_X1 g679(.A(KEYINPUT122), .B(KEYINPUT62), .C1(new_n876_), .C2(new_n324_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n879_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n873_), .A2(new_n875_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n701_), .A2(new_n342_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(KEYINPUT123), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n886_), .ZN(G1348gat));
  AOI21_X1  g686(.A(G176gat), .B1(new_n883_), .B2(new_n579_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n875_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n852_), .A2(new_n325_), .A3(new_n819_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n888_), .B1(new_n889_), .B2(new_n890_), .ZN(G1349gat));
  NOR3_X1   g690(.A1(new_n619_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n892_));
  INV_X1    g691(.A(G183gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n869_), .A2(new_n631_), .A3(new_n889_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n883_), .A2(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1350gat));
  INV_X1    g694(.A(new_n632_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n883_), .B(new_n896_), .C1(new_n334_), .C2(new_n333_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n832_), .A2(new_n605_), .A3(new_n889_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n898_), .A2(new_n899_), .A3(G190gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(G190gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n897_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(KEYINPUT125), .B(new_n897_), .C1(new_n900_), .C2(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1351gat));
  NAND3_X1  g705(.A1(new_n853_), .A2(new_n701_), .A3(new_n874_), .ZN(new_n907_));
  OR3_X1    g706(.A1(new_n907_), .A2(KEYINPUT126), .A3(new_n474_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n474_), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT126), .B1(new_n907_), .B2(new_n474_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n908_), .A2(new_n909_), .A3(new_n910_), .ZN(G1352gat));
  AND2_X1   g710(.A1(new_n853_), .A2(new_n874_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n579_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g713(.A(KEYINPUT63), .B(G211gat), .C1(new_n912_), .C2(new_n631_), .ZN(new_n915_));
  XOR2_X1   g714(.A(KEYINPUT63), .B(G211gat), .Z(new_n916_));
  AND3_X1   g715(.A1(new_n912_), .A2(new_n631_), .A3(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n915_), .A2(new_n917_), .ZN(G1354gat));
  AOI21_X1  g717(.A(G218gat), .B1(new_n912_), .B2(new_n896_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n605_), .A2(G218gat), .ZN(new_n920_));
  XOR2_X1   g719(.A(new_n920_), .B(KEYINPUT127), .Z(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n912_), .B2(new_n921_), .ZN(G1355gat));
endmodule


