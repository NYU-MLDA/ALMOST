//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n985_, new_n987_, new_n988_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1013_,
    new_n1014_, new_n1015_, new_n1017_, new_n1018_, new_n1020_, new_n1021_,
    new_n1023_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT87), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT29), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT85), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT1), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n210_), .B2(KEYINPUT1), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT84), .ZN(new_n215_));
  INV_X1    g014(.A(G155gat), .ZN(new_n216_));
  INV_X1    g015(.A(G162gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n220_));
  AND2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n218_), .A2(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n209_), .B1(new_n214_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224_));
  INV_X1    g023(.A(G141gat), .ZN(new_n225_));
  INV_X1    g024(.A(G148gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n205_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n227_), .A2(new_n229_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n218_), .A2(new_n219_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n210_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT86), .B1(new_n223_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT85), .B1(new_n221_), .B2(new_n220_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT1), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n221_), .A2(new_n220_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n219_), .ZN(new_n240_));
  NOR3_X1   g039(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n208_), .B1(new_n238_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT86), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n232_), .A2(new_n233_), .A3(new_n210_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n204_), .B1(new_n235_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT88), .ZN(new_n248_));
  INV_X1    g047(.A(G197gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n248_), .B1(new_n249_), .B2(G204gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G211gat), .A2(G218gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G211gat), .A2(G218gat), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n252_), .A2(new_n253_), .A3(KEYINPUT89), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT89), .ZN(new_n255_));
  INV_X1    g054(.A(G211gat), .ZN(new_n256_));
  INV_X1    g055(.A(G218gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n255_), .B1(new_n258_), .B2(new_n251_), .ZN(new_n259_));
  OAI211_X1 g058(.A(KEYINPUT21), .B(new_n250_), .C1(new_n254_), .C2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G197gat), .B(G204gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT89), .B1(new_n252_), .B2(new_n253_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n258_), .A2(new_n255_), .A3(new_n251_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n265_), .A2(KEYINPUT21), .ZN(new_n266_));
  INV_X1    g065(.A(new_n261_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n265_), .A2(KEYINPUT21), .A3(new_n267_), .A4(new_n250_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n262_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n203_), .B1(new_n247_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT29), .B1(new_n223_), .B2(new_n234_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT90), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n203_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n269_), .A2(KEYINPUT91), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT91), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n262_), .A2(new_n266_), .A3(new_n275_), .A4(new_n268_), .ZN(new_n276_));
  OAI211_X1 g075(.A(KEYINPUT90), .B(KEYINPUT29), .C1(new_n223_), .C2(new_n234_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n273_), .A2(new_n274_), .A3(new_n276_), .A4(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G78gat), .B(G106gat), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n270_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n279_), .B1(new_n270_), .B2(new_n278_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT92), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n270_), .A2(new_n278_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n279_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT92), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n270_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n235_), .A2(new_n204_), .A3(new_n246_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n289_), .A2(G50gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT28), .B(G22gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(G50gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n292_), .B1(new_n290_), .B2(new_n293_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n282_), .A2(new_n288_), .A3(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n289_), .B(G50gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n291_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n294_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n301_), .B(KEYINPUT92), .C1(new_n280_), .C2(new_n281_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n298_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G226gat), .A2(G233gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT19), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n309_));
  NOR2_X1   g108(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(KEYINPUT23), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n306_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G176gat), .ZN(new_n314_));
  AND2_X1   g113(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n313_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n307_), .A2(KEYINPUT23), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n309_), .A2(new_n310_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n321_), .B1(new_n322_), .B2(new_n307_), .ZN(new_n323_));
  INV_X1    g122(.A(G190gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(KEYINPUT26), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(KEYINPUT74), .A3(KEYINPUT75), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(KEYINPUT26), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT26), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(G190gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n327_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n327_), .B1(new_n329_), .B2(G190gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n326_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n336_));
  NOR2_X1   g135(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n323_), .B1(new_n335_), .B2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT24), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n318_), .A2(KEYINPUT24), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n342_), .B1(new_n343_), .B2(new_n340_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n320_), .B1(new_n339_), .B2(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n346_), .A2(new_n269_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n310_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n307_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n321_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n306_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n319_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT26), .B(G190gat), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n338_), .A2(new_n355_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n353_), .A2(new_n354_), .B1(new_n356_), .B2(new_n345_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT20), .B1(new_n269_), .B2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n305_), .B1(new_n347_), .B2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n305_), .B1(new_n269_), .B2(new_n357_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n360_), .B(KEYINPUT20), .C1(new_n269_), .C2(new_n346_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT18), .B(G64gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(G92gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  NAND3_X1  g164(.A1(new_n359_), .A2(new_n361_), .A3(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n366_), .A2(KEYINPUT27), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n338_), .A2(new_n355_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n311_), .A2(new_n312_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  OAI22_X1  g169(.A1(new_n370_), .A2(new_n344_), .B1(new_n352_), .B2(new_n319_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT20), .B1(new_n346_), .B2(new_n269_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n305_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n346_), .A2(new_n269_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n305_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n371_), .A2(new_n262_), .A3(new_n266_), .A4(new_n268_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n375_), .A2(KEYINPUT20), .A3(new_n376_), .A4(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT95), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n262_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(new_n371_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n383_), .A2(KEYINPUT95), .A3(new_n376_), .A4(new_n375_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n374_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n365_), .B(KEYINPUT97), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n365_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n376_), .B1(new_n383_), .B2(new_n375_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n376_), .B1(new_n382_), .B2(new_n371_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(new_n373_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n388_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n366_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT27), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n367_), .A2(new_n387_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n303_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT98), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n303_), .A2(KEYINPUT98), .A3(new_n395_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G227gat), .A2(G233gat), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n401_), .B(KEYINPUT77), .Z(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G71gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G15gat), .B(G43gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n350_), .A2(new_n351_), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n330_), .A2(new_n327_), .A3(new_n333_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n329_), .A2(G190gat), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT74), .B1(new_n409_), .B2(new_n325_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT75), .B1(new_n328_), .B2(new_n327_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n338_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n345_), .B(new_n407_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT30), .ZN(new_n415_));
  INV_X1    g214(.A(new_n320_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n415_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n417_), .A2(new_n418_), .A3(G99gat), .ZN(new_n419_));
  INV_X1    g218(.A(G99gat), .ZN(new_n420_));
  AOI211_X1 g219(.A(new_n344_), .B(new_n323_), .C1(new_n335_), .C2(new_n338_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT30), .B1(new_n421_), .B2(new_n320_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n414_), .A2(new_n416_), .A3(new_n415_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n420_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n406_), .B1(new_n419_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G113gat), .B(G120gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G127gat), .A2(G134gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G127gat), .A2(G134gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT79), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  OR2_X1    g230(.A1(G127gat), .A2(G134gat), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT79), .B1(new_n432_), .B2(new_n427_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n426_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT80), .ZN(new_n435_));
  INV_X1    g234(.A(new_n426_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n430_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n432_), .A2(KEYINPUT79), .A3(new_n427_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n434_), .A2(new_n435_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT81), .ZN(new_n441_));
  OAI211_X1 g240(.A(KEYINPUT80), .B(new_n426_), .C1(new_n431_), .C2(new_n433_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT31), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n441_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n440_), .A2(new_n442_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT81), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT31), .B1(new_n449_), .B2(new_n443_), .ZN(new_n450_));
  OAI22_X1  g249(.A1(new_n447_), .A2(new_n450_), .B1(KEYINPUT78), .B2(KEYINPUT82), .ZN(new_n451_));
  OAI21_X1  g250(.A(G99gat), .B1(new_n417_), .B2(new_n418_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n422_), .A2(new_n420_), .A3(new_n423_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n453_), .A3(new_n405_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n425_), .A2(new_n451_), .A3(new_n454_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n452_), .A2(new_n453_), .A3(new_n405_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n405_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT82), .B1(new_n447_), .B2(new_n450_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n445_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n449_), .A2(KEYINPUT31), .A3(new_n443_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(KEYINPUT78), .A3(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n455_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT83), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n467_), .B(new_n455_), .C1(new_n458_), .C2(new_n464_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n244_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n448_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT4), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G225gat), .A2(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n434_), .A2(new_n439_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n476_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n235_), .A2(new_n246_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n477_), .B1(new_n478_), .B2(new_n448_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n473_), .B(new_n475_), .C1(new_n479_), .C2(new_n472_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n235_), .A2(new_n246_), .B1(new_n442_), .B2(new_n440_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n474_), .B1(new_n481_), .B2(new_n477_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT0), .B(G57gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(G85gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(G1gat), .B(G29gat), .Z(new_n485_));
  XOR2_X1   g284(.A(new_n484_), .B(new_n485_), .Z(new_n486_));
  NAND3_X1  g285(.A1(new_n480_), .A2(new_n482_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT96), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n486_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n480_), .A2(new_n482_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n486_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(KEYINPUT96), .A3(new_n487_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n466_), .A2(new_n468_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n466_), .A2(new_n468_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n493_), .B1(KEYINPUT96), .B2(new_n487_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n488_), .A2(new_n489_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n395_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n303_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n496_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT93), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT33), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n503_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n504_));
  AOI211_X1 g303(.A(KEYINPUT33), .B(new_n486_), .C1(new_n480_), .C2(new_n482_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT4), .B1(new_n481_), .B2(new_n477_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n475_), .B1(new_n507_), .B2(new_n473_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n481_), .A2(new_n477_), .A3(new_n474_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n486_), .A3(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(new_n366_), .A3(new_n392_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n502_), .B1(new_n506_), .B2(new_n513_), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n508_), .A2(new_n492_), .A3(new_n510_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n393_), .A2(new_n515_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n516_), .B(KEYINPUT93), .C1(new_n504_), .C2(new_n505_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n365_), .A2(KEYINPUT32), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n359_), .A2(new_n361_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT94), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(KEYINPUT32), .B(new_n365_), .C1(new_n519_), .C2(KEYINPUT94), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n521_), .B1(new_n522_), .B2(new_n385_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(new_n490_), .A3(new_n494_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n514_), .A2(new_n517_), .A3(new_n303_), .A4(new_n524_), .ZN(new_n525_));
  AOI22_X1  g324(.A1(new_n400_), .A2(new_n495_), .B1(new_n501_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT9), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT9), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT64), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G99gat), .A2(G106gat), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT6), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT10), .B(G99gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(G106gat), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n539_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT64), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n530_), .A2(new_n544_), .A3(new_n532_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n534_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT65), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n547_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n548_));
  OR2_X1    g347(.A1(G85gat), .A2(G92gat), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(KEYINPUT65), .A3(new_n527_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT8), .ZN(new_n552_));
  OR3_X1    g351(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n553_), .A2(new_n537_), .A3(new_n538_), .A4(new_n554_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n551_), .A2(new_n552_), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n552_), .B1(new_n551_), .B2(new_n555_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n546_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(G57gat), .ZN(new_n559_));
  INV_X1    g358(.A(G64gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G57gat), .A2(G64gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT11), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G71gat), .B(G78gat), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT11), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n561_), .A2(new_n567_), .A3(new_n562_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n564_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n563_), .A2(new_n565_), .A3(KEYINPUT11), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT66), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n558_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n575_), .B1(new_n558_), .B2(new_n572_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n546_), .B(new_n571_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n574_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n576_), .A2(new_n577_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G230gat), .A2(G233gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n558_), .A2(new_n572_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n578_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n582_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(G120gat), .B(G148gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(G204gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT5), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(new_n314_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n583_), .A2(new_n587_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT67), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n583_), .A2(KEYINPUT67), .A3(new_n587_), .A4(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n583_), .A2(new_n587_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n591_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT13), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n596_), .A2(new_n602_), .A3(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G15gat), .B(G22gat), .ZN(new_n605_));
  INV_X1    g404(.A(G1gat), .ZN(new_n606_));
  INV_X1    g405(.A(G8gat), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT14), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G1gat), .B(G8gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n609_), .B(new_n610_), .Z(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(G43gat), .B(G50gat), .Z(new_n613_));
  XOR2_X1   g412(.A(G29gat), .B(G36gat), .Z(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G43gat), .B(G50gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G29gat), .B(G36gat), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n615_), .A2(new_n616_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n616_), .B1(new_n615_), .B2(new_n619_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n612_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n615_), .A2(new_n619_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n616_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n615_), .A2(new_n616_), .A3(new_n619_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n611_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n623_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G229gat), .A2(G233gat), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT15), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n634_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n626_), .A2(KEYINPUT15), .A3(new_n627_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n631_), .B(new_n629_), .C1(new_n637_), .C2(new_n611_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G113gat), .B(G141gat), .ZN(new_n639_));
  INV_X1    g438(.A(G169gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(new_n249_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n633_), .A2(new_n638_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n643_), .B1(new_n633_), .B2(new_n638_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n604_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT72), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT37), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT73), .Z(new_n652_));
  INV_X1    g451(.A(KEYINPUT71), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT70), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n654_), .B1(new_n558_), .B2(new_n622_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(G232gat), .A2(G233gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT34), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(KEYINPUT35), .A3(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n628_), .B(new_n546_), .C1(new_n557_), .C2(new_n556_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n657_), .A2(KEYINPUT35), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n558_), .A2(new_n636_), .A3(new_n635_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n664_), .A2(KEYINPUT35), .A3(new_n657_), .A4(new_n655_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n653_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(G190gat), .B(G218gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(G134gat), .B(G162gat), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n663_), .A2(new_n665_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(KEYINPUT36), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT36), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n669_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n666_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n671_), .A2(KEYINPUT71), .ZN(new_n676_));
  INV_X1    g475(.A(new_n674_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n673_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n676_), .B(new_n677_), .C1(new_n678_), .C2(new_n670_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n675_), .A2(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n650_), .A2(KEYINPUT37), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n652_), .B1(new_n680_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n652_), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n681_), .B(new_n684_), .C1(new_n675_), .C2(new_n679_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n611_), .B(new_n571_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(G231gat), .A2(G233gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT17), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT16), .B(G183gat), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(G211gat), .ZN(new_n693_));
  XOR2_X1   g492(.A(G127gat), .B(G155gat), .Z(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  OR3_X1    g494(.A1(new_n690_), .A2(new_n691_), .A3(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(KEYINPUT17), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n690_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  NOR4_X1   g498(.A1(new_n526_), .A2(new_n649_), .A3(new_n686_), .A4(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n497_), .A2(new_n498_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n606_), .A3(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT38), .ZN(new_n703_));
  OR3_X1    g502(.A1(new_n649_), .A2(KEYINPUT99), .A3(new_n699_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT99), .B1(new_n649_), .B2(new_n699_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n501_), .A2(new_n525_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n303_), .A2(KEYINPUT98), .A3(new_n395_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT98), .B1(new_n303_), .B2(new_n395_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n495_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT100), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n658_), .B(new_n664_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n669_), .B1(new_n712_), .B2(new_n673_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n676_), .B1(new_n713_), .B2(new_n677_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n672_), .A2(new_n666_), .A3(new_n674_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n711_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n675_), .A2(KEYINPUT100), .A3(new_n679_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n704_), .A2(new_n705_), .A3(new_n710_), .A4(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n701_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G1gat), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n703_), .A2(new_n721_), .ZN(G1324gat));
  AND3_X1   g521(.A1(new_n704_), .A2(new_n710_), .A3(new_n718_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n724_));
  INV_X1    g523(.A(new_n395_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n723_), .A2(new_n724_), .A3(new_n705_), .A4(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT101), .B1(new_n719_), .B2(new_n395_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(G8gat), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT39), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT39), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n726_), .A2(new_n730_), .A3(new_n727_), .A4(G8gat), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n700_), .A2(new_n607_), .A3(new_n725_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT40), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n732_), .A2(KEYINPUT40), .A3(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1325gat));
  INV_X1    g537(.A(new_n496_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G15gat), .B1(new_n719_), .B2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT41), .Z(new_n741_));
  INV_X1    g540(.A(G15gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n700_), .A2(new_n742_), .A3(new_n496_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1326gat));
  OAI21_X1  g543(.A(G22gat), .B1(new_n719_), .B2(new_n303_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT42), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n303_), .A2(G22gat), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT102), .Z(new_n748_));
  NAND2_X1  g547(.A1(new_n700_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n746_), .A2(new_n749_), .ZN(G1327gat));
  NAND3_X1  g549(.A1(new_n604_), .A2(new_n648_), .A3(new_n699_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n683_), .A2(new_n685_), .ZN(new_n752_));
  OAI21_X1  g551(.A(KEYINPUT43), .B1(new_n526_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n710_), .A2(new_n754_), .A3(new_n686_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n751_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n756_), .B2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(G29gat), .A3(new_n701_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n751_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n717_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT100), .B1(new_n675_), .B2(new_n679_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(new_n710_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT104), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n762_), .A2(new_n710_), .A3(new_n768_), .A4(new_n765_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n720_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n761_), .B1(G29gat), .B2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT105), .ZN(G1328gat));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n775_));
  INV_X1    g574(.A(G36gat), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n767_), .A2(new_n776_), .A3(new_n725_), .A4(new_n769_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(KEYINPUT106), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(KEYINPUT106), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n753_), .A2(new_n755_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n781_), .A2(new_n762_), .A3(new_n757_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n759_), .B1(new_n781_), .B2(new_n762_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n725_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(G36gat), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT106), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n770_), .A2(new_n786_), .A3(new_n776_), .A4(new_n725_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n777_), .A2(KEYINPUT106), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(KEYINPUT45), .A3(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n780_), .A2(new_n785_), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n790_), .B(new_n791_), .ZN(G1329gat));
  OAI211_X1 g591(.A(G43gat), .B(new_n496_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT107), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n760_), .A2(KEYINPUT107), .A3(G43gat), .A4(new_n496_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT108), .B(G43gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n771_), .B2(new_n739_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n796_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT47), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n795_), .A2(new_n796_), .A3(new_n801_), .A4(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1330gat));
  INV_X1    g602(.A(G50gat), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n770_), .A2(new_n804_), .A3(new_n500_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n760_), .A2(new_n500_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n804_), .ZN(G1331gat));
  INV_X1    g606(.A(new_n604_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n699_), .A2(new_n648_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n710_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n718_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n811_), .A2(new_n559_), .A3(new_n720_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n752_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n813_), .A2(KEYINPUT109), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(KEYINPUT109), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n701_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n812_), .B1(new_n816_), .B2(new_n559_), .ZN(new_n817_));
  XOR2_X1   g616(.A(new_n817_), .B(KEYINPUT110), .Z(G1332gat));
  OAI21_X1  g617(.A(G64gat), .B1(new_n811_), .B2(new_n395_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT48), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n725_), .A2(new_n560_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n813_), .B2(new_n821_), .ZN(G1333gat));
  OR3_X1    g621(.A1(new_n813_), .A2(G71gat), .A3(new_n739_), .ZN(new_n823_));
  OAI21_X1  g622(.A(G71gat), .B1(new_n811_), .B2(new_n739_), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n824_), .A2(KEYINPUT111), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(KEYINPUT111), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n825_), .A2(KEYINPUT49), .A3(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT49), .B1(new_n825_), .B2(new_n826_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n823_), .B1(new_n827_), .B2(new_n828_), .ZN(G1334gat));
  OAI21_X1  g628(.A(G78gat), .B1(new_n811_), .B2(new_n303_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT50), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n303_), .A2(G78gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n813_), .B2(new_n832_), .ZN(G1335gat));
  NOR2_X1   g632(.A1(new_n526_), .A2(new_n718_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n699_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n604_), .A2(new_n648_), .A3(new_n835_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(G85gat), .B1(new_n837_), .B2(new_n701_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n710_), .A2(new_n754_), .A3(new_n686_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n754_), .B1(new_n710_), .B2(new_n686_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT112), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n836_), .B(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n753_), .A2(new_n844_), .A3(new_n755_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n841_), .A2(new_n843_), .A3(new_n845_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n846_), .A2(G85gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n838_), .B1(new_n847_), .B2(new_n701_), .ZN(G1336gat));
  AOI21_X1  g647(.A(G92gat), .B1(new_n837_), .B2(new_n725_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n846_), .A2(new_n725_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(G92gat), .ZN(G1337gat));
  NAND4_X1  g650(.A1(new_n841_), .A2(new_n496_), .A3(new_n843_), .A4(new_n845_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n852_), .A2(KEYINPUT114), .A3(G99gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT114), .B1(new_n852_), .B2(G99gat), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n834_), .A2(new_n541_), .A3(new_n496_), .A4(new_n836_), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(KEYINPUT115), .Z(new_n857_));
  NAND4_X1  g656(.A1(new_n855_), .A2(KEYINPUT116), .A3(KEYINPUT51), .A4(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n852_), .A2(G99gat), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n852_), .A2(KEYINPUT114), .A3(G99gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n857_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n864_));
  OR2_X1    g663(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n858_), .A2(new_n866_), .ZN(G1338gat));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n781_), .A2(new_n500_), .A3(new_n843_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(G106gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n869_), .B2(G106gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n868_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n873_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(KEYINPUT52), .A3(new_n871_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n837_), .A2(new_n542_), .A3(new_n500_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n874_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT53), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n874_), .A2(new_n876_), .A3(new_n880_), .A4(new_n877_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(G1339gat));
  NOR2_X1   g681(.A1(new_n739_), .A2(new_n720_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n647_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT55), .B1(new_n581_), .B2(new_n582_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n583_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n575_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n584_), .A2(new_n887_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n578_), .A2(new_n579_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n558_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT55), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n586_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n886_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(KEYINPUT56), .B1(new_n895_), .B2(new_n598_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n897_));
  AOI211_X1 g696(.A(new_n897_), .B(new_n591_), .C1(new_n886_), .C2(new_n894_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n884_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n630_), .A2(new_n631_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n632_), .B(new_n629_), .C1(new_n637_), .C2(new_n611_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n900_), .A2(new_n901_), .A3(new_n642_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n902_), .A2(new_n903_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n904_), .A2(new_n905_), .A3(new_n645_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n600_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n899_), .A2(new_n907_), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n908_), .A2(new_n718_), .A3(KEYINPUT57), .ZN(new_n909_));
  AOI21_X1  g708(.A(KEYINPUT57), .B1(new_n908_), .B2(new_n718_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n892_), .B1(new_n891_), .B2(new_n586_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n891_), .A2(new_n586_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n598_), .B1(new_n915_), .B2(new_n893_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n897_), .ZN(new_n917_));
  OAI211_X1 g716(.A(KEYINPUT56), .B(new_n598_), .C1(new_n915_), .C2(new_n893_), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n917_), .A2(KEYINPUT119), .A3(new_n918_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n906_), .B(new_n596_), .C1(new_n918_), .C2(KEYINPUT119), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n912_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n920_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n917_), .A2(KEYINPUT119), .A3(new_n918_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n922_), .A2(KEYINPUT58), .A3(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n686_), .A2(new_n921_), .A3(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n835_), .B1(new_n911_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n752_), .A2(new_n927_), .A3(new_n604_), .A4(new_n809_), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n604_), .B(new_n809_), .C1(new_n683_), .C2(new_n685_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(KEYINPUT54), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n928_), .A2(new_n930_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n400_), .B(new_n883_), .C1(new_n926_), .C2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(G113gat), .B1(new_n933_), .B2(new_n648_), .ZN(new_n934_));
  OR2_X1    g733(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n935_));
  NAND2_X1  g734(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n932_), .A2(new_n935_), .A3(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n400_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT57), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n917_), .A2(new_n918_), .ZN(new_n940_));
  AOI22_X1  g739(.A1(new_n940_), .A2(new_n884_), .B1(new_n600_), .B2(new_n906_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n939_), .B1(new_n765_), .B2(new_n941_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n908_), .A2(new_n718_), .A3(KEYINPUT57), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n925_), .A2(new_n942_), .A3(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n699_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n928_), .A2(new_n930_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n938_), .B1(new_n945_), .B2(new_n946_), .ZN(new_n947_));
  NAND4_X1  g746(.A1(new_n947_), .A2(KEYINPUT120), .A3(KEYINPUT59), .A4(new_n883_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n647_), .B1(new_n937_), .B2(new_n948_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n934_), .B1(new_n949_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g749(.A(G120gat), .ZN(new_n951_));
  OR2_X1    g750(.A1(new_n951_), .A2(KEYINPUT60), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n604_), .B2(KEYINPUT60), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n933_), .A2(new_n952_), .A3(new_n953_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(KEYINPUT121), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n604_), .B1(new_n937_), .B2(new_n948_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n951_), .B2(new_n956_), .ZN(G1341gat));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n958_));
  INV_X1    g757(.A(G127gat), .ZN(new_n959_));
  AOI211_X1 g758(.A(new_n959_), .B(new_n699_), .C1(new_n937_), .C2(new_n948_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT122), .ZN(new_n961_));
  AOI22_X1  g760(.A1(new_n944_), .A2(new_n699_), .B1(new_n928_), .B2(new_n930_), .ZN(new_n962_));
  INV_X1    g761(.A(new_n883_), .ZN(new_n963_));
  NOR4_X1   g762(.A1(new_n962_), .A2(new_n699_), .A3(new_n938_), .A4(new_n963_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n961_), .B1(new_n964_), .B2(G127gat), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n947_), .A2(new_n835_), .A3(new_n883_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n966_), .A2(KEYINPUT122), .A3(new_n959_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n965_), .A2(new_n967_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n958_), .B1(new_n960_), .B2(new_n968_), .ZN(new_n969_));
  NOR3_X1   g768(.A1(new_n964_), .A2(new_n961_), .A3(G127gat), .ZN(new_n970_));
  AOI21_X1  g769(.A(KEYINPUT122), .B1(new_n966_), .B2(new_n959_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n970_), .A2(new_n971_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n937_), .A2(new_n948_), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n973_), .A2(G127gat), .A3(new_n835_), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n972_), .A2(new_n974_), .A3(KEYINPUT123), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n969_), .A2(new_n975_), .ZN(G1342gat));
  AOI21_X1  g775(.A(G134gat), .B1(new_n933_), .B2(new_n765_), .ZN(new_n977_));
  AND2_X1   g776(.A1(new_n973_), .A2(G134gat), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n977_), .B1(new_n978_), .B2(new_n686_), .ZN(G1343gat));
  NAND2_X1  g778(.A1(new_n739_), .A2(new_n500_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n962_), .A2(new_n980_), .ZN(new_n981_));
  NAND3_X1  g780(.A1(new_n981_), .A2(new_n701_), .A3(new_n395_), .ZN(new_n982_));
  NOR2_X1   g781(.A1(new_n982_), .A2(new_n647_), .ZN(new_n983_));
  XNOR2_X1  g782(.A(new_n983_), .B(new_n225_), .ZN(G1344gat));
  NOR2_X1   g783(.A1(new_n982_), .A2(new_n604_), .ZN(new_n985_));
  XNOR2_X1  g784(.A(new_n985_), .B(new_n226_), .ZN(G1345gat));
  NOR2_X1   g785(.A1(new_n982_), .A2(new_n699_), .ZN(new_n987_));
  XOR2_X1   g786(.A(KEYINPUT61), .B(G155gat), .Z(new_n988_));
  XNOR2_X1  g787(.A(new_n987_), .B(new_n988_), .ZN(G1346gat));
  NOR3_X1   g788(.A1(new_n982_), .A2(new_n217_), .A3(new_n752_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n217_), .B1(new_n982_), .B2(new_n718_), .ZN(new_n991_));
  INV_X1    g790(.A(KEYINPUT124), .ZN(new_n992_));
  OR2_X1    g791(.A1(new_n991_), .A2(new_n992_), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n991_), .A2(new_n992_), .ZN(new_n994_));
  AOI21_X1  g793(.A(new_n990_), .B1(new_n993_), .B2(new_n994_), .ZN(G1347gat));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n996_));
  OAI21_X1  g795(.A(new_n303_), .B1(new_n926_), .B2(new_n931_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n495_), .A2(new_n725_), .ZN(new_n998_));
  NOR2_X1   g797(.A1(new_n997_), .A2(new_n998_), .ZN(new_n999_));
  NAND2_X1  g798(.A1(new_n999_), .A2(new_n648_), .ZN(new_n1000_));
  AOI21_X1  g799(.A(new_n996_), .B1(new_n1000_), .B2(G169gat), .ZN(new_n1001_));
  AOI211_X1 g800(.A(KEYINPUT62), .B(new_n640_), .C1(new_n999_), .C2(new_n648_), .ZN(new_n1002_));
  INV_X1    g801(.A(new_n999_), .ZN(new_n1003_));
  OAI21_X1  g802(.A(new_n648_), .B1(new_n316_), .B2(new_n315_), .ZN(new_n1004_));
  XOR2_X1   g803(.A(new_n1004_), .B(KEYINPUT125), .Z(new_n1005_));
  OAI22_X1  g804(.A1(new_n1001_), .A2(new_n1002_), .B1(new_n1003_), .B2(new_n1005_), .ZN(G1348gat));
  AOI21_X1  g805(.A(G176gat), .B1(new_n999_), .B2(new_n808_), .ZN(new_n1007_));
  OR2_X1    g806(.A1(new_n997_), .A2(KEYINPUT126), .ZN(new_n1008_));
  INV_X1    g807(.A(new_n998_), .ZN(new_n1009_));
  NAND2_X1  g808(.A1(new_n997_), .A2(KEYINPUT126), .ZN(new_n1010_));
  AND4_X1   g809(.A1(G176gat), .A2(new_n1008_), .A3(new_n1009_), .A4(new_n1010_), .ZN(new_n1011_));
  AOI21_X1  g810(.A(new_n1007_), .B1(new_n1011_), .B2(new_n808_), .ZN(G1349gat));
  NOR3_X1   g811(.A1(new_n1003_), .A2(new_n699_), .A3(new_n338_), .ZN(new_n1013_));
  NAND4_X1  g812(.A1(new_n1008_), .A2(new_n835_), .A3(new_n1009_), .A4(new_n1010_), .ZN(new_n1014_));
  INV_X1    g813(.A(G183gat), .ZN(new_n1015_));
  AOI21_X1  g814(.A(new_n1013_), .B1(new_n1014_), .B2(new_n1015_), .ZN(G1350gat));
  OAI21_X1  g815(.A(G190gat), .B1(new_n1003_), .B2(new_n752_), .ZN(new_n1017_));
  NAND3_X1  g816(.A1(new_n999_), .A2(new_n355_), .A3(new_n765_), .ZN(new_n1018_));
  NAND2_X1  g817(.A1(new_n1017_), .A2(new_n1018_), .ZN(G1351gat));
  NOR4_X1   g818(.A1(new_n962_), .A2(new_n701_), .A3(new_n395_), .A4(new_n980_), .ZN(new_n1020_));
  NAND2_X1  g819(.A1(new_n1020_), .A2(new_n648_), .ZN(new_n1021_));
  XNOR2_X1  g820(.A(new_n1021_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g821(.A1(new_n1020_), .A2(new_n808_), .ZN(new_n1023_));
  XNOR2_X1  g822(.A(new_n1023_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g823(.A1(new_n1020_), .A2(new_n835_), .ZN(new_n1025_));
  NOR2_X1   g824(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1026_));
  AND2_X1   g825(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1027_));
  NOR3_X1   g826(.A1(new_n1025_), .A2(new_n1026_), .A3(new_n1027_), .ZN(new_n1028_));
  AOI21_X1  g827(.A(new_n1028_), .B1(new_n1025_), .B2(new_n1026_), .ZN(G1354gat));
  INV_X1    g828(.A(new_n1020_), .ZN(new_n1030_));
  OAI21_X1  g829(.A(new_n257_), .B1(new_n1030_), .B2(new_n718_), .ZN(new_n1031_));
  NAND3_X1  g830(.A1(new_n1020_), .A2(G218gat), .A3(new_n686_), .ZN(new_n1032_));
  NAND2_X1  g831(.A1(new_n1031_), .A2(new_n1032_), .ZN(new_n1033_));
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1034_));
  NAND2_X1  g833(.A1(new_n1033_), .A2(new_n1034_), .ZN(new_n1035_));
  NAND3_X1  g834(.A1(new_n1031_), .A2(KEYINPUT127), .A3(new_n1032_), .ZN(new_n1036_));
  NAND2_X1  g835(.A1(new_n1035_), .A2(new_n1036_), .ZN(G1355gat));
endmodule


