//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT68), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n208_));
  INV_X1    g007(.A(G99gat), .ZN(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT7), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT6), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G99gat), .A3(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n208_), .A2(new_n218_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n212_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT65), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n212_), .A2(new_n217_), .A3(new_n222_), .A4(new_n219_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G85gat), .B(G92gat), .Z(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT66), .B(KEYINPUT8), .Z(new_n225_));
  AND2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n221_), .A2(new_n223_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n220_), .A2(new_n228_), .A3(new_n224_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT8), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n220_), .B2(new_n224_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n227_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT10), .B(G99gat), .Z(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(new_n210_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n224_), .A2(KEYINPUT9), .ZN(new_n235_));
  INV_X1    g034(.A(G85gat), .ZN(new_n236_));
  INV_X1    g035(.A(G92gat), .ZN(new_n237_));
  OR3_X1    g036(.A1(new_n236_), .A2(new_n237_), .A3(KEYINPUT9), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n234_), .A2(new_n235_), .A3(new_n217_), .A4(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n232_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G64gat), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n243_));
  XOR2_X1   g042(.A(G71gat), .B(G78gat), .Z(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n243_), .A2(new_n244_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n240_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n232_), .A2(new_n247_), .A3(new_n239_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G230gat), .A2(G233gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n207_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n232_), .A2(new_n247_), .A3(new_n239_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n247_), .B1(new_n232_), .B2(new_n239_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n207_), .B(new_n253_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT12), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n255_), .A2(new_n256_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n260_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n252_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n206_), .B1(new_n259_), .B2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n253_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT68), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n264_), .A2(new_n257_), .A3(new_n267_), .A4(new_n206_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n259_), .A2(KEYINPUT69), .A3(new_n264_), .A4(new_n206_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n265_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n272_), .A2(KEYINPUT13), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(KEYINPUT13), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G15gat), .B(G22gat), .ZN(new_n275_));
  INV_X1    g074(.A(G1gat), .ZN(new_n276_));
  INV_X1    g075(.A(G8gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT14), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G8gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n247_), .B(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G231gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT17), .ZN(new_n285_));
  XOR2_X1   g084(.A(G127gat), .B(G155gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT16), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G183gat), .B(G211gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  OR3_X1    g088(.A1(new_n284_), .A2(new_n285_), .A3(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(KEYINPUT17), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n284_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G190gat), .B(G218gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT71), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G134gat), .B(G162gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT36), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G232gat), .A2(G233gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT34), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT35), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n239_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n220_), .A2(new_n224_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT67), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(KEYINPUT8), .A3(new_n229_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n307_), .B1(new_n310_), .B2(new_n227_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G29gat), .B(G36gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G43gat), .B(G50gat), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n313_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n311_), .A2(new_n316_), .B1(new_n304_), .B2(new_n303_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n314_), .A2(new_n315_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT15), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n311_), .A2(new_n319_), .A3(KEYINPUT70), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n316_), .B(KEYINPUT15), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n321_), .B1(new_n240_), .B2(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n306_), .B(new_n317_), .C1(new_n320_), .C2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT70), .B1(new_n311_), .B2(new_n319_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n240_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n306_), .B1(new_n328_), .B2(new_n317_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n300_), .B1(new_n325_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT37), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n317_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n305_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n298_), .A2(KEYINPUT36), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n335_), .A3(new_n324_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n330_), .A2(new_n331_), .A3(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n299_), .B(KEYINPUT72), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n325_), .B2(new_n329_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n331_), .B1(new_n339_), .B2(new_n336_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n294_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n273_), .A2(new_n274_), .A3(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT73), .ZN(new_n343_));
  XOR2_X1   g142(.A(G127gat), .B(G134gat), .Z(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT83), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G127gat), .B(G134gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT83), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G113gat), .B(G120gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n345_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(KEYINPUT84), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G141gat), .A2(G148gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT2), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n361_));
  OAI22_X1  g160(.A1(new_n361_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n357_), .A2(new_n360_), .A3(new_n362_), .A4(new_n363_), .ZN(new_n364_));
  OR2_X1    g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n355_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n368_), .A2(new_n358_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(KEYINPUT1), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT1), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(G155gat), .A3(G162gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n372_), .A3(new_n365_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n364_), .A2(new_n367_), .B1(new_n369_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT97), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n354_), .A2(new_n375_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n352_), .A2(KEYINPUT97), .A3(new_n374_), .A4(new_n353_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(KEYINPUT4), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n364_), .A2(new_n367_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n369_), .A2(new_n373_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n354_), .A2(new_n381_), .A3(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n378_), .A2(new_n380_), .A3(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G85gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT0), .B(G57gat), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n388_), .B(new_n389_), .Z(new_n390_));
  NAND3_X1  g189(.A1(new_n376_), .A2(new_n379_), .A3(new_n377_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n386_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n390_), .B1(new_n386_), .B2(new_n391_), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(G176gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT22), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(G169gat), .ZN(new_n400_));
  AND2_X1   g199(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n401_));
  NOR2_X1   g200(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n402_));
  OAI21_X1  g201(.A(G169gat), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n400_), .B1(new_n403_), .B2(KEYINPUT79), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n405_), .B(G169gat), .C1(new_n401_), .C2(new_n402_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n397_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(G183gat), .ZN(new_n408_));
  INV_X1    g207(.A(G190gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT76), .B(KEYINPUT23), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G183gat), .A2(G190gat), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(KEYINPUT77), .A2(G183gat), .A3(G190gat), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT77), .B1(G183gat), .B2(G190gat), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT23), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n410_), .B1(new_n413_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n407_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT26), .B(G190gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT75), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT25), .B1(new_n421_), .B2(new_n408_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  OR3_X1    g222(.A1(new_n421_), .A2(new_n408_), .A3(KEYINPUT25), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G169gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n398_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(KEYINPUT24), .A3(new_n396_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(KEYINPUT24), .B2(new_n427_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n411_), .A2(new_n412_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n416_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n425_), .A2(new_n430_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n419_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G15gat), .B(G43gat), .Z(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT31), .ZN(new_n440_));
  XOR2_X1   g239(.A(KEYINPUT81), .B(KEYINPUT82), .Z(new_n441_));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G71gat), .B(G99gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n443_), .B(new_n444_), .Z(new_n445_));
  XOR2_X1   g244(.A(new_n445_), .B(new_n354_), .Z(new_n446_));
  NAND2_X1  g245(.A1(new_n440_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT31), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n439_), .B(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n446_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n395_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G8gat), .B(G36gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT18), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G64gat), .B(G92gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n454_), .B(new_n455_), .Z(new_n456_));
  INV_X1    g255(.A(KEYINPUT95), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n429_), .B1(new_n424_), .B2(new_n423_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n433_), .A2(new_n458_), .B1(new_n407_), .B2(new_n418_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G197gat), .B(G204gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT21), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G218gat), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n463_), .A2(G211gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(G211gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT89), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G211gat), .B(G218gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT89), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n462_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT90), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT90), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n462_), .A2(new_n466_), .A3(new_n469_), .A4(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n466_), .A2(new_n469_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n460_), .B(KEYINPUT21), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n471_), .A2(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n457_), .B1(new_n459_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n471_), .A2(new_n473_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n474_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(new_n435_), .A3(KEYINPUT95), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G226gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT19), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT20), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT25), .B(G183gat), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n429_), .B1(new_n420_), .B2(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n413_), .A2(new_n417_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n433_), .A2(new_n410_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT22), .B(G169gat), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n397_), .B1(new_n491_), .B2(new_n398_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n488_), .A2(new_n489_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n486_), .B1(new_n476_), .B2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n482_), .A2(new_n485_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT94), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n488_), .A2(new_n489_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n490_), .A2(new_n492_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n486_), .B1(new_n480_), .B2(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n478_), .A2(new_n419_), .A3(new_n479_), .A4(new_n434_), .ZN(new_n501_));
  AOI211_X1 g300(.A(new_n496_), .B(new_n485_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n501_), .B(KEYINPUT20), .C1(new_n476_), .C2(new_n493_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT94), .B1(new_n503_), .B2(new_n484_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n456_), .B(new_n495_), .C1(new_n502_), .C2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT96), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT20), .B1(new_n476_), .B2(new_n493_), .ZN(new_n508_));
  AND4_X1   g307(.A1(new_n478_), .A2(new_n419_), .A3(new_n479_), .A4(new_n434_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n484_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n496_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n503_), .A2(KEYINPUT94), .A3(new_n484_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n513_), .A2(KEYINPUT96), .A3(new_n456_), .A4(new_n495_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n495_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n456_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n507_), .A2(new_n514_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT27), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n485_), .B1(new_n482_), .B2(new_n494_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n503_), .A2(new_n484_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n516_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n505_), .A2(KEYINPUT27), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT28), .B1(new_n384_), .B2(KEYINPUT29), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT28), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT29), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n374_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G22gat), .B(G50gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT93), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n526_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n534_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT86), .B(G228gat), .Z(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT87), .B(G233gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n384_), .A2(KEYINPUT29), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n480_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n541_), .A2(new_n542_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n539_), .B(new_n540_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G78gat), .B(G106gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT92), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n541_), .A2(KEYINPUT85), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n539_), .A2(new_n540_), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT88), .Z(new_n552_));
  NAND2_X1  g351(.A1(new_n541_), .A2(KEYINPUT85), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n550_), .A2(new_n480_), .A3(new_n552_), .A4(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n546_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n549_), .B1(new_n546_), .B2(new_n554_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n538_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n546_), .A2(new_n554_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n548_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n546_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n537_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  AND4_X1   g361(.A1(KEYINPUT99), .A2(new_n520_), .A3(new_n525_), .A4(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n524_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT99), .B1(new_n564_), .B2(new_n562_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n452_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n393_), .A2(new_n394_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n557_), .A2(new_n561_), .A3(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n524_), .A2(new_n568_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n520_), .A2(new_n569_), .A3(KEYINPUT98), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT98), .B1(new_n520_), .B2(new_n569_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n562_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n378_), .A2(new_n379_), .A3(new_n385_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n390_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n376_), .A2(new_n380_), .A3(new_n377_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n392_), .A2(KEYINPUT33), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT33), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n386_), .A2(new_n578_), .A3(new_n390_), .A4(new_n391_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n576_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n507_), .A2(new_n517_), .A3(new_n514_), .A4(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n456_), .A2(KEYINPUT32), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n395_), .B(new_n584_), .C1(new_n515_), .C2(new_n583_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n572_), .B1(new_n581_), .B2(new_n585_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n570_), .A2(new_n571_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n447_), .A2(new_n451_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n566_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n281_), .A2(new_n318_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n322_), .A2(new_n281_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n281_), .B(new_n318_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n592_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n593_), .A2(new_n594_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G113gat), .B(G141gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(G169gat), .B(G197gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n597_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT74), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n597_), .A2(new_n600_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  NOR3_X1   g403(.A1(new_n343_), .A2(new_n590_), .A3(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(new_n276_), .A3(new_n395_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT38), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n273_), .A2(new_n274_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n604_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n330_), .A2(new_n336_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n589_), .A2(new_n611_), .A3(new_n294_), .A4(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n613_), .B2(new_n567_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n606_), .A2(new_n607_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n608_), .A2(new_n614_), .A3(new_n615_), .ZN(G1324gat));
  INV_X1    g415(.A(new_n564_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n605_), .A2(new_n277_), .A3(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n613_), .A2(new_n564_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n277_), .B1(new_n619_), .B2(KEYINPUT100), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(new_n613_), .B2(new_n564_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n620_), .A2(new_n621_), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n621_), .B1(new_n620_), .B2(new_n623_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n618_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(KEYINPUT40), .B(new_n618_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1325gat));
  INV_X1    g429(.A(G15gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n605_), .A2(new_n631_), .A3(new_n588_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT101), .Z(new_n633_));
  INV_X1    g432(.A(new_n588_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G15gat), .B1(new_n613_), .B2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT41), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n635_), .A2(KEYINPUT41), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n633_), .A2(new_n636_), .A3(new_n637_), .ZN(G1326gat));
  OAI21_X1  g437(.A(G22gat), .B1(new_n613_), .B2(new_n562_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT42), .ZN(new_n640_));
  INV_X1    g439(.A(G22gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n605_), .A2(new_n641_), .A3(new_n572_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(G1327gat));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n339_), .A2(new_n336_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT37), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n330_), .A2(new_n331_), .A3(new_n336_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT102), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n520_), .A2(new_n569_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n586_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n520_), .A2(new_n569_), .A3(KEYINPUT98), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n588_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n588_), .A2(new_n567_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n520_), .A2(new_n525_), .A3(new_n562_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n564_), .A2(KEYINPUT99), .A3(new_n562_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n649_), .B1(new_n654_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n648_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI22_X1  g464(.A1(new_n661_), .A2(KEYINPUT43), .B1(new_n589_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n611_), .A2(new_n293_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n644_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n667_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n663_), .B1(new_n589_), .B2(new_n649_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n654_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n664_), .B1(new_n671_), .B2(new_n566_), .ZN(new_n672_));
  OAI211_X1 g471(.A(KEYINPUT44), .B(new_n669_), .C1(new_n670_), .C2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n668_), .A2(new_n395_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(G29gat), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n610_), .A2(new_n294_), .A3(new_n612_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n604_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(new_n589_), .A3(new_n677_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n567_), .A2(G29gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(G1328gat));
  NOR3_X1   g479(.A1(new_n678_), .A2(G36gat), .A3(new_n564_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT45), .Z(new_n682_));
  NAND3_X1  g481(.A1(new_n668_), .A2(new_n617_), .A3(new_n673_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT103), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n668_), .A2(new_n685_), .A3(new_n673_), .A4(new_n617_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G36gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n682_), .B1(new_n684_), .B2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT104), .B(KEYINPUT46), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n682_), .B(new_n689_), .C1(new_n684_), .C2(new_n687_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1329gat));
  INV_X1    g492(.A(G43gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n634_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n668_), .A2(new_n673_), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n668_), .A2(KEYINPUT105), .A3(new_n673_), .A4(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n694_), .B1(new_n678_), .B2(new_n634_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT106), .Z(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT47), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n700_), .A2(new_n705_), .A3(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1330gat));
  OR3_X1    g506(.A1(new_n678_), .A2(G50gat), .A3(new_n562_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n668_), .A2(new_n572_), .A3(new_n673_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n709_), .A2(KEYINPUT107), .A3(G50gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT107), .B1(new_n709_), .B2(G50gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n708_), .B1(new_n710_), .B2(new_n711_), .ZN(G1331gat));
  AOI21_X1  g511(.A(new_n293_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n610_), .A2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT108), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n590_), .A2(new_n677_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT109), .Z(new_n718_));
  INV_X1    g517(.A(G57gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n395_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n609_), .A2(new_n677_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n589_), .A2(new_n294_), .A3(new_n612_), .A4(new_n721_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT110), .Z(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(new_n395_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n719_), .B2(new_n724_), .ZN(G1332gat));
  INV_X1    g524(.A(G64gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n718_), .A2(new_n726_), .A3(new_n617_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n723_), .A2(new_n617_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G64gat), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT48), .B(new_n726_), .C1(new_n723_), .C2(new_n617_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1333gat));
  INV_X1    g531(.A(G71gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n718_), .A2(new_n733_), .A3(new_n588_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT49), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n723_), .A2(new_n588_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G71gat), .ZN(new_n737_));
  AOI211_X1 g536(.A(KEYINPUT49), .B(new_n733_), .C1(new_n723_), .C2(new_n588_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1334gat));
  INV_X1    g538(.A(G78gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n718_), .A2(new_n740_), .A3(new_n572_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n723_), .A2(new_n572_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(G78gat), .ZN(new_n744_));
  AOI211_X1 g543(.A(KEYINPUT50), .B(new_n740_), .C1(new_n723_), .C2(new_n572_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1335gat));
  INV_X1    g545(.A(new_n612_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n716_), .A2(new_n610_), .A3(new_n293_), .A4(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(new_n236_), .A3(new_n395_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n721_), .A2(new_n293_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n666_), .A2(new_n567_), .A3(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n752_), .B2(new_n236_), .ZN(G1336gat));
  NAND3_X1  g552(.A1(new_n749_), .A2(new_n237_), .A3(new_n617_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n666_), .A2(new_n564_), .A3(new_n751_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(new_n237_), .ZN(G1337gat));
  NAND3_X1  g555(.A1(new_n749_), .A2(new_n588_), .A3(new_n233_), .ZN(new_n757_));
  OR3_X1    g556(.A1(new_n666_), .A2(new_n634_), .A3(new_n751_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n758_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT111), .B1(new_n758_), .B2(G99gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT51), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n763_), .B(new_n757_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1338gat));
  NAND3_X1  g564(.A1(new_n749_), .A2(new_n210_), .A3(new_n572_), .ZN(new_n766_));
  OR3_X1    g565(.A1(new_n666_), .A2(new_n562_), .A3(new_n751_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n767_), .A2(G106gat), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n767_), .B2(G106gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT53), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(new_n766_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1339gat));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n342_), .A2(new_n776_), .A3(new_n777_), .A4(new_n604_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n270_), .A2(new_n271_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n265_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT13), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n272_), .A2(KEYINPUT13), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n783_), .A2(new_n713_), .A3(new_n604_), .A4(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT114), .B1(new_n785_), .B2(KEYINPUT113), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n778_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT54), .B1(new_n785_), .B2(KEYINPUT113), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n778_), .A2(new_n786_), .A3(new_n788_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n600_), .B1(new_n595_), .B2(new_n592_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n594_), .A2(new_n591_), .A3(new_n596_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n601_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n796_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n264_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n249_), .A2(KEYINPUT12), .A3(new_n250_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n253_), .B1(new_n801_), .B2(new_n262_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT55), .B1(new_n802_), .B2(KEYINPUT115), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n801_), .A2(new_n253_), .A3(new_n262_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n801_), .A2(KEYINPUT116), .A3(new_n253_), .A4(new_n262_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n800_), .A2(new_n803_), .A3(new_n806_), .A4(new_n807_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n808_), .A2(KEYINPUT56), .A3(new_n205_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT56), .B1(new_n808_), .B2(new_n205_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n797_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n648_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT58), .B(new_n797_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n814_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n604_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n796_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT118), .B1(new_n781_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n272_), .A2(new_n825_), .A3(new_n796_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n819_), .B(KEYINPUT117), .C1(new_n809_), .C2(new_n810_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n822_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n612_), .ZN(new_n830_));
  XOR2_X1   g629(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(KEYINPUT57), .A3(new_n612_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n818_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n792_), .B1(new_n834_), .B2(new_n293_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n658_), .A2(new_n659_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n836_), .A2(new_n395_), .A3(new_n588_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT59), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n792_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n829_), .A2(KEYINPUT57), .A3(new_n612_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n831_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n829_), .B2(new_n612_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n813_), .A2(new_n815_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n840_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n839_), .B1(new_n844_), .B2(new_n294_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n837_), .A2(KEYINPUT59), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n838_), .A2(new_n847_), .A3(new_n677_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G113gat), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n835_), .A2(new_n837_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n604_), .A2(G113gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n849_), .B1(new_n851_), .B2(new_n852_), .ZN(G1340gat));
  NAND3_X1  g652(.A1(new_n838_), .A2(new_n847_), .A3(new_n610_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G120gat), .ZN(new_n855_));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n609_), .B2(KEYINPUT60), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(KEYINPUT60), .B2(new_n856_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n855_), .B1(new_n851_), .B2(new_n858_), .ZN(G1341gat));
  AOI21_X1  g658(.A(G127gat), .B1(new_n850_), .B2(new_n294_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n838_), .A2(new_n847_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n294_), .A2(G127gat), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(KEYINPUT121), .Z(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n861_), .B2(new_n863_), .ZN(G1342gat));
  NAND3_X1  g663(.A1(new_n838_), .A2(new_n847_), .A3(new_n662_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G134gat), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n612_), .A2(G134gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n851_), .B2(new_n867_), .ZN(G1343gat));
  NOR4_X1   g667(.A1(new_n617_), .A2(new_n588_), .A3(new_n562_), .A4(new_n567_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n781_), .A2(KEYINPUT118), .A3(new_n823_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n825_), .B1(new_n272_), .B2(new_n796_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n821_), .B2(new_n820_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n747_), .B1(new_n874_), .B2(new_n828_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n833_), .B1(new_n875_), .B2(new_n841_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n816_), .A2(new_n817_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n293_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n870_), .B1(new_n878_), .B2(new_n839_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n677_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n879_), .B2(new_n610_), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n835_), .A2(KEYINPUT123), .A3(new_n609_), .A4(new_n870_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT122), .B(G148gat), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n883_), .A2(new_n884_), .A3(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n840_), .A2(new_n842_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n294_), .B1(new_n888_), .B2(new_n818_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n610_), .B(new_n869_), .C1(new_n889_), .C2(new_n792_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT123), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n879_), .A2(new_n882_), .A3(new_n610_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n885_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n887_), .A2(new_n893_), .ZN(G1345gat));
  NAND2_X1  g693(.A1(new_n879_), .A2(new_n294_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1346gat));
  AND3_X1   g696(.A1(new_n879_), .A2(G162gat), .A3(new_n649_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n835_), .A2(new_n612_), .A3(new_n870_), .ZN(new_n899_));
  OR3_X1    g698(.A1(new_n899_), .A2(KEYINPUT124), .A3(G162gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT124), .B1(new_n899_), .B2(G162gat), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n898_), .B1(new_n900_), .B2(new_n901_), .ZN(G1347gat));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n655_), .A2(new_n564_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n572_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n845_), .A2(new_n677_), .A3(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n903_), .B1(new_n908_), .B2(new_n426_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n907_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n491_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .ZN(G1348gat));
  INV_X1    g711(.A(new_n844_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n792_), .B1(new_n913_), .B2(new_n293_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n906_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G176gat), .B1(new_n916_), .B2(new_n610_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n878_), .A2(new_n839_), .ZN(new_n918_));
  AOI21_X1  g717(.A(KEYINPUT125), .B1(new_n918_), .B2(new_n562_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n835_), .A2(new_n920_), .A3(new_n572_), .ZN(new_n921_));
  OR2_X1    g720(.A1(new_n919_), .A2(new_n921_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n905_), .A2(new_n609_), .A3(new_n398_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n917_), .B1(new_n922_), .B2(new_n923_), .ZN(G1349gat));
  NOR2_X1   g723(.A1(new_n293_), .A2(new_n487_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n845_), .A2(new_n906_), .A3(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT126), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n845_), .A2(new_n928_), .A3(new_n906_), .A4(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n294_), .B(new_n904_), .C1(new_n919_), .C2(new_n921_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(new_n408_), .ZN(G1350gat));
  NAND3_X1  g731(.A1(new_n916_), .A2(new_n420_), .A3(new_n747_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n914_), .A2(new_n648_), .A3(new_n915_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n934_), .B2(new_n409_), .ZN(G1351gat));
  NOR3_X1   g734(.A1(new_n588_), .A2(new_n564_), .A3(new_n568_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n918_), .A2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n937_), .A2(new_n604_), .ZN(new_n938_));
  XOR2_X1   g737(.A(KEYINPUT127), .B(G197gat), .Z(new_n939_));
  XNOR2_X1  g738(.A(new_n938_), .B(new_n939_), .ZN(G1352gat));
  NOR2_X1   g739(.A1(new_n937_), .A2(new_n609_), .ZN(new_n941_));
  INV_X1    g740(.A(G204gat), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n941_), .B(new_n942_), .ZN(G1353gat));
  NOR2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  AND2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  NOR4_X1   g744(.A1(new_n937_), .A2(new_n293_), .A3(new_n944_), .A4(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n937_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n294_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n946_), .B1(new_n948_), .B2(new_n944_), .ZN(G1354gat));
  OAI21_X1  g748(.A(G218gat), .B1(new_n937_), .B2(new_n648_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n747_), .A2(new_n463_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n937_), .B2(new_n951_), .ZN(G1355gat));
endmodule


