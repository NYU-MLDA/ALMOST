//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n203_), .B(KEYINPUT64), .Z(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT65), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT10), .B(G99gat), .Z(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT6), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G85gat), .B(G92gat), .Z(new_n217_));
  OAI21_X1  g016(.A(new_n216_), .B1(new_n217_), .B2(new_n213_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT66), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n220_), .B(new_n216_), .C1(new_n217_), .C2(new_n213_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n212_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G57gat), .B(G64gat), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n223_), .A2(KEYINPUT11), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(KEYINPUT11), .ZN(new_n225_));
  XOR2_X1   g024(.A(G71gat), .B(G78gat), .Z(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n225_), .A2(new_n226_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  OR3_X1    g029(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n211_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n217_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n232_), .B2(new_n217_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n222_), .B(new_n229_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n232_), .A2(new_n217_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT8), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n234_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n229_), .B1(new_n241_), .B2(new_n222_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n206_), .B1(new_n238_), .B2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G120gat), .B(G148gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G176gat), .B(G204gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT12), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n241_), .A2(new_n222_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(KEYINPUT68), .B(new_n250_), .C1(new_n252_), .C2(new_n229_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n242_), .B2(KEYINPUT12), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n237_), .A2(new_n205_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT69), .ZN(new_n258_));
  INV_X1    g057(.A(new_n229_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n251_), .A2(KEYINPUT12), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT67), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n242_), .A2(new_n262_), .A3(KEYINPUT12), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  AND4_X1   g063(.A1(KEYINPUT70), .A2(new_n256_), .A3(new_n258_), .A4(new_n264_), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n253_), .A2(new_n255_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT70), .B1(new_n266_), .B2(new_n258_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n243_), .B(new_n249_), .C1(new_n265_), .C2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n243_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n256_), .A2(new_n258_), .A3(new_n264_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n266_), .A2(KEYINPUT70), .A3(new_n258_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n271_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n276_), .A2(new_n249_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n270_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT13), .ZN(new_n279_));
  NOR3_X1   g078(.A1(new_n276_), .A2(new_n269_), .A3(new_n249_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n243_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(new_n248_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(new_n269_), .A3(new_n268_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT13), .B1(new_n282_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n202_), .B1(new_n281_), .B2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n279_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n282_), .A2(new_n285_), .A3(KEYINPUT13), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(KEYINPUT73), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT74), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G15gat), .B(G22gat), .ZN(new_n293_));
  INV_X1    g092(.A(G1gat), .ZN(new_n294_));
  INV_X1    g093(.A(G8gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT14), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G231gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(new_n259_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT79), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT16), .B(G183gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(G211gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(G127gat), .B(G155gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT17), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n303_), .B(new_n309_), .Z(new_n310_));
  INV_X1    g109(.A(new_n302_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(new_n308_), .A3(new_n307_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT80), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G29gat), .B(G36gat), .ZN(new_n315_));
  INV_X1    g114(.A(G43gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G50gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT15), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n251_), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n321_), .B(KEYINPUT76), .Z(new_n322_));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G232gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT34), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT75), .B(KEYINPUT35), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT77), .ZN(new_n328_));
  AOI211_X1 g127(.A(new_n323_), .B(new_n328_), .C1(new_n252_), .C2(new_n319_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n322_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n325_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n326_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G190gat), .B(G218gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G134gat), .ZN(new_n336_));
  INV_X1    g135(.A(G162gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT36), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n322_), .B(new_n329_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n334_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n334_), .A2(new_n342_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n338_), .B(KEYINPUT36), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(KEYINPUT37), .B(new_n343_), .C1(new_n344_), .C2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT37), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n334_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n346_), .B1(new_n334_), .B2(new_n342_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n292_), .A2(new_n314_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(G169gat), .ZN(new_n354_));
  INV_X1    g153(.A(G176gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(KEYINPUT24), .A3(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT25), .B(G183gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT26), .B(G190gat), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n359_), .A2(new_n360_), .A3(KEYINPUT83), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT83), .B1(new_n359_), .B2(new_n360_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n358_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT84), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n356_), .A2(KEYINPUT24), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT23), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n367_), .A2(KEYINPUT23), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n366_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(KEYINPUT84), .B(new_n358_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n365_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G204gat), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n373_), .A2(G197gat), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(G197gat), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT21), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G197gat), .B(G204gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT21), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G211gat), .B(G218gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT95), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n376_), .A2(new_n380_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT95), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n376_), .A2(new_n379_), .A3(new_n384_), .A4(new_n380_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(G169gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n354_), .A2(KEYINPUT85), .A3(KEYINPUT22), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(new_n355_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT86), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n369_), .A2(new_n368_), .ZN(new_n393_));
  INV_X1    g192(.A(G183gat), .ZN(new_n394_));
  INV_X1    g193(.A(G190gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n393_), .A2(new_n396_), .B1(G169gat), .B2(G176gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n392_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n372_), .A2(new_n387_), .A3(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT22), .B(G169gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n355_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n359_), .A2(new_n360_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n370_), .A2(new_n403_), .A3(new_n358_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n386_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT99), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT99), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n386_), .A3(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n399_), .A2(new_n407_), .A3(KEYINPUT20), .A4(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G226gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT19), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT18), .B(G64gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(G92gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G8gat), .B(G36gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT20), .B1(new_n405_), .B2(new_n386_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n372_), .A2(new_n398_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n419_), .B2(new_n386_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n412_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n413_), .A2(new_n417_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n417_), .B1(new_n413_), .B2(new_n422_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT100), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n413_), .A2(new_n422_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n417_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT100), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n413_), .A2(new_n417_), .A3(new_n422_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n425_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT0), .B(G57gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(G85gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(G1gat), .B(G29gat), .Z(new_n435_));
  XOR2_X1   g234(.A(new_n434_), .B(new_n435_), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G155gat), .A2(G162gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT90), .B1(new_n439_), .B2(KEYINPUT1), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT90), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT1), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(G155gat), .A4(G162gat), .ZN(new_n443_));
  OR2_X1    g242(.A1(G155gat), .A2(G162gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(KEYINPUT1), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n440_), .A2(new_n443_), .A3(new_n444_), .A4(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(G141gat), .ZN(new_n447_));
  INV_X1    g246(.A(G148gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G141gat), .A2(G148gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n452_));
  NOR2_X1   g251(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n449_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  AND3_X1   g253(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n454_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n444_), .A2(new_n439_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n460_), .A2(KEYINPUT92), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT92), .B1(new_n460_), .B2(new_n461_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n451_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G127gat), .A2(G134gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(G127gat), .A2(G134gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(G113gat), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G127gat), .ZN(new_n469_));
  INV_X1    g268(.A(G134gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G113gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n465_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n468_), .A2(new_n473_), .A3(G120gat), .ZN(new_n474_));
  AOI21_X1  g273(.A(G120gat), .B1(new_n468_), .B2(new_n473_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n464_), .A2(new_n477_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n451_), .B(new_n476_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(KEYINPUT4), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n460_), .A2(new_n461_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT92), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n460_), .A2(KEYINPUT92), .A3(new_n461_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n476_), .B1(new_n485_), .B2(new_n451_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT4), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n438_), .B1(new_n480_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n438_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n437_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT33), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n494_), .B(new_n437_), .C1(new_n489_), .C2(new_n491_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT101), .ZN(new_n497_));
  INV_X1    g296(.A(new_n479_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n497_), .B1(new_n486_), .B2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n478_), .A2(KEYINPUT101), .A3(new_n479_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n490_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n436_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT102), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n480_), .A2(new_n488_), .A3(new_n438_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(KEYINPUT102), .A3(new_n436_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n496_), .A2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT103), .B1(new_n432_), .B2(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n501_), .A2(KEYINPUT102), .A3(new_n436_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT102), .B1(new_n501_), .B2(new_n436_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n512_), .A2(new_n505_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT103), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n425_), .A4(new_n431_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n407_), .A2(new_n409_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n516_), .A2(KEYINPUT20), .A3(new_n421_), .A4(new_n399_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n421_), .B2(new_n420_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n417_), .A2(KEYINPUT32), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  OR3_X1    g319(.A1(new_n489_), .A2(new_n437_), .A3(new_n491_), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n518_), .A2(new_n520_), .B1(new_n521_), .B2(new_n492_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(new_n426_), .B2(new_n520_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n509_), .A2(new_n515_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n451_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT29), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n386_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT96), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n386_), .A2(new_n529_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n528_), .A2(G228gat), .A3(G233gat), .A4(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n387_), .B1(KEYINPUT29), .B2(new_n464_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(G228gat), .A3(G233gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G78gat), .B(G106gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n536_), .B(KEYINPUT97), .Z(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT94), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n539_));
  OAI21_X1  g338(.A(new_n539_), .B1(new_n464_), .B2(KEYINPUT29), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n526_), .A2(new_n527_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G22gat), .B(G50gat), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n540_), .A2(new_n542_), .A3(new_n544_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n537_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n531_), .A2(new_n534_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n538_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(KEYINPUT98), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI211_X1 g353(.A(KEYINPUT94), .B(new_n554_), .C1(new_n535_), .C2(new_n537_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n546_), .A2(new_n547_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n552_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n535_), .A2(new_n537_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n558_), .B1(new_n556_), .B2(KEYINPUT98), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n524_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT27), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n518_), .B2(new_n427_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n430_), .A2(KEYINPUT105), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n430_), .A2(KEYINPUT105), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n562_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT106), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT106), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n569_), .B(new_n562_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n521_), .A2(KEYINPUT104), .A3(new_n492_), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT104), .B1(new_n521_), .B2(new_n492_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n557_), .B(new_n559_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n561_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n419_), .A2(KEYINPUT87), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G15gat), .B(G43gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G227gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT87), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n372_), .A2(new_n583_), .A3(new_n398_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n578_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n582_), .B1(new_n578_), .B2(new_n584_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G71gat), .B(G99gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT30), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  OR3_X1    g388(.A1(new_n585_), .A2(new_n586_), .A3(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n589_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT88), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT89), .B1(new_n592_), .B2(KEYINPUT88), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n476_), .B(KEYINPUT31), .Z(new_n595_));
  INV_X1    g394(.A(KEYINPUT88), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT89), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n590_), .A2(new_n596_), .A3(new_n597_), .A4(new_n591_), .ZN(new_n598_));
  AND4_X1   g397(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .A4(new_n598_), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n594_), .A2(new_n598_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n577_), .A2(KEYINPUT107), .A3(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n572_), .A2(new_n573_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT108), .ZN(new_n606_));
  INV_X1    g405(.A(new_n571_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n607_), .B2(new_n560_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n560_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n571_), .A2(new_n609_), .A3(KEYINPUT108), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n601_), .B(new_n605_), .C1(new_n608_), .C2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT107), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n575_), .B1(new_n524_), .B2(new_n560_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n612_), .B1(new_n613_), .B2(new_n601_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n603_), .A2(new_n611_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n319_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n616_), .A2(new_n299_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n320_), .B2(new_n299_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G229gat), .A2(G233gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n319_), .B(new_n299_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(new_n619_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G113gat), .B(G141gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(G197gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT81), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(new_n354_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n620_), .A2(new_n622_), .A3(new_n627_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT82), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n615_), .A2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n353_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n294_), .A3(new_n604_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT38), .ZN(new_n637_));
  INV_X1    g436(.A(new_n631_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT109), .B1(new_n291_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT109), .ZN(new_n640_));
  AOI211_X1 g439(.A(new_n640_), .B(new_n631_), .C1(new_n287_), .C2(new_n290_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n349_), .A2(new_n350_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n615_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n642_), .A2(new_n313_), .A3(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G1gat), .B1(new_n646_), .B2(new_n605_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n637_), .A2(new_n647_), .ZN(G1324gat));
  OAI21_X1  g447(.A(G8gat), .B1(new_n646_), .B2(new_n607_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT39), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n635_), .A2(new_n295_), .A3(new_n571_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n650_), .A2(KEYINPUT40), .A3(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1325gat));
  OAI21_X1  g455(.A(G15gat), .B1(new_n646_), .B2(new_n602_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT41), .Z(new_n658_));
  INV_X1    g457(.A(G15gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n635_), .A2(new_n659_), .A3(new_n601_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(G1326gat));
  OAI21_X1  g460(.A(G22gat), .B1(new_n646_), .B2(new_n560_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT42), .ZN(new_n663_));
  INV_X1    g462(.A(G22gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n635_), .A2(new_n664_), .A3(new_n609_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(G1327gat));
  INV_X1    g465(.A(new_n314_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n644_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n634_), .A2(new_n291_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n604_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n615_), .A2(new_n672_), .A3(new_n352_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n615_), .B2(new_n352_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n642_), .B(new_n314_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(G29gat), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n615_), .A2(new_n352_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT43), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n615_), .A2(new_n672_), .A3(new_n352_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n682_), .A2(KEYINPUT44), .A3(new_n642_), .A4(new_n314_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(new_n604_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n671_), .B1(new_n678_), .B2(new_n684_), .ZN(G1328gat));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n634_), .A2(new_n291_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n607_), .A2(G36gat), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n687_), .A2(KEYINPUT45), .A3(new_n668_), .A4(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT45), .ZN(new_n690_));
  INV_X1    g489(.A(new_n688_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n669_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n677_), .A2(new_n683_), .A3(new_n571_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(G36gat), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT110), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n686_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n607_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n683_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT110), .B(KEYINPUT46), .C1(new_n700_), .C2(new_n693_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n697_), .A2(new_n701_), .ZN(G1329gat));
  OAI21_X1  g501(.A(new_n316_), .B1(new_n669_), .B2(new_n602_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n677_), .A2(G43gat), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n683_), .A2(new_n601_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n703_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g506(.A1(new_n677_), .A2(new_n683_), .A3(new_n609_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G50gat), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n609_), .A2(new_n318_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT111), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n709_), .B1(new_n669_), .B2(new_n711_), .ZN(G1331gat));
  NAND4_X1  g511(.A1(new_n292_), .A2(new_n645_), .A3(new_n632_), .A4(new_n667_), .ZN(new_n713_));
  INV_X1    g512(.A(G57gat), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n605_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n615_), .A2(new_n631_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n291_), .A2(new_n314_), .A3(new_n352_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n719_), .A2(KEYINPUT112), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(KEYINPUT112), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n604_), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n715_), .B1(new_n722_), .B2(new_n714_), .ZN(G1332gat));
  OAI21_X1  g522(.A(G64gat), .B1(new_n713_), .B2(new_n607_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT48), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n607_), .A2(G64gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n718_), .B2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n713_), .B2(new_n602_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  OR3_X1    g528(.A1(new_n718_), .A2(G71gat), .A3(new_n602_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n729_), .A2(KEYINPUT113), .A3(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1334gat));
  OR3_X1    g534(.A1(new_n718_), .A2(G78gat), .A3(new_n560_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G78gat), .B1(new_n713_), .B2(new_n560_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(KEYINPUT50), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(KEYINPUT50), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n736_), .B1(new_n740_), .B2(new_n741_), .ZN(G1335gat));
  AND2_X1   g541(.A1(new_n292_), .A2(new_n668_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n716_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G85gat), .B1(new_n745_), .B2(new_n604_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n291_), .A2(new_n638_), .A3(new_n667_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n682_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT115), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT115), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n682_), .A2(new_n750_), .A3(new_n747_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n605_), .A2(new_n214_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n746_), .B1(new_n752_), .B2(new_n753_), .ZN(G1336gat));
  NAND4_X1  g553(.A1(new_n749_), .A2(G92gat), .A3(new_n571_), .A4(new_n751_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n215_), .B1(new_n744_), .B2(new_n607_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(G1337gat));
  NAND3_X1  g558(.A1(new_n749_), .A2(new_n601_), .A3(new_n751_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G99gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n745_), .A2(new_n207_), .A3(new_n601_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT51), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n765_), .A3(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1338gat));
  OAI211_X1 g566(.A(new_n747_), .B(new_n609_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(G106gat), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(KEYINPUT117), .A3(G106gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(KEYINPUT52), .A3(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n745_), .A2(new_n208_), .A3(new_n609_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n769_), .A2(new_n770_), .A3(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n773_), .A2(new_n774_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT53), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n773_), .A2(new_n779_), .A3(new_n774_), .A4(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1339gat));
  AOI21_X1  g580(.A(new_n633_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n352_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n667_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n784_), .B(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n266_), .A2(KEYINPUT55), .A3(new_n258_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n266_), .A2(new_n237_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n206_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n265_), .A2(new_n267_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n787_), .B(new_n789_), .C1(new_n790_), .C2(KEYINPUT55), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n248_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n792_), .A2(KEYINPUT56), .B1(new_n276_), .B2(new_n249_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n619_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n627_), .B1(new_n618_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n794_), .B2(new_n621_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n796_), .A2(new_n630_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n791_), .A2(new_n798_), .A3(new_n248_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n793_), .A2(new_n797_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n793_), .A2(KEYINPUT58), .A3(new_n797_), .A4(new_n799_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n352_), .A3(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT118), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n793_), .A2(new_n638_), .A3(new_n799_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n282_), .A2(new_n285_), .A3(new_n797_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n643_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n805_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n313_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n786_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n601_), .B(new_n604_), .C1(new_n608_), .C2(new_n610_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n472_), .B1(new_n815_), .B2(new_n631_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT59), .B1(new_n813_), .B2(new_n814_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n806_), .A2(new_n807_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n809_), .B1(new_n818_), .B2(new_n643_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n808_), .A2(KEYINPUT57), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n804_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n786_), .B1(new_n821_), .B2(new_n314_), .ZN(new_n822_));
  XOR2_X1   g621(.A(new_n814_), .B(KEYINPUT119), .Z(new_n823_));
  OR3_X1    g622(.A1(new_n822_), .A2(KEYINPUT59), .A3(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n817_), .A2(G113gat), .A3(new_n633_), .A4(new_n824_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n816_), .A2(new_n825_), .ZN(G1340gat));
  INV_X1    g625(.A(G120gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n291_), .B2(KEYINPUT60), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT120), .B1(new_n827_), .B2(KEYINPUT60), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n814_), .B(new_n813_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n828_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n817_), .A2(new_n292_), .A3(new_n824_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G120gat), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(G1341gat));
  OAI21_X1  g634(.A(new_n469_), .B1(new_n815_), .B2(new_n314_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n817_), .A2(G127gat), .A3(new_n313_), .A4(new_n824_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1342gat));
  OAI21_X1  g637(.A(new_n470_), .B1(new_n815_), .B2(new_n644_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n817_), .A2(G134gat), .A3(new_n352_), .A4(new_n824_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1343gat));
  NOR4_X1   g640(.A1(new_n601_), .A2(new_n605_), .A3(new_n560_), .A4(new_n571_), .ZN(new_n842_));
  XOR2_X1   g641(.A(new_n842_), .B(KEYINPUT121), .Z(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n813_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n638_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n292_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g648(.A1(new_n845_), .A2(new_n667_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT61), .B(G155gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1346gat));
  INV_X1    g651(.A(new_n813_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n843_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n854_), .A2(new_n337_), .A3(new_n783_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n813_), .A2(new_n644_), .A3(new_n844_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT122), .B1(new_n856_), .B2(G162gat), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n858_), .B(new_n337_), .C1(new_n854_), .C2(new_n644_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n855_), .B1(new_n857_), .B2(new_n859_), .ZN(G1347gat));
  NAND2_X1  g659(.A1(new_n821_), .A2(new_n314_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n786_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n601_), .A2(new_n605_), .A3(new_n571_), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(KEYINPUT123), .Z(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n560_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n863_), .A2(new_n864_), .A3(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT125), .B1(new_n822_), .B2(new_n867_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n638_), .A3(new_n400_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n667_), .B1(new_n810_), .B2(new_n804_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n638_), .B(new_n868_), .C1(new_n873_), .C2(new_n786_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT124), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n863_), .A2(new_n876_), .A3(new_n638_), .A4(new_n868_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(G169gat), .A3(new_n877_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n878_), .A2(KEYINPUT62), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(KEYINPUT62), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n872_), .B1(new_n879_), .B2(new_n880_), .ZN(G1348gat));
  NAND3_X1  g680(.A1(new_n292_), .A2(G176gat), .A3(new_n866_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n813_), .A2(new_n609_), .A3(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n871_), .A2(new_n290_), .A3(new_n287_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n355_), .ZN(G1349gat));
  NAND4_X1  g684(.A1(new_n853_), .A2(new_n560_), .A3(new_n667_), .A4(new_n866_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n812_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n359_), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n886_), .A2(new_n394_), .B1(new_n887_), .B2(new_n888_), .ZN(G1350gat));
  NAND3_X1  g688(.A1(new_n871_), .A2(new_n643_), .A3(new_n360_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT126), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n871_), .A2(new_n352_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(G190gat), .ZN(new_n893_));
  AOI211_X1 g692(.A(KEYINPUT126), .B(new_n395_), .C1(new_n871_), .C2(new_n352_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n890_), .B1(new_n893_), .B2(new_n894_), .ZN(G1351gat));
  NAND3_X1  g694(.A1(new_n602_), .A2(new_n609_), .A3(new_n571_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n813_), .A2(new_n604_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n638_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n292_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  AND2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n897_), .B(new_n313_), .C1(new_n902_), .C2(new_n903_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n897_), .A2(new_n313_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n902_), .ZN(G1354gat));
  AOI21_X1  g705(.A(G218gat), .B1(new_n897_), .B2(new_n643_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n352_), .A2(G218gat), .ZN(new_n908_));
  XOR2_X1   g707(.A(new_n908_), .B(KEYINPUT127), .Z(new_n909_));
  AOI21_X1  g708(.A(new_n907_), .B1(new_n897_), .B2(new_n909_), .ZN(G1355gat));
endmodule


