//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT71), .ZN(new_n203_));
  INV_X1    g002(.A(G230gat), .ZN(new_n204_));
  INV_X1    g003(.A(G233gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  OAI22_X1  g010(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n213_));
  INV_X1    g012(.A(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n211_), .A2(new_n212_), .A3(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT9), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n219_), .A2(KEYINPUT64), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n229_), .A2(new_n218_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232_));
  INV_X1    g031(.A(new_n219_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n232_), .B1(new_n233_), .B2(KEYINPUT9), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT10), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n214_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n215_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n211_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n217_), .A2(new_n225_), .A3(new_n221_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n227_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G71gat), .B(G78gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G57gat), .B(G64gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT67), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n248_), .B2(KEYINPUT11), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n247_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT11), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n251_), .A2(KEYINPUT68), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n254_), .B1(new_n248_), .B2(KEYINPUT11), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n249_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT68), .B1(new_n251_), .B2(new_n252_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n245_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n248_), .A2(new_n254_), .A3(KEYINPUT11), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n244_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(KEYINPUT69), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n256_), .A2(new_n244_), .A3(new_n260_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(new_n261_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n206_), .B1(new_n263_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT12), .ZN(new_n270_));
  INV_X1    g069(.A(new_n206_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT12), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n264_), .A2(new_n268_), .A3(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n270_), .A2(new_n271_), .A3(new_n273_), .A4(new_n262_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G120gat), .B(G148gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT5), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G176gat), .B(G204gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n267_), .A2(new_n274_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n279_), .B1(new_n267_), .B2(new_n274_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n203_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n281_), .A2(new_n203_), .A3(new_n282_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n202_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n285_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(KEYINPUT13), .A3(new_n283_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n286_), .A2(new_n288_), .A3(KEYINPUT72), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G229gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G29gat), .B(G36gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G43gat), .B(G50gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n295_), .ZN(new_n298_));
  XOR2_X1   g097(.A(G43gat), .B(G50gat), .Z(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G1gat), .A2(G8gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT14), .ZN(new_n302_));
  NOR2_X1   g101(.A1(G15gat), .A2(G22gat), .ZN(new_n303_));
  AND2_X1   g102(.A1(G15gat), .A2(G22gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT78), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT79), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT78), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n302_), .B(new_n308_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G1gat), .B(G8gat), .Z(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n307_), .B1(new_n306_), .B2(new_n309_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n311_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n314_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n312_), .B1(new_n316_), .B2(new_n310_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n297_), .B(new_n300_), .C1(new_n315_), .C2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n313_), .B1(new_n311_), .B2(new_n314_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n316_), .A2(new_n312_), .A3(new_n310_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n300_), .A2(new_n297_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT82), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n318_), .A2(KEYINPUT82), .A3(new_n322_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n294_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n317_), .A2(new_n315_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT15), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n321_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n300_), .A2(KEYINPUT15), .A3(new_n297_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n294_), .A3(new_n322_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n327_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT84), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G113gat), .B(G141gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G169gat), .B(G197gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n338_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n294_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n326_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT82), .B1(new_n318_), .B2(new_n322_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n343_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(new_n335_), .A3(new_n341_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT84), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n342_), .A2(new_n348_), .ZN(new_n349_));
  OR3_X1    g148(.A1(new_n327_), .A2(new_n336_), .A3(KEYINPUT83), .ZN(new_n350_));
  INV_X1    g149(.A(new_n341_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT83), .B1(new_n327_), .B2(new_n336_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(G134gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G127gat), .ZN(new_n357_));
  INV_X1    g156(.A(G127gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(G134gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G120gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(G113gat), .ZN(new_n362_));
  INV_X1    g161(.A(G113gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(G120gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n360_), .A2(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n357_), .A2(new_n359_), .A3(new_n362_), .A4(new_n364_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT86), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT87), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n369_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n366_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n368_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT87), .ZN(new_n374_));
  INV_X1    g173(.A(new_n366_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n372_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G71gat), .B(G99gat), .ZN(new_n379_));
  INV_X1    g178(.A(G43gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT30), .ZN(new_n382_));
  NOR2_X1   g181(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G169gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G183gat), .A2(G190gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT23), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n387_), .B(new_n388_), .C1(G183gat), .C2(G190gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n384_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n388_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(G169gat), .B2(G176gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(G190gat), .ZN(new_n398_));
  OR3_X1    g197(.A1(new_n398_), .A2(KEYINPUT85), .A3(KEYINPUT26), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT25), .B(G183gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT26), .B1(new_n398_), .B2(KEYINPUT85), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n390_), .B1(new_n397_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n382_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT30), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n381_), .B(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n404_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n411_), .B(G15gat), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT88), .B1(new_n410_), .B2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n414_), .B1(new_n413_), .B2(new_n410_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n415_), .A2(KEYINPUT31), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(KEYINPUT31), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n378_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n415_), .A2(KEYINPUT31), .ZN(new_n419_));
  INV_X1    g218(.A(new_n378_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(KEYINPUT31), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n424_));
  INV_X1    g223(.A(G141gat), .ZN(new_n425_));
  INV_X1    g224(.A(G148gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT90), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n424_), .B1(new_n427_), .B2(KEYINPUT3), .ZN(new_n428_));
  NAND3_X1  g227(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT91), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT91), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n431_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT3), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n434_), .A2(new_n425_), .A3(new_n426_), .A4(KEYINPUT90), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n428_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G155gat), .A2(G162gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT89), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT89), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(G155gat), .B2(G162gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G155gat), .A2(G162gat), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n438_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n436_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(KEYINPUT1), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT1), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(G155gat), .A3(G162gat), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n438_), .A2(new_n440_), .A3(new_n444_), .A4(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G141gat), .B(G148gat), .Z(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT92), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT92), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n443_), .A2(new_n452_), .A3(new_n449_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n451_), .A2(new_n453_), .A3(new_n377_), .A4(new_n372_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G225gat), .A2(G233gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT100), .B1(new_n366_), .B2(new_n367_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n366_), .A2(KEYINPUT100), .A3(new_n367_), .ZN(new_n457_));
  OR3_X1    g256(.A1(new_n450_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(new_n455_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT101), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT101), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n454_), .A2(new_n458_), .A3(new_n461_), .A4(new_n455_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  AOI221_X4 g262(.A(KEYINPUT92), .B1(new_n447_), .B2(new_n448_), .C1(new_n436_), .C2(new_n442_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n452_), .B1(new_n443_), .B2(new_n449_), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n378_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n450_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT4), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT4), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n454_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n455_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n463_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT102), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G29gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(G85gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT0), .B(G57gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n472_), .A2(new_n473_), .A3(KEYINPUT33), .A4(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n455_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n469_), .B1(new_n454_), .B2(new_n458_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n464_), .A2(new_n465_), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT4), .B1(new_n482_), .B2(new_n420_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n480_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n484_), .A2(new_n478_), .A3(new_n460_), .A4(new_n462_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT102), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n486_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT20), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G211gat), .B(G218gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G197gat), .B(G204gat), .ZN(new_n491_));
  INV_X1    g290(.A(G204gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT95), .B1(new_n492_), .B2(G197gat), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n490_), .A2(new_n491_), .A3(KEYINPUT21), .A4(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n490_), .A2(KEYINPUT21), .A3(new_n493_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n490_), .A2(KEYINPUT21), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(new_n491_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n495_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT26), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G190gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n398_), .A2(KEYINPUT26), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n501_), .A2(new_n502_), .A3(KEYINPUT97), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT97), .B1(new_n501_), .B2(new_n502_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n400_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n395_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n505_), .A2(new_n506_), .B1(new_n389_), .B2(new_n384_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n489_), .B1(new_n499_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G226gat), .A2(G233gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT19), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n491_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(KEYINPUT21), .B2(new_n490_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n496_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n494_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT98), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n404_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n516_), .B1(new_n404_), .B2(new_n515_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n508_), .B(new_n511_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n499_), .A2(new_n507_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT20), .B1(new_n404_), .B2(new_n515_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n510_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G8gat), .B(G36gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G64gat), .B(G92gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n523_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n519_), .A2(new_n528_), .A3(new_n522_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n454_), .A2(new_n480_), .A3(new_n458_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT103), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n477_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n533_), .B2(new_n477_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n455_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n532_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n479_), .A2(new_n487_), .A3(new_n488_), .A4(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n528_), .A2(KEYINPUT32), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n541_), .B1(new_n523_), .B2(KEYINPUT104), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n508_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n510_), .ZN(new_n544_));
  OR3_X1    g343(.A1(new_n520_), .A2(new_n521_), .A3(new_n510_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(KEYINPUT32), .A3(new_n528_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n519_), .A2(KEYINPUT104), .A3(new_n522_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n542_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n477_), .B1(new_n463_), .B2(new_n471_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n485_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n540_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n451_), .A2(new_n453_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT28), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT29), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n555_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G22gat), .B(G50gat), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT93), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  OR3_X1    g361(.A1(new_n558_), .A2(new_n559_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT94), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(G228gat), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(G228gat), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n205_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n499_), .A2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n556_), .B1(new_n443_), .B2(new_n449_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n568_), .B1(new_n571_), .B2(new_n499_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G78gat), .B(G106gat), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n570_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT96), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n562_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n563_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n570_), .A2(new_n572_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n573_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n575_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n579_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n553_), .A2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n579_), .B(new_n582_), .Z(new_n585_));
  OAI211_X1 g384(.A(KEYINPUT27), .B(new_n531_), .C1(new_n546_), .C2(new_n528_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT27), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n532_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n551_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n585_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n423_), .B1(new_n584_), .B2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n423_), .A2(new_n583_), .A3(new_n590_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(new_n551_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n293_), .A2(new_n355_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT76), .ZN(new_n598_));
  XOR2_X1   g397(.A(G190gat), .B(G218gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT75), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(KEYINPUT36), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n227_), .A2(new_n242_), .A3(new_n243_), .A4(new_n321_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n217_), .A2(new_n225_), .A3(new_n221_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n240_), .B1(new_n234_), .B2(new_n231_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n225_), .B1(new_n217_), .B2(new_n221_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n605_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n331_), .A2(new_n332_), .ZN(new_n609_));
  OAI211_X1 g408(.A(KEYINPUT74), .B(new_n604_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT73), .B(KEYINPUT35), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n333_), .A2(new_n244_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT34), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(new_n604_), .A3(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n614_), .A2(KEYINPUT74), .A3(new_n604_), .A4(new_n611_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n613_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n616_), .B1(new_n613_), .B2(new_n619_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n603_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n613_), .A2(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n617_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n613_), .A2(new_n619_), .A3(new_n618_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n602_), .B(KEYINPUT36), .Z(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n598_), .B1(new_n622_), .B2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n620_), .A2(new_n621_), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT76), .B1(new_n629_), .B2(new_n626_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n628_), .A2(new_n630_), .A3(KEYINPUT37), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT37), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n622_), .B2(new_n627_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n631_), .A2(KEYINPUT77), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT77), .ZN(new_n635_));
  INV_X1    g434(.A(new_n626_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n620_), .A2(new_n636_), .A3(new_n621_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n603_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT76), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n627_), .A2(new_n598_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n632_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n633_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n635_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n634_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n256_), .A2(new_n260_), .ZN(new_n646_));
  INV_X1    g445(.A(G231gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n647_), .B2(new_n205_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n256_), .A2(G231gat), .A3(new_n260_), .A4(G233gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT80), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n650_), .A2(KEYINPUT80), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n329_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n653_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n328_), .A3(new_n651_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(G127gat), .B(G155gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT16), .ZN(new_n659_));
  XOR2_X1   g458(.A(G183gat), .B(G211gat), .Z(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT17), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT81), .B1(new_n657_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n657_), .A2(new_n662_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT17), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n661_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n664_), .B1(new_n667_), .B2(new_n657_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n663_), .B1(new_n668_), .B2(KEYINPUT81), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n645_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n597_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n673_), .A2(G1gat), .A3(new_n591_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT38), .Z(new_n675_));
  INV_X1    g474(.A(new_n669_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n628_), .A2(new_n630_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n597_), .A2(new_n551_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G1gat), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n675_), .A2(new_n680_), .ZN(G1324gat));
  OR3_X1    g480(.A1(new_n673_), .A2(G8gat), .A3(new_n590_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n597_), .A2(new_n589_), .A3(new_n678_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT39), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(new_n684_), .A3(G8gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n683_), .B2(G8gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT40), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1325gat));
  NAND3_X1  g488(.A1(new_n597_), .A2(new_n423_), .A3(new_n678_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n690_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT41), .B1(new_n690_), .B2(G15gat), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n418_), .A2(new_n422_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n693_), .A2(G15gat), .ZN(new_n694_));
  OAI22_X1  g493(.A1(new_n691_), .A2(new_n692_), .B1(new_n673_), .B2(new_n694_), .ZN(G1326gat));
  NAND3_X1  g494(.A1(new_n597_), .A2(new_n585_), .A3(new_n678_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G22gat), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(KEYINPUT42), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(KEYINPUT42), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n583_), .A2(G22gat), .ZN(new_n700_));
  OAI22_X1  g499(.A1(new_n698_), .A2(new_n699_), .B1(new_n673_), .B2(new_n700_), .ZN(G1327gat));
  OAI21_X1  g500(.A(KEYINPUT77), .B1(new_n631_), .B2(new_n633_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n642_), .A2(new_n635_), .A3(new_n643_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(KEYINPUT105), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n705_), .B1(new_n634_), .B2(new_n644_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n704_), .B(new_n706_), .C1(new_n593_), .C2(new_n595_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT43), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n585_), .B1(new_n552_), .B2(new_n540_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n583_), .A2(new_n589_), .A3(new_n551_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n693_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n594_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n591_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n645_), .A2(KEYINPUT43), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n708_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n291_), .A2(new_n676_), .A3(new_n292_), .A4(new_n354_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n717_), .A2(new_n718_), .A3(new_n719_), .A4(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n718_), .A2(new_n719_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n707_), .A2(KEYINPUT43), .B1(new_n714_), .B2(new_n715_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n723_), .B(new_n724_), .C1(new_n725_), .C2(new_n720_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n591_), .B1(new_n722_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(G29gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n676_), .A2(new_n677_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n597_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n551_), .A2(new_n728_), .ZN(new_n732_));
  OAI22_X1  g531(.A1(new_n727_), .A2(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(G1328gat));
  NOR2_X1   g532(.A1(new_n590_), .A2(G36gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n597_), .A2(new_n730_), .A3(new_n734_), .ZN(new_n735_));
  XOR2_X1   g534(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n722_), .A2(new_n726_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(new_n739_), .A3(new_n589_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G36gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n738_), .B2(new_n589_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n737_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OAI211_X1 g544(.A(KEYINPUT46), .B(new_n737_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1329gat));
  NOR2_X1   g546(.A1(new_n693_), .A2(new_n380_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n738_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n597_), .A2(new_n423_), .A3(new_n730_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT109), .B1(new_n750_), .B2(new_n380_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n738_), .A2(new_n753_), .A3(new_n748_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT47), .B1(new_n752_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n754_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n756_), .B(new_n757_), .C1(new_n749_), .C2(new_n751_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(new_n758_), .ZN(G1330gat));
  INV_X1    g558(.A(G50gat), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n583_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n597_), .A2(new_n585_), .A3(new_n730_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n738_), .A2(new_n761_), .B1(new_n760_), .B2(new_n762_), .ZN(G1331gat));
  NOR2_X1   g562(.A1(new_n596_), .A2(new_n354_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n678_), .A3(new_n293_), .ZN(new_n765_));
  INV_X1    g564(.A(G57gat), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n591_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n293_), .A2(new_n671_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT110), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n764_), .B(KEYINPUT111), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n771_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n768_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n775_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(KEYINPUT113), .A3(new_n773_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n776_), .A2(new_n778_), .A3(new_n551_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n767_), .B1(new_n779_), .B2(new_n766_), .ZN(G1332gat));
  NOR2_X1   g579(.A1(new_n774_), .A2(new_n775_), .ZN(new_n781_));
  INV_X1    g580(.A(G64gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n589_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G64gat), .B1(new_n765_), .B2(new_n590_), .ZN(new_n784_));
  XOR2_X1   g583(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n785_));
  XNOR2_X1  g584(.A(new_n784_), .B(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n783_), .A2(new_n786_), .ZN(G1333gat));
  INV_X1    g586(.A(G71gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n781_), .A2(new_n788_), .A3(new_n423_), .ZN(new_n789_));
  OAI21_X1  g588(.A(G71gat), .B1(new_n765_), .B2(new_n693_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT49), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1334gat));
  INV_X1    g591(.A(G78gat), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n781_), .A2(new_n793_), .A3(new_n585_), .ZN(new_n794_));
  OAI21_X1  g593(.A(G78gat), .B1(new_n765_), .B2(new_n583_), .ZN(new_n795_));
  XOR2_X1   g594(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n797_), .ZN(G1335gat));
  AOI211_X1 g597(.A(new_n354_), .B(new_n669_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n717_), .A2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(G85gat), .B1(new_n800_), .B2(new_n591_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n293_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(new_n729_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n772_), .A2(new_n803_), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n591_), .A2(G85gat), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n801_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n806_), .B(KEYINPUT116), .Z(G1336gat));
  INV_X1    g606(.A(new_n804_), .ZN(new_n808_));
  AOI21_X1  g607(.A(G92gat), .B1(new_n808_), .B2(new_n589_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n800_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n589_), .A2(G92gat), .ZN(new_n811_));
  XOR2_X1   g610(.A(new_n811_), .B(KEYINPUT117), .Z(new_n812_));
  AOI21_X1  g611(.A(new_n809_), .B1(new_n810_), .B2(new_n812_), .ZN(G1337gat));
  OAI21_X1  g612(.A(G99gat), .B1(new_n800_), .B2(new_n693_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n423_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n804_), .B2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g616(.A1(new_n808_), .A2(new_n215_), .A3(new_n585_), .ZN(new_n818_));
  OAI21_X1  g617(.A(G106gat), .B1(new_n800_), .B2(new_n583_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(KEYINPUT52), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(KEYINPUT52), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n818_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g622(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n294_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n334_), .A2(new_n343_), .A3(new_n322_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n826_), .A2(new_n351_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n342_), .A2(new_n348_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n270_), .A2(new_n273_), .A3(new_n262_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n206_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT55), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n274_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n274_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(new_n833_), .A3(KEYINPUT55), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n279_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n828_), .B(new_n280_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n836_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n824_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n645_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n828_), .A2(new_n280_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n830_), .A2(new_n833_), .A3(KEYINPUT55), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n833_), .B1(KEYINPUT55), .B2(new_n830_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n278_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT56), .ZN(new_n846_));
  INV_X1    g645(.A(new_n824_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n842_), .A2(new_n846_), .A3(new_n847_), .A4(new_n838_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n840_), .A2(new_n841_), .A3(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n836_), .B1(new_n835_), .B2(KEYINPUT118), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n845_), .A2(new_n851_), .A3(KEYINPUT56), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n281_), .B1(new_n349_), .B2(new_n353_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n850_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n287_), .A2(new_n828_), .A3(new_n283_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n677_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n849_), .B1(new_n856_), .B2(KEYINPUT57), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(KEYINPUT57), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n676_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n289_), .A2(new_n355_), .ZN(new_n861_));
  OR3_X1    g660(.A1(new_n861_), .A2(new_n670_), .A3(KEYINPUT54), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT54), .B1(new_n861_), .B2(new_n670_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n860_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n551_), .A3(new_n712_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n363_), .A3(new_n354_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(KEYINPUT59), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n866_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n355_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n868_), .B1(new_n872_), .B2(new_n363_), .ZN(G1340gat));
  OAI21_X1  g672(.A(new_n361_), .B1(new_n802_), .B2(KEYINPUT60), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n867_), .B(new_n874_), .C1(KEYINPUT60), .C2(new_n361_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n802_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n361_), .ZN(G1341gat));
  NAND3_X1  g676(.A1(new_n867_), .A2(new_n358_), .A3(new_n669_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n676_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n358_), .ZN(G1342gat));
  NAND3_X1  g679(.A1(new_n867_), .A2(new_n356_), .A3(new_n677_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n645_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(new_n356_), .ZN(G1343gat));
  OR2_X1    g682(.A1(new_n856_), .A2(KEYINPUT57), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(new_n858_), .A3(new_n849_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n885_), .A2(new_n676_), .B1(new_n863_), .B2(new_n862_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n591_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n423_), .A2(new_n583_), .A3(new_n589_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n355_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n425_), .ZN(G1344gat));
  NOR2_X1   g690(.A1(new_n889_), .A2(new_n802_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT120), .B(G148gat), .Z(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1345gat));
  NOR2_X1   g693(.A1(new_n889_), .A2(new_n676_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n895_), .B(new_n897_), .ZN(G1346gat));
  AND2_X1   g697(.A1(new_n887_), .A2(new_n888_), .ZN(new_n899_));
  AOI21_X1  g698(.A(G162gat), .B1(new_n899_), .B2(new_n677_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n706_), .A2(G162gat), .A3(new_n704_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT121), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n900_), .B1(new_n899_), .B2(new_n902_), .ZN(G1347gat));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n585_), .A2(new_n693_), .A3(new_n551_), .A4(new_n590_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n865_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n355_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT22), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n904_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(G169gat), .ZN(new_n910_));
  INV_X1    g709(.A(G169gat), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(new_n907_), .B2(new_n904_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n909_), .B2(new_n912_), .ZN(G1348gat));
  NOR2_X1   g712(.A1(new_n906_), .A2(new_n802_), .ZN(new_n914_));
  INV_X1    g713(.A(G176gat), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n915_), .A2(KEYINPUT122), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(KEYINPUT122), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n914_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n914_), .B2(new_n917_), .ZN(G1349gat));
  NOR2_X1   g718(.A1(new_n906_), .A2(new_n676_), .ZN(new_n920_));
  MUX2_X1   g719(.A(G183gat), .B(new_n400_), .S(new_n920_), .Z(G1350gat));
  NOR2_X1   g720(.A1(new_n503_), .A2(new_n504_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n865_), .A2(new_n923_), .A3(new_n677_), .A4(new_n905_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n906_), .A2(new_n645_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n398_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  OAI211_X1 g727(.A(KEYINPUT123), .B(new_n924_), .C1(new_n925_), .C2(new_n398_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1351gat));
  NOR3_X1   g729(.A1(new_n423_), .A2(new_n583_), .A3(new_n551_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT124), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n589_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(KEYINPUT125), .B1(new_n865_), .B2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936_));
  AOI211_X1 g735(.A(new_n936_), .B(new_n933_), .C1(new_n860_), .C2(new_n864_), .ZN(new_n937_));
  OAI211_X1 g736(.A(G197gat), .B(new_n354_), .C1(new_n935_), .C2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(KEYINPUT126), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n936_), .B1(new_n886_), .B2(new_n933_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n865_), .A2(KEYINPUT125), .A3(new_n934_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943_));
  NAND4_X1  g742(.A1(new_n942_), .A2(new_n943_), .A3(G197gat), .A4(new_n354_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n354_), .B1(new_n935_), .B2(new_n937_), .ZN(new_n945_));
  INV_X1    g744(.A(G197gat), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  AND3_X1   g746(.A1(new_n939_), .A2(new_n944_), .A3(new_n947_), .ZN(G1352gat));
  NAND2_X1  g747(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n942_), .A2(new_n293_), .A3(new_n949_), .ZN(new_n950_));
  INV_X1    g749(.A(new_n942_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n951_), .A2(new_n802_), .ZN(new_n952_));
  XOR2_X1   g751(.A(KEYINPUT127), .B(G204gat), .Z(new_n953_));
  OAI21_X1  g752(.A(new_n950_), .B1(new_n952_), .B2(new_n953_), .ZN(G1353gat));
  NOR2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  AND2_X1   g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  OAI211_X1 g755(.A(new_n942_), .B(new_n669_), .C1(new_n955_), .C2(new_n956_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n951_), .A2(new_n676_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n958_), .B2(new_n955_), .ZN(G1354gat));
  OAI21_X1  g758(.A(G218gat), .B1(new_n951_), .B2(new_n645_), .ZN(new_n960_));
  INV_X1    g759(.A(G218gat), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n942_), .A2(new_n961_), .A3(new_n677_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n960_), .A2(new_n962_), .ZN(G1355gat));
endmodule


