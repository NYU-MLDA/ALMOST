//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n601_, new_n602_, new_n603_, new_n604_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT71), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G50gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT71), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n203_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G50gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n205_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT15), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n205_), .A2(new_n209_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT15), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT10), .B(G99gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT6), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G85gat), .B(G92gat), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT9), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(G85gat), .A3(G92gat), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n220_), .A2(new_n224_), .A3(new_n226_), .A4(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT8), .ZN(new_n231_));
  INV_X1    g030(.A(G99gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n219_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT7), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT65), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT65), .B(KEYINPUT7), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n236_), .B1(new_n237_), .B2(new_n233_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n231_), .B(new_n225_), .C1(new_n238_), .C2(new_n223_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n225_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n223_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n236_), .B(KEYINPUT66), .C1(new_n237_), .C2(new_n233_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n240_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n239_), .B1(new_n244_), .B2(new_n231_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n230_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(KEYINPUT68), .B(new_n239_), .C1(new_n244_), .C2(new_n231_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT69), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT7), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n233_), .B1(new_n251_), .B2(new_n235_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n232_), .A2(new_n219_), .B1(new_n234_), .B2(KEYINPUT65), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n241_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(new_n243_), .A3(new_n224_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n231_), .B1(new_n255_), .B2(new_n225_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n239_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n246_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n258_), .A2(KEYINPUT69), .A3(new_n229_), .A4(new_n248_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n215_), .B1(new_n249_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G232gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT34), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT35), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n212_), .A2(new_n245_), .A3(new_n229_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n261_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n264_), .A2(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n261_), .A2(new_n271_), .A3(new_n266_), .A4(new_n267_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G190gat), .B(G218gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G134gat), .B(G162gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(KEYINPUT72), .B(KEYINPUT73), .Z(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n278_), .A2(KEYINPUT36), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT74), .B1(new_n273_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT74), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n270_), .A2(new_n282_), .A3(new_n279_), .A4(new_n272_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT37), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n278_), .B(KEYINPUT36), .Z(new_n286_));
  NAND2_X1  g085(.A1(new_n273_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n286_), .B(KEYINPUT75), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n281_), .A2(new_n283_), .B1(new_n273_), .B2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n285_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT17), .ZN(new_n293_));
  XOR2_X1   g092(.A(G15gat), .B(G22gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT76), .B(G8gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G1gat), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(new_n296_), .B2(KEYINPUT14), .ZN(new_n297_));
  INV_X1    g096(.A(G1gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(G8gat), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n300_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G231gat), .A2(G233gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n303_), .B(new_n304_), .Z(new_n305_));
  INV_X1    g104(.A(G64gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G57gat), .ZN(new_n307_));
  INV_X1    g106(.A(G57gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G64gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT11), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G71gat), .B(G78gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n307_), .A2(new_n309_), .A3(KEYINPUT11), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n313_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n305_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n305_), .A2(new_n317_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G183gat), .B(G211gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G127gat), .B(G155gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  OR4_X1    g123(.A1(new_n293_), .A2(new_n318_), .A3(new_n319_), .A4(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT67), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n313_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n327_));
  AND4_X1   g126(.A1(KEYINPUT11), .A2(new_n311_), .A3(new_n307_), .A4(new_n309_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n326_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n315_), .A2(KEYINPUT67), .A3(new_n316_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n305_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n305_), .A2(new_n332_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n324_), .B(KEYINPUT17), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n325_), .A2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n292_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT12), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n317_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n258_), .A2(new_n229_), .A3(new_n248_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT69), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n341_), .B1(new_n344_), .B2(new_n259_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n331_), .B(new_n229_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G230gat), .A2(G233gat), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n245_), .A2(new_n229_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT12), .B1(new_n352_), .B2(new_n332_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n345_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n332_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n348_), .B1(new_n355_), .B2(new_n346_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G120gat), .B(G148gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G204gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT5), .B(G176gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n357_), .B(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n363_), .A2(KEYINPUT13), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(KEYINPUT13), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n338_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G127gat), .B(G134gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT84), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(G113gat), .ZN(new_n372_));
  INV_X1    g171(.A(G120gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  OR2_X1    g173(.A1(G141gat), .A2(G148gat), .ZN(new_n375_));
  NAND3_X1  g174(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G141gat), .A2(G148gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G155gat), .B(G162gat), .Z(new_n379_));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n378_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT85), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n375_), .B(KEYINPUT3), .Z(new_n383_));
  XNOR2_X1  g182(.A(new_n377_), .B(KEYINPUT2), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n382_), .B1(new_n379_), .B2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n374_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n369_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT90), .B1(new_n374_), .B2(new_n386_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n374_), .A2(new_n386_), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT4), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n393_), .A2(KEYINPUT91), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(KEYINPUT91), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n389_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n396_), .A2(KEYINPUT92), .B1(new_n392_), .B2(new_n369_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n394_), .A2(new_n395_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT92), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n399_), .A3(new_n389_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(G1gat), .B(G29gat), .Z(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT94), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G57gat), .B(G85gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n403_), .B(new_n406_), .Z(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n401_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n397_), .A2(new_n400_), .A3(new_n407_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT22), .B(G169gat), .ZN(new_n413_));
  INV_X1    g212(.A(G176gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT81), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G183gat), .A2(G190gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(KEYINPUT23), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n417_), .B(KEYINPUT80), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n419_), .B1(new_n420_), .B2(KEYINPUT23), .ZN(new_n421_));
  NOR2_X1   g220(.A1(G183gat), .A2(G190gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G169gat), .A2(G176gat), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n416_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT25), .B(G183gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT26), .B(G190gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(G169gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n414_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(KEYINPUT24), .A3(new_n425_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT79), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT23), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n420_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(new_n435_), .B2(new_n418_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n431_), .A2(KEYINPUT24), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n426_), .B1(new_n434_), .B2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT82), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT30), .ZN(new_n442_));
  XOR2_X1   g241(.A(G15gat), .B(G43gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G227gat), .A2(G233gat), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n445_), .B(KEYINPUT83), .Z(new_n446_));
  XNOR2_X1  g245(.A(new_n444_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n374_), .B(KEYINPUT31), .ZN(new_n448_));
  XOR2_X1   g247(.A(G71gat), .B(G99gat), .Z(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n447_), .A2(new_n450_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G197gat), .B(G204gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(G211gat), .B(G218gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n455_), .B1(KEYINPUT21), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(KEYINPUT21), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT29), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n460_), .B1(new_n386_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G228gat), .A2(G233gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(G78gat), .B(G106gat), .Z(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT86), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n386_), .A2(new_n461_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G22gat), .B(G50gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT28), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n468_), .B(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n467_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n464_), .B(new_n465_), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n472_), .B(new_n473_), .Z(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n454_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n453_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n451_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n474_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n438_), .A2(new_n432_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n427_), .B(KEYINPUT87), .ZN(new_n483_));
  INV_X1    g282(.A(new_n428_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n421_), .B(new_n482_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n485_), .B(KEYINPUT88), .Z(new_n486_));
  NAND2_X1  g285(.A1(new_n437_), .A2(new_n423_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n487_), .A2(new_n425_), .A3(new_n415_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n481_), .B1(new_n490_), .B2(new_n460_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n491_), .B1(new_n460_), .B2(new_n441_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G226gat), .A2(G233gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT19), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n441_), .A2(new_n460_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n488_), .A2(new_n460_), .ZN(new_n496_));
  AOI211_X1 g295(.A(new_n481_), .B(new_n494_), .C1(new_n486_), .C2(new_n496_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n492_), .A2(new_n494_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n499_));
  XNOR2_X1  g298(.A(G8gat), .B(G36gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G64gat), .B(G92gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n498_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT27), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n498_), .B2(new_n504_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n492_), .A2(new_n494_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n496_), .B2(new_n485_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n495_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n509_), .B1(new_n494_), .B2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n508_), .B1(new_n513_), .B2(new_n504_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n507_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n412_), .A2(new_n480_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT33), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n410_), .A2(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n397_), .A2(new_n400_), .A3(KEYINPUT33), .A4(new_n407_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n369_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n398_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n407_), .B1(new_n392_), .B2(new_n521_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT95), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n505_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n519_), .A2(new_n520_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n519_), .A2(KEYINPUT96), .A3(new_n520_), .A4(new_n526_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n504_), .A2(KEYINPUT32), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n498_), .A2(new_n531_), .ZN(new_n532_));
  OAI22_X1  g331(.A1(new_n532_), .A2(KEYINPUT97), .B1(new_n513_), .B2(new_n531_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n533_), .B1(KEYINPUT97), .B2(new_n532_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n411_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n529_), .A2(new_n530_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n478_), .A2(new_n475_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n517_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT99), .ZN(new_n540_));
  INV_X1    g339(.A(new_n303_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n215_), .A2(KEYINPUT78), .A3(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n211_), .A2(new_n541_), .A3(new_n214_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT78), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n303_), .A2(new_n212_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n546_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n541_), .A2(new_n210_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n547_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n548_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G113gat), .B(G141gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(G169gat), .ZN(new_n557_));
  INV_X1    g356(.A(G197gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n551_), .A2(new_n555_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n549_), .B1(new_n542_), .B2(new_n545_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n555_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n539_), .A2(new_n540_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n540_), .B1(new_n539_), .B2(new_n566_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n368_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n570_), .A2(new_n298_), .A3(new_n411_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT38), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n536_), .A2(new_n538_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n517_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n284_), .A2(new_n287_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n337_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n366_), .A2(new_n566_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .A4(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(G1gat), .B1(new_n579_), .B2(new_n412_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n571_), .A2(KEYINPUT38), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n581_), .A2(KEYINPUT100), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(KEYINPUT100), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n572_), .B(new_n580_), .C1(new_n582_), .C2(new_n583_), .ZN(G1324gat));
  OAI21_X1  g383(.A(G8gat), .B1(new_n579_), .B2(new_n516_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT39), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT39), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n587_), .B(G8gat), .C1(new_n579_), .C2(new_n516_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n295_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n570_), .A2(new_n590_), .A3(new_n515_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT101), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT101), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n589_), .A2(new_n594_), .A3(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT40), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n593_), .A2(KEYINPUT40), .A3(new_n595_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(G1325gat));
  OAI21_X1  g399(.A(G15gat), .B1(new_n579_), .B2(new_n478_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT41), .Z(new_n602_));
  INV_X1    g401(.A(G15gat), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n570_), .A2(new_n603_), .A3(new_n454_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(G1326gat));
  OAI21_X1  g404(.A(G22gat), .B1(new_n579_), .B2(new_n475_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT42), .ZN(new_n607_));
  INV_X1    g406(.A(G22gat), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n570_), .A2(new_n608_), .A3(new_n474_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(G1327gat));
  NOR2_X1   g409(.A1(new_n576_), .A2(new_n577_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(new_n366_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT99), .B1(new_n575_), .B2(new_n565_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n613_), .B1(new_n614_), .B2(new_n567_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(G29gat), .B1(new_n616_), .B2(new_n411_), .ZN(new_n617_));
  OAI21_X1  g416(.A(KEYINPUT43), .B1(new_n291_), .B2(KEYINPUT102), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n619_), .B1(new_n539_), .B2(new_n291_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n527_), .A2(new_n528_), .B1(new_n411_), .B2(new_n534_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n537_), .B1(new_n621_), .B2(new_n530_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n292_), .B(new_n618_), .C1(new_n622_), .C2(new_n517_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n624_), .A2(KEYINPUT44), .A3(new_n337_), .A4(new_n578_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n625_), .A2(G29gat), .A3(new_n411_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n577_), .B1(new_n620_), .B2(new_n623_), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT44), .B1(new_n627_), .B2(new_n578_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n617_), .B1(new_n626_), .B2(new_n629_), .ZN(G1328gat));
  INV_X1    g429(.A(KEYINPUT46), .ZN(new_n631_));
  INV_X1    g430(.A(new_n625_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n632_), .A2(new_n628_), .A3(new_n516_), .ZN(new_n633_));
  INV_X1    g432(.A(G36gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT45), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n515_), .B(KEYINPUT103), .Z(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(G36gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n636_), .B1(new_n616_), .B2(new_n638_), .ZN(new_n639_));
  NOR4_X1   g438(.A1(new_n615_), .A2(KEYINPUT45), .A3(G36gat), .A4(new_n637_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n631_), .B1(new_n635_), .B2(new_n641_), .ZN(new_n642_));
  OAI221_X1 g441(.A(KEYINPUT46), .B1(new_n639_), .B2(new_n640_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1329gat));
  INV_X1    g443(.A(G43gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n615_), .B2(new_n478_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n478_), .A2(new_n645_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n625_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n648_), .B2(new_n628_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT104), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n646_), .B(new_n651_), .C1(new_n648_), .C2(new_n628_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n650_), .A2(KEYINPUT47), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT47), .B1(new_n650_), .B2(new_n652_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1330gat));
  AOI21_X1  g454(.A(G50gat), .B1(new_n616_), .B2(new_n474_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n632_), .A2(new_n208_), .A3(new_n475_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(new_n629_), .ZN(G1331gat));
  NOR2_X1   g457(.A1(new_n367_), .A2(new_n565_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n575_), .A2(new_n659_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n660_), .A2(new_n292_), .A3(new_n337_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n308_), .A3(new_n411_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .A4(new_n659_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G57gat), .B1(new_n663_), .B2(new_n412_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1332gat));
  OAI21_X1  g464(.A(G64gat), .B1(new_n663_), .B2(new_n637_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT48), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n637_), .A2(G64gat), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT105), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n661_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(G1333gat));
  INV_X1    g470(.A(G71gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n661_), .A2(new_n672_), .A3(new_n454_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G71gat), .B1(new_n663_), .B2(new_n478_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT106), .Z(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(KEYINPUT49), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(KEYINPUT49), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(G1334gat));
  OAI21_X1  g477(.A(G78gat), .B1(new_n663_), .B2(new_n475_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT50), .ZN(new_n680_));
  INV_X1    g479(.A(G78gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n661_), .A2(new_n681_), .A3(new_n474_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(G1335gat));
  NOR2_X1   g482(.A1(new_n660_), .A2(new_n612_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G85gat), .B1(new_n684_), .B2(new_n411_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n627_), .A2(new_n659_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n411_), .A2(G85gat), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT107), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n685_), .B1(new_n686_), .B2(new_n688_), .ZN(G1336gat));
  INV_X1    g488(.A(G92gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n684_), .A2(new_n690_), .A3(new_n515_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n637_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n686_), .A2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n693_), .B2(new_n690_), .ZN(G1337gat));
  INV_X1    g493(.A(KEYINPUT108), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n627_), .A2(new_n454_), .A3(new_n659_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G99gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n684_), .A2(new_n454_), .A3(new_n218_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n695_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n697_), .A2(new_n695_), .A3(new_n698_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n700_), .A2(KEYINPUT51), .A3(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT51), .B1(new_n700_), .B2(new_n701_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1338gat));
  NAND4_X1  g503(.A1(new_n624_), .A2(new_n474_), .A3(new_n337_), .A4(new_n659_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n627_), .A2(KEYINPUT109), .A3(new_n474_), .A4(new_n659_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n219_), .B1(KEYINPUT110), .B2(KEYINPUT52), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n711_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .A4(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n684_), .A2(new_n219_), .A3(new_n474_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n712_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT53), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT53), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n712_), .A2(new_n718_), .A3(new_n714_), .A4(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1339gat));
  NOR3_X1   g519(.A1(new_n412_), .A2(new_n476_), .A3(new_n515_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT115), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n546_), .A2(new_n547_), .A3(new_n554_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n559_), .B1(new_n553_), .B2(new_n548_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n560_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(new_n363_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n340_), .B1(new_n249_), .B2(new_n260_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n353_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n346_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n348_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(KEYINPUT113), .A3(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT113), .B1(new_n732_), .B2(new_n733_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n354_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n350_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n730_), .A2(new_n731_), .A3(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n739_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(KEYINPUT112), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n354_), .A2(KEYINPUT55), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n740_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  OAI211_X1 g547(.A(KEYINPUT56), .B(new_n362_), .C1(new_n737_), .C2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n751_));
  INV_X1    g550(.A(new_n346_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n345_), .A2(new_n752_), .A3(new_n353_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n751_), .B1(new_n753_), .B2(new_n348_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n734_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756_));
  NOR4_X1   g555(.A1(new_n345_), .A2(new_n351_), .A3(new_n756_), .A4(new_n353_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n744_), .A2(new_n745_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(new_n738_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n759_), .A3(new_n746_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT56), .B1(new_n760_), .B2(new_n362_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n750_), .A2(new_n761_), .A3(KEYINPUT114), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n357_), .A2(new_n361_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n565_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n362_), .B1(new_n737_), .B2(new_n748_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n729_), .B1(new_n762_), .B2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT57), .B1(new_n771_), .B2(new_n576_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n768_), .A2(new_n769_), .A3(new_n749_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n764_), .B1(new_n761_), .B2(KEYINPUT114), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n728_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT57), .ZN(new_n776_));
  INV_X1    g575(.A(new_n576_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n723_), .B1(new_n772_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n776_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT115), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n560_), .A2(new_n726_), .A3(new_n763_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n768_), .B2(new_n749_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT58), .ZN(new_n784_));
  INV_X1    g583(.A(new_n782_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n750_), .B2(new_n761_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT58), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n783_), .A2(KEYINPUT116), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n291_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n784_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  AOI211_X1 g591(.A(KEYINPUT117), .B(new_n291_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n779_), .B(new_n781_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT118), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n788_), .A2(new_n789_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n292_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT117), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n790_), .A2(new_n791_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n784_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n779_), .A4(new_n781_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n795_), .A2(new_n802_), .A3(new_n337_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT54), .B1(new_n368_), .B2(new_n565_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n338_), .A2(new_n805_), .A3(new_n566_), .A4(new_n367_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n722_), .B1(new_n803_), .B2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(G113gat), .B1(new_n808_), .B2(new_n565_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT119), .ZN(new_n810_));
  INV_X1    g609(.A(new_n807_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n577_), .B1(new_n794_), .B2(KEYINPUT118), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n802_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT59), .B1(new_n813_), .B2(new_n722_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n772_), .A2(new_n778_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n800_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n807_), .B1(new_n816_), .B2(new_n577_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n722_), .A2(KEYINPUT59), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n814_), .A2(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n565_), .A2(G113gat), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n810_), .B1(new_n820_), .B2(new_n821_), .ZN(G1340gat));
  INV_X1    g621(.A(KEYINPUT121), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n367_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n824_), .B(new_n825_), .C1(new_n808_), .C2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n825_), .B1(new_n814_), .B2(new_n824_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n373_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n367_), .A2(G120gat), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(KEYINPUT60), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(KEYINPUT60), .B2(new_n373_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n808_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n823_), .B1(new_n830_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n829_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(G120gat), .A3(new_n827_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(KEYINPUT121), .A3(new_n834_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(G1341gat));
  INV_X1    g639(.A(G127gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n808_), .A2(new_n841_), .A3(new_n577_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n820_), .A2(new_n577_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n844_), .B2(new_n841_), .ZN(G1342gat));
  INV_X1    g644(.A(G134gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n808_), .A2(new_n846_), .A3(new_n777_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n820_), .A2(new_n292_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n849_), .B2(new_n846_), .ZN(G1343gat));
  NOR4_X1   g649(.A1(new_n813_), .A2(new_n412_), .A3(new_n479_), .A4(new_n692_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n565_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT122), .B(G141gat), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1344gat));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n366_), .ZN(new_n855_));
  XOR2_X1   g654(.A(KEYINPUT123), .B(G148gat), .Z(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1345gat));
  NAND2_X1  g656(.A1(new_n851_), .A2(new_n577_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT61), .B(G155gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1346gat));
  INV_X1    g659(.A(G162gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n851_), .A2(new_n861_), .A3(new_n777_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n851_), .A2(new_n292_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n861_), .ZN(G1347gat));
  NAND2_X1  g663(.A1(new_n412_), .A2(new_n692_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  AND4_X1   g665(.A1(new_n475_), .A2(new_n817_), .A3(new_n454_), .A4(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n430_), .B1(new_n867_), .B2(new_n565_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n868_), .A2(KEYINPUT62), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(KEYINPUT62), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n867_), .A2(new_n565_), .A3(new_n413_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .ZN(G1348gat));
  AOI21_X1  g671(.A(G176gat), .B1(new_n867_), .B2(new_n366_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n813_), .A2(new_n474_), .ZN(new_n874_));
  NOR4_X1   g673(.A1(new_n865_), .A2(new_n414_), .A3(new_n478_), .A4(new_n367_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(G1349gat));
  NAND4_X1  g675(.A1(new_n874_), .A2(new_n454_), .A3(new_n577_), .A4(new_n866_), .ZN(new_n877_));
  INV_X1    g676(.A(G183gat), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n577_), .A2(new_n483_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n877_), .A2(new_n878_), .B1(new_n867_), .B2(new_n879_), .ZN(G1350gat));
  NAND2_X1  g679(.A1(new_n867_), .A2(new_n292_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(G190gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n867_), .A2(new_n428_), .A3(new_n777_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1351gat));
  NAND2_X1  g683(.A1(new_n803_), .A2(new_n807_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n865_), .A2(new_n479_), .ZN(new_n886_));
  AOI21_X1  g685(.A(KEYINPUT124), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888_));
  INV_X1    g687(.A(new_n886_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n813_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  OAI211_X1 g689(.A(G197gat), .B(new_n565_), .C1(new_n887_), .C2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n885_), .A2(KEYINPUT124), .A3(new_n886_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n888_), .B1(new_n813_), .B2(new_n889_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n896_), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n565_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n893_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n896_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n558_), .B1(new_n899_), .B2(new_n566_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT126), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n902_), .B(new_n558_), .C1(new_n899_), .C2(new_n566_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n898_), .B1(new_n901_), .B2(new_n903_), .ZN(G1352gat));
  NOR2_X1   g703(.A1(new_n899_), .A2(new_n367_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n906_), .A2(G204gat), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(G204gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n905_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n905_), .B2(new_n908_), .ZN(G1353gat));
  NAND2_X1  g709(.A1(new_n896_), .A2(new_n577_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  AND2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n911_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n911_), .B2(new_n912_), .ZN(G1354gat));
  OR3_X1    g714(.A1(new_n899_), .A2(G218gat), .A3(new_n576_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G218gat), .B1(new_n899_), .B2(new_n291_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1355gat));
endmodule


