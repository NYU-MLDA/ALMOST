//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_;
  INV_X1    g000(.A(G228gat), .ZN(new_n202_));
  INV_X1    g001(.A(G233gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT88), .B(G211gat), .Z(new_n205_));
  INV_X1    g004(.A(G218gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT88), .B(G211gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G218gat), .ZN(new_n209_));
  XOR2_X1   g008(.A(G197gat), .B(G204gat), .Z(new_n210_));
  OAI211_X1 g009(.A(new_n207_), .B(new_n209_), .C1(KEYINPUT21), .C2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(KEYINPUT89), .A3(KEYINPUT21), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n212_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(new_n209_), .A3(new_n207_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT83), .ZN(new_n218_));
  AND2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  INV_X1    g018(.A(G141gat), .ZN(new_n220_));
  INV_X1    g019(.A(G148gat), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n219_), .A2(KEYINPUT1), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G155gat), .B(G162gat), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n218_), .B(new_n222_), .C1(KEYINPUT1), .C2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT84), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n223_), .A2(KEYINPUT1), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT84), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(new_n218_), .A4(new_n222_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n217_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n220_), .A2(new_n221_), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n230_), .A2(KEYINPUT2), .B1(new_n231_), .B2(KEYINPUT3), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT83), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n217_), .B(new_n233_), .ZN(new_n234_));
  OAI221_X1 g033(.A(new_n232_), .B1(KEYINPUT3), .B2(new_n231_), .C1(new_n234_), .C2(KEYINPUT2), .ZN(new_n235_));
  INV_X1    g034(.A(new_n223_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n229_), .A2(new_n237_), .ZN(new_n238_));
  AOI211_X1 g037(.A(new_n204_), .B(new_n216_), .C1(new_n238_), .C2(KEYINPUT29), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT91), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n216_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n213_), .A2(KEYINPUT91), .A3(new_n215_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n242_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT92), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n204_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n246_), .B2(new_n204_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n240_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G78gat), .B(G106gat), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(KEYINPUT93), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n253_), .B(new_n240_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G22gat), .B(G50gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT86), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n256_), .B1(new_n238_), .B2(KEYINPUT29), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n225_), .A2(new_n228_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259_));
  INV_X1    g058(.A(new_n256_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n257_), .A2(new_n263_), .A3(new_n261_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n254_), .A2(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n252_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n267_), .B(KEYINPUT87), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n246_), .A2(new_n204_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT92), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n246_), .A2(new_n247_), .A3(new_n204_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n239_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(new_n253_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n254_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n270_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT94), .ZN(new_n278_));
  INV_X1    g077(.A(new_n253_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n250_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n254_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT94), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(new_n270_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n269_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G225gat), .A2(G233gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n287_));
  XOR2_X1   g086(.A(G127gat), .B(G134gat), .Z(new_n288_));
  XOR2_X1   g087(.A(G113gat), .B(G120gat), .Z(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  NAND3_X1  g089(.A1(new_n238_), .A2(new_n287_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n238_), .A2(new_n290_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n290_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n258_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n286_), .B(new_n291_), .C1(new_n295_), .C2(new_n287_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n294_), .A3(new_n285_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G1gat), .B(G29gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(G85gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT0), .B(G57gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n296_), .A2(new_n297_), .A3(new_n302_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT24), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  MUX2_X1   g108(.A(new_n308_), .B(KEYINPUT24), .S(new_n309_), .Z(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT26), .B(G190gat), .ZN(new_n311_));
  INV_X1    g110(.A(G183gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT25), .B1(new_n312_), .B2(KEYINPUT75), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n312_), .A2(KEYINPUT25), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n311_), .B(new_n313_), .C1(new_n314_), .C2(KEYINPUT75), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(G183gat), .B2(G190gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n318_), .B1(new_n321_), .B2(new_n317_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n316_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n321_), .B2(KEYINPUT23), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(G169gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT22), .B1(new_n329_), .B2(KEYINPUT77), .ZN(new_n330_));
  INV_X1    g129(.A(G176gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT22), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(G169gat), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n330_), .B(new_n331_), .C1(KEYINPUT77), .C2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n307_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT78), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n328_), .A2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n335_), .A2(KEYINPUT78), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n323_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT30), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT80), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G227gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(G15gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(G71gat), .ZN(new_n346_));
  INV_X1    g145(.A(G99gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT79), .B(G43gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n342_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n350_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n352_), .B1(new_n353_), .B2(new_n341_), .ZN(new_n354_));
  XOR2_X1   g153(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n355_));
  XOR2_X1   g154(.A(new_n355_), .B(KEYINPUT82), .Z(new_n356_));
  XNOR2_X1  g155(.A(new_n290_), .B(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  OR3_X1    g157(.A1(new_n351_), .A2(new_n354_), .A3(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n358_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n306_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT27), .ZN(new_n362_));
  INV_X1    g161(.A(new_n216_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n329_), .A2(KEYINPUT22), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n333_), .A2(new_n364_), .ZN(new_n365_));
  OAI221_X1 g164(.A(new_n307_), .B1(G176gat), .B2(new_n365_), .C1(new_n322_), .C2(new_n326_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT25), .B(G183gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT96), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n311_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n325_), .B(new_n310_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n363_), .A2(new_n372_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n216_), .B(new_n323_), .C1(new_n338_), .C2(new_n337_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n373_), .A2(new_n374_), .A3(KEYINPUT20), .A4(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT20), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n339_), .B2(new_n363_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n216_), .A2(new_n366_), .A3(new_n371_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n377_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G8gat), .B(G36gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(G64gat), .B(G92gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  NOR3_X1   g187(.A1(new_n379_), .A2(new_n383_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n388_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n381_), .A2(new_n382_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n377_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n390_), .B1(new_n393_), .B2(new_n378_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n362_), .B1(new_n389_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n245_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT91), .B1(new_n213_), .B2(new_n215_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n366_), .B(new_n371_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n392_), .B1(new_n398_), .B2(new_n381_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n373_), .A2(new_n374_), .A3(KEYINPUT20), .A4(new_n392_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT100), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n381_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n377_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT100), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n388_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n388_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT27), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n395_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT102), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT102), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n395_), .B(new_n412_), .C1(new_n407_), .C2(new_n409_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n284_), .A2(new_n361_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT98), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n305_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n393_), .A2(new_n378_), .A3(new_n390_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n408_), .A3(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n285_), .B(new_n291_), .C1(new_n295_), .C2(new_n287_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n421_), .B(new_n303_), .C1(new_n285_), .C2(new_n295_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n296_), .A2(new_n297_), .A3(KEYINPUT33), .A4(new_n302_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n416_), .B1(new_n420_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n389_), .A2(new_n394_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(KEYINPUT98), .A4(new_n418_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n388_), .A2(KEYINPUT32), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n405_), .B1(new_n404_), .B2(new_n400_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n399_), .A2(KEYINPUT100), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n430_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT99), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT99), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n437_), .B(new_n430_), .C1(new_n379_), .C2(new_n383_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n434_), .A2(new_n439_), .A3(new_n306_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT101), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT101), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n434_), .A2(new_n439_), .A3(new_n442_), .A4(new_n306_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n429_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n284_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n269_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n281_), .A2(new_n282_), .A3(new_n270_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n282_), .B1(new_n281_), .B2(new_n270_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n306_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n450_), .B(new_n395_), .C1(new_n407_), .C2(new_n409_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n445_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n359_), .A2(new_n360_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n415_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G29gat), .B(G36gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G43gat), .B(G50gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT15), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G15gat), .B(G22gat), .ZN(new_n463_));
  INV_X1    g262(.A(G1gat), .ZN(new_n464_));
  INV_X1    g263(.A(G8gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT14), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G1gat), .B(G8gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n462_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n461_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G229gat), .A2(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT72), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n469_), .B(new_n471_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n475_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT72), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n470_), .A2(new_n479_), .A3(new_n474_), .A4(new_n472_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n476_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G113gat), .B(G141gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT73), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G169gat), .B(G197gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n485_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n476_), .A2(new_n478_), .A3(new_n480_), .A4(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT74), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n458_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT37), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT70), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n494_), .B(KEYINPUT71), .Z(new_n495_));
  INV_X1    g294(.A(G106gat), .ZN(new_n496_));
  AND2_X1   g295(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT64), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT64), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n496_), .B1(new_n500_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT6), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(G99gat), .A3(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(G85gat), .ZN(new_n510_));
  INV_X1    g309(.A(G92gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(KEYINPUT9), .A3(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n513_), .A2(KEYINPUT9), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n509_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT65), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n504_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n501_), .A2(KEYINPUT64), .A3(new_n502_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n499_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n520_));
  AOI21_X1  g319(.A(G106gat), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n509_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT65), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT7), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(new_n347_), .A3(new_n496_), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT66), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT66), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n526_), .A2(new_n530_), .A3(new_n527_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n509_), .A3(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n512_), .A2(new_n513_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n533_), .A2(KEYINPUT8), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n506_), .A2(new_n508_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n535_), .B2(new_n528_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT8), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n532_), .A2(new_n534_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n524_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n462_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G232gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT34), .ZN(new_n542_));
  OAI221_X1 g341(.A(new_n540_), .B1(KEYINPUT35), .B2(new_n542_), .C1(new_n471_), .C2(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(KEYINPUT35), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G190gat), .B(G218gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G134gat), .B(G162gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(KEYINPUT36), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n543_), .A2(new_n545_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n546_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n549_), .B(KEYINPUT36), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n546_), .B2(new_n551_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n493_), .A2(KEYINPUT70), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n495_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n495_), .ZN(new_n560_));
  NOR4_X1   g359(.A1(new_n552_), .A2(new_n555_), .A3(new_n557_), .A4(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G57gat), .B(G64gat), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n564_), .A2(KEYINPUT11), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(KEYINPUT11), .ZN(new_n566_));
  XOR2_X1   g365(.A(G71gat), .B(G78gat), .Z(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n566_), .A2(new_n567_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n469_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n574_));
  XOR2_X1   g373(.A(G127gat), .B(G155gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT16), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  OR3_X1    g377(.A1(new_n573_), .A2(new_n574_), .A3(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(KEYINPUT17), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n573_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n563_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585_));
  INV_X1    g384(.A(new_n570_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n539_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n524_), .A2(new_n570_), .A3(new_n538_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n585_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT67), .Z(new_n590_));
  NAND2_X1  g389(.A1(KEYINPUT68), .A2(KEYINPUT12), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT68), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n539_), .A2(new_n586_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n594_), .ZN(new_n596_));
  AOI211_X1 g395(.A(new_n596_), .B(new_n570_), .C1(new_n524_), .C2(new_n538_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n592_), .B(new_n585_), .C1(new_n595_), .C2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n590_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G120gat), .B(G148gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT5), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n603_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n590_), .A2(new_n598_), .A3(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n607_));
  AND3_X1   g406(.A1(new_n604_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT13), .ZN(new_n609_));
  AOI22_X1  g408(.A1(new_n604_), .A2(new_n606_), .B1(KEYINPUT69), .B2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n584_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n492_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n464_), .A3(new_n306_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT38), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n556_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n489_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n611_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(new_n583_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n458_), .A2(new_n618_), .A3(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n623_), .B2(new_n450_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n615_), .A2(new_n616_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n617_), .A2(new_n624_), .A3(new_n625_), .ZN(G1324gat));
  OAI21_X1  g425(.A(G8gat), .B1(new_n623_), .B2(new_n414_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT39), .ZN(new_n628_));
  INV_X1    g427(.A(new_n414_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n614_), .A2(new_n465_), .A3(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n628_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1325gat));
  OAI21_X1  g433(.A(G15gat), .B1(new_n623_), .B2(new_n456_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT41), .Z(new_n636_));
  NAND3_X1  g435(.A1(new_n614_), .A2(new_n344_), .A3(new_n455_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1326gat));
  XNOR2_X1  g437(.A(new_n449_), .B(KEYINPUT104), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  OR3_X1    g439(.A1(new_n613_), .A2(G22gat), .A3(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n642_));
  INV_X1    g441(.A(new_n623_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n639_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n642_), .B1(new_n644_), .B2(G22gat), .ZN(new_n645_));
  OAI211_X1 g444(.A(G22gat), .B(new_n642_), .C1(new_n623_), .C2(new_n640_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n641_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT106), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n641_), .B(new_n650_), .C1(new_n645_), .C2(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(G1327gat));
  NAND2_X1  g451(.A1(new_n556_), .A2(new_n582_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n611_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n492_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n306_), .ZN(new_n657_));
  OAI21_X1  g456(.A(KEYINPUT43), .B1(new_n457_), .B2(new_n563_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n455_), .B1(new_n445_), .B2(new_n453_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n659_), .B(new_n562_), .C1(new_n660_), .C2(new_n415_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n620_), .A2(new_n582_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT44), .B1(new_n662_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  AOI211_X1 g465(.A(new_n666_), .B(new_n663_), .C1(new_n658_), .C2(new_n661_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n306_), .A2(G29gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n657_), .B1(new_n668_), .B2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  INV_X1    g470(.A(G36gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n668_), .B2(new_n629_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n414_), .A2(G36gat), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n674_), .B1(new_n655_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n674_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n492_), .A2(new_n654_), .A3(new_n678_), .A4(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n671_), .B1(new_n673_), .B2(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n677_), .A2(new_n679_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n665_), .A2(new_n667_), .A3(new_n414_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n682_), .B(KEYINPUT46), .C1(new_n672_), .C2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(G1329gat));
  NAND2_X1  g484(.A1(new_n455_), .A2(G43gat), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n665_), .A2(new_n667_), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G43gat), .B1(new_n656_), .B2(new_n455_), .ZN(new_n688_));
  OR3_X1    g487(.A1(new_n687_), .A2(new_n688_), .A3(KEYINPUT47), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT47), .B1(new_n687_), .B2(new_n688_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1330gat));
  AOI21_X1  g490(.A(G50gat), .B1(new_n656_), .B2(new_n639_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n449_), .A2(G50gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n668_), .B2(new_n693_), .ZN(G1331gat));
  NOR2_X1   g493(.A1(new_n491_), .A2(new_n582_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n458_), .A2(new_n611_), .A3(new_n618_), .A4(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G57gat), .B1(new_n696_), .B2(new_n450_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n608_), .A2(new_n610_), .ZN(new_n698_));
  OR4_X1    g497(.A1(new_n457_), .A2(new_n489_), .A3(new_n698_), .A4(new_n584_), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n450_), .A2(G57gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n697_), .B1(new_n699_), .B2(new_n700_), .ZN(G1332gat));
  OAI21_X1  g500(.A(G64gat), .B1(new_n696_), .B2(new_n414_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT48), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n414_), .A2(G64gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n699_), .B2(new_n704_), .ZN(G1333gat));
  OAI21_X1  g504(.A(G71gat), .B1(new_n696_), .B2(new_n456_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT49), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n456_), .A2(G71gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n699_), .B2(new_n708_), .ZN(G1334gat));
  OAI21_X1  g508(.A(G78gat), .B1(new_n696_), .B2(new_n640_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT50), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n640_), .A2(G78gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n699_), .B2(new_n712_), .ZN(G1335gat));
  NOR2_X1   g512(.A1(new_n698_), .A2(new_n653_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n458_), .A2(new_n619_), .A3(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT108), .ZN(new_n716_));
  AOI21_X1  g515(.A(G85gat), .B1(new_n716_), .B2(new_n306_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n611_), .A2(new_n619_), .A3(new_n582_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n662_), .A2(KEYINPUT109), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n658_), .A2(new_n720_), .A3(new_n661_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n718_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n306_), .A2(G85gat), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT110), .Z(new_n724_));
  AOI21_X1  g523(.A(new_n717_), .B1(new_n722_), .B2(new_n724_), .ZN(G1336gat));
  NAND3_X1  g524(.A1(new_n716_), .A2(new_n511_), .A3(new_n629_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n722_), .A2(new_n629_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(new_n511_), .ZN(G1337gat));
  NAND2_X1  g527(.A1(new_n722_), .A2(new_n455_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(G99gat), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n456_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n716_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(new_n731_), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n347_), .B1(new_n722_), .B2(new_n455_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n733_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT51), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(G1338gat));
  NAND3_X1  g537(.A1(new_n716_), .A2(new_n496_), .A3(new_n449_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n718_), .A2(new_n284_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n496_), .B1(new_n662_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n741_), .A2(new_n742_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n739_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT53), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n739_), .B(new_n747_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1339gat));
  AND2_X1   g548(.A1(new_n606_), .A2(new_n489_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n588_), .A2(new_n591_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n587_), .A2(new_n596_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n539_), .A2(new_n593_), .A3(new_n594_), .A4(new_n586_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n751_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT55), .B1(new_n754_), .B2(new_n585_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n598_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n592_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758_));
  INV_X1    g557(.A(new_n585_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n756_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT56), .B1(new_n762_), .B2(new_n603_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n758_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n598_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OAI211_X1 g565(.A(KEYINPUT56), .B(new_n603_), .C1(new_n766_), .C2(new_n760_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n750_), .B1(new_n763_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n604_), .A2(new_n606_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n487_), .B1(new_n477_), .B2(new_n474_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(new_n474_), .B2(new_n473_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n488_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT112), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n488_), .A2(new_n775_), .A3(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n770_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n556_), .B1(new_n769_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT57), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT57), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n603_), .B1(new_n766_), .B2(new_n760_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n767_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n786_), .A2(new_n750_), .B1(new_n770_), .B2(new_n777_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT113), .B(new_n782_), .C1(new_n787_), .C2(new_n556_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n781_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n785_), .A2(new_n790_), .A3(new_n767_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n783_), .A2(KEYINPUT114), .A3(new_n784_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n777_), .A2(new_n606_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n791_), .A2(KEYINPUT58), .A3(new_n792_), .A4(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n562_), .ZN(new_n795_));
  XOR2_X1   g594(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n796_));
  NAND3_X1  g595(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(KEYINPUT115), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n791_), .A2(new_n799_), .A3(new_n792_), .A4(new_n793_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n795_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n582_), .B1(new_n789_), .B2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n695_), .B(KEYINPUT111), .C1(new_n608_), .C2(new_n610_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n563_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT111), .B1(new_n698_), .B2(new_n695_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT54), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n807_));
  INV_X1    g606(.A(new_n695_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n611_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n563_), .A4(new_n803_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n806_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n802_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n284_), .A2(new_n455_), .A3(new_n306_), .A4(new_n414_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n814_), .A2(KEYINPUT118), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(KEYINPUT118), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(KEYINPUT59), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n813_), .A2(KEYINPUT119), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT119), .B1(new_n813_), .B2(new_n818_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT59), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n813_), .A2(KEYINPUT117), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n802_), .A2(new_n812_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n817_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n821_), .B(new_n491_), .C1(new_n822_), .C2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G113gat), .ZN(new_n828_));
  INV_X1    g627(.A(new_n826_), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n619_), .A2(G113gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n828_), .B1(new_n829_), .B2(new_n830_), .ZN(G1340gat));
  OAI21_X1  g630(.A(new_n821_), .B1(new_n822_), .B2(new_n826_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G120gat), .B1(new_n832_), .B2(new_n698_), .ZN(new_n833_));
  INV_X1    g632(.A(G120gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n698_), .B2(KEYINPUT60), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n826_), .B(new_n835_), .C1(KEYINPUT60), .C2(new_n834_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n836_), .ZN(G1341gat));
  NAND2_X1  g636(.A1(new_n823_), .A2(new_n825_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n817_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n583_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(G127gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n840_), .A2(KEYINPUT120), .A3(new_n841_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n820_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n813_), .A2(KEYINPUT119), .A3(new_n818_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(KEYINPUT59), .B2(new_n829_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n582_), .A2(new_n841_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n844_), .A2(new_n845_), .B1(new_n849_), .B2(new_n850_), .ZN(G1342gat));
  OAI21_X1  g650(.A(G134gat), .B1(new_n832_), .B2(new_n563_), .ZN(new_n852_));
  OR3_X1    g651(.A1(new_n829_), .A2(G134gat), .A3(new_n618_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1343gat));
  NOR2_X1   g653(.A1(new_n284_), .A2(new_n455_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n306_), .A3(new_n414_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT121), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n489_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT122), .B(G141gat), .Z(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1344gat));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n611_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g663(.A1(new_n859_), .A2(new_n583_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT61), .B(G155gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  INV_X1    g666(.A(G162gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n859_), .B2(new_n562_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n618_), .A2(G162gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n859_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(KEYINPUT123), .A3(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n874_));
  INV_X1    g673(.A(new_n872_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n869_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n876_), .ZN(G1347gat));
  AND2_X1   g676(.A1(new_n802_), .A2(new_n812_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n414_), .A2(new_n306_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n455_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n639_), .A2(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n878_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n489_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(G169gat), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT124), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n886_), .A3(G169gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n885_), .A2(KEYINPUT62), .A3(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n883_), .A2(new_n365_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n886_), .B1(new_n883_), .B2(G169gat), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n888_), .A2(new_n892_), .ZN(G1348gat));
  AOI21_X1  g692(.A(G176gat), .B1(new_n882_), .B2(new_n611_), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n894_), .A2(KEYINPUT125), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(KEYINPUT125), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n449_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n880_), .A2(new_n331_), .A3(new_n698_), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n895_), .A2(new_n896_), .B1(new_n897_), .B2(new_n898_), .ZN(G1349gat));
  AND3_X1   g698(.A1(new_n882_), .A2(new_n369_), .A3(new_n583_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n897_), .A2(new_n455_), .A3(new_n583_), .A4(new_n879_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n312_), .ZN(G1350gat));
  NAND3_X1  g701(.A1(new_n882_), .A2(new_n311_), .A3(new_n556_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n878_), .A2(new_n563_), .A3(new_n881_), .ZN(new_n904_));
  INV_X1    g703(.A(G190gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT126), .ZN(G1351gat));
  NAND2_X1  g706(.A1(new_n855_), .A2(new_n879_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n802_), .A2(new_n824_), .A3(new_n812_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n824_), .B1(new_n802_), .B2(new_n812_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT127), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT127), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n914_), .B(new_n909_), .C1(new_n910_), .C2(new_n911_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G197gat), .B1(new_n916_), .B2(new_n489_), .ZN(new_n917_));
  INV_X1    g716(.A(G197gat), .ZN(new_n918_));
  AOI211_X1 g717(.A(new_n918_), .B(new_n619_), .C1(new_n913_), .C2(new_n915_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1352gat));
  AOI21_X1  g719(.A(new_n914_), .B1(new_n838_), .B2(new_n909_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n915_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n611_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(G204gat), .ZN(new_n924_));
  INV_X1    g723(.A(G204gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n916_), .A2(new_n925_), .A3(new_n611_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1353gat));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n582_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n916_), .B2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n930_), .ZN(new_n932_));
  AOI211_X1 g731(.A(new_n928_), .B(new_n932_), .C1(new_n913_), .C2(new_n915_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n931_), .A2(new_n933_), .ZN(G1354gat));
  NAND3_X1  g733(.A1(new_n916_), .A2(new_n206_), .A3(new_n556_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n563_), .B1(new_n913_), .B2(new_n915_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n206_), .B2(new_n936_), .ZN(G1355gat));
endmodule


