//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_;
  NAND2_X1  g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G85gat), .A2(G92gat), .ZN(new_n204_));
  NOR3_X1   g003(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT67), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT67), .ZN(new_n206_));
  INV_X1    g005(.A(G85gat), .ZN(new_n207_));
  INV_X1    g006(.A(G92gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n206_), .B1(new_n209_), .B2(new_n202_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n205_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  OR3_X1    g015(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI211_X1 g019(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n216_), .A2(new_n217_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n211_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT8), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT8), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n211_), .A2(new_n222_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT10), .ZN(new_n228_));
  INV_X1    g027(.A(G99gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n230_), .A2(KEYINPUT64), .A3(new_n231_), .A4(new_n232_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n209_), .A2(KEYINPUT9), .A3(new_n202_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n202_), .A2(KEYINPUT9), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n216_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT65), .B1(new_n237_), .B2(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n216_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n227_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G29gat), .B(G36gat), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n247_), .A2(KEYINPUT69), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(KEYINPUT69), .ZN(new_n249_));
  XOR2_X1   g048(.A(G43gat), .B(G50gat), .Z(new_n250_));
  OR3_X1    g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n250_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n246_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G232gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT34), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT35), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n253_), .B(KEYINPUT15), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n260_), .B1(new_n262_), .B2(new_n246_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(KEYINPUT70), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n257_), .A2(new_n258_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n267_));
  INV_X1    g066(.A(new_n265_), .ZN(new_n268_));
  OAI221_X1 g067(.A(new_n260_), .B1(KEYINPUT70), .B2(new_n268_), .C1(new_n262_), .C2(new_n246_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G190gat), .B(G218gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G134gat), .B(G162gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(KEYINPUT36), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n266_), .A2(new_n267_), .A3(new_n269_), .A4(new_n274_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n266_), .A2(new_n269_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n273_), .A2(KEYINPUT36), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT37), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT37), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n278_), .A2(new_n281_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G57gat), .B(G64gat), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n287_), .A2(KEYINPUT11), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(KEYINPUT11), .ZN(new_n289_));
  XOR2_X1   g088(.A(G71gat), .B(G78gat), .Z(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n289_), .A2(new_n290_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G231gat), .A2(G233gat), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n293_), .B(new_n294_), .Z(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT72), .B(G8gat), .ZN(new_n296_));
  INV_X1    g095(.A(G1gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT14), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G15gat), .B(G22gat), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G1gat), .B(G8gat), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n301_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n295_), .B(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G127gat), .B(G155gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT16), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G183gat), .B(G211gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT17), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n306_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n295_), .B(new_n304_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n310_), .B(KEYINPUT17), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT73), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n286_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G120gat), .B(G148gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT5), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G176gat), .B(G204gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  NAND2_X1  g125(.A1(G230gat), .A2(G233gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n227_), .A2(new_n245_), .A3(new_n293_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n293_), .B1(new_n227_), .B2(new_n245_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT68), .ZN(new_n332_));
  AND2_X1   g131(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT64), .B1(new_n335_), .B2(new_n231_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n236_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n243_), .B1(new_n338_), .B2(new_n242_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n237_), .A2(KEYINPUT65), .A3(new_n240_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n211_), .A2(new_n222_), .A3(new_n225_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n225_), .B1(new_n211_), .B2(new_n222_), .ZN(new_n342_));
  OAI22_X1  g141(.A1(new_n339_), .A2(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n293_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n227_), .A2(new_n245_), .A3(new_n293_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(KEYINPUT12), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT12), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n330_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n328_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n326_), .B1(new_n332_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n332_), .A2(new_n350_), .A3(new_n326_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT13), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT13), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n356_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n322_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(G71gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT80), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT23), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT79), .B(KEYINPUT23), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n366_), .B2(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(KEYINPUT77), .B(G190gat), .Z(new_n371_));
  OAI21_X1  g170(.A(new_n370_), .B1(G183gat), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT22), .ZN(new_n374_));
  INV_X1    g173(.A(G176gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377_));
  AOI22_X1  g176(.A1(new_n376_), .A2(G169gat), .B1(new_n377_), .B2(new_n374_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n372_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n369_), .A2(new_n366_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n380_), .B1(new_n367_), .B2(KEYINPUT23), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT24), .ZN(new_n383_));
  MUX2_X1   g182(.A(new_n383_), .B(KEYINPUT24), .S(new_n377_), .Z(new_n384_));
  AND2_X1   g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT25), .B(G183gat), .ZN(new_n386_));
  AND2_X1   g185(.A1(KEYINPUT78), .A2(KEYINPUT26), .ZN(new_n387_));
  OAI21_X1  g186(.A(G190gat), .B1(KEYINPUT78), .B2(KEYINPUT26), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT26), .ZN(new_n389_));
  OAI221_X1 g188(.A(new_n386_), .B1(new_n387_), .B2(new_n388_), .C1(new_n371_), .C2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n385_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n379_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n372_), .A2(new_n378_), .B1(new_n385_), .B2(new_n390_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n393_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n395_), .A2(new_n229_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n229_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n365_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n400_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n364_), .A3(new_n398_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n361_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G127gat), .B(G134gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G113gat), .B(G120gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(new_n409_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n413_), .B(KEYINPUT31), .Z(new_n414_));
  XNOR2_X1  g213(.A(G15gat), .B(G43gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n401_), .A2(new_n403_), .A3(new_n361_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n405_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n416_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n417_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n419_), .B1(new_n420_), .B2(new_n404_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G85gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT0), .B(G57gat), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n425_), .B(new_n426_), .Z(new_n427_));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G155gat), .A2(G162gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n431_), .A2(KEYINPUT1), .ZN(new_n432_));
  NOR2_X1   g231(.A1(G155gat), .A2(G162gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n433_), .B2(KEYINPUT1), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT86), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n432_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OAI211_X1 g235(.A(KEYINPUT86), .B(new_n431_), .C1(new_n433_), .C2(KEYINPUT1), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G141gat), .B(G148gat), .ZN(new_n439_));
  OR2_X1    g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT2), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT3), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n445_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n433_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n431_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n440_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n413_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n440_), .A2(new_n451_), .A3(new_n408_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n430_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT4), .B1(new_n452_), .B2(new_n413_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n429_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n453_), .A2(new_n428_), .A3(new_n454_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n427_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n427_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n460_), .B2(KEYINPUT100), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n457_), .A2(new_n458_), .A3(new_n427_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT100), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT101), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n459_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n457_), .A2(new_n458_), .A3(KEYINPUT100), .A4(new_n427_), .ZN(new_n467_));
  AND4_X1   g266(.A1(KEYINPUT101), .A2(new_n464_), .A3(new_n466_), .A4(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT27), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G211gat), .B(G218gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT21), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(G197gat), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT89), .B1(new_n474_), .B2(G204gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n476_));
  INV_X1    g275(.A(G204gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n477_), .A3(G197gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(G204gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n475_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n473_), .A2(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n480_), .A2(KEYINPUT21), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n482_), .A2(new_n471_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(G197gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n472_), .B1(new_n484_), .B2(new_n479_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT88), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n483_), .A2(KEYINPUT90), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT90), .B1(new_n483_), .B2(new_n486_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n481_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n392_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT94), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT94), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n489_), .A2(new_n492_), .A3(new_n392_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n381_), .B1(G183gat), .B2(G190gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n382_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT22), .B(G169gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n497_), .B2(new_n375_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT26), .B(G190gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n386_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n384_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n370_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT20), .B1(new_n489_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G226gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT19), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n494_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G8gat), .B(G36gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT18), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G64gat), .B(G92gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n512_), .B(new_n513_), .Z(new_n514_));
  INV_X1    g313(.A(KEYINPUT20), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n489_), .B2(new_n505_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n396_), .B(new_n481_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n508_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n510_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n514_), .B1(new_n510_), .B2(new_n519_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n470_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT103), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(KEYINPUT102), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n510_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT102), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n470_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n514_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n508_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT97), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n491_), .A2(new_n493_), .B1(new_n506_), .B2(new_n531_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n506_), .A2(new_n531_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n530_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT98), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n518_), .B2(new_n508_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n516_), .A2(KEYINPUT98), .A3(new_n530_), .A4(new_n517_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n529_), .B1(new_n534_), .B2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n525_), .A2(new_n528_), .A3(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(KEYINPUT103), .B(new_n470_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n469_), .A2(new_n524_), .A3(new_n540_), .A4(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n452_), .A2(KEYINPUT29), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT28), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G22gat), .B(G50gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G78gat), .B(G106gat), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n452_), .A2(KEYINPUT29), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n489_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n489_), .A2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(G228gat), .A2(G233gat), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n552_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n555_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n489_), .B(new_n551_), .C1(new_n553_), .C2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n550_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n548_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(new_n558_), .A3(new_n550_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT93), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n559_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AOI211_X1 g366(.A(KEYINPUT92), .B(new_n550_), .C1(new_n556_), .C2(new_n558_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n563_), .B1(new_n570_), .B2(new_n548_), .ZN(new_n571_));
  AOI211_X1 g370(.A(KEYINPUT93), .B(new_n547_), .C1(new_n567_), .C2(new_n569_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n562_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n423_), .B1(new_n542_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n514_), .A2(KEYINPUT32), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n534_), .B2(new_n538_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT99), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n461_), .A2(new_n464_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT99), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n580_), .B(new_n576_), .C1(new_n534_), .C2(new_n538_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n510_), .A2(new_n519_), .A3(new_n575_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n578_), .A2(new_n579_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n559_), .B1(new_n564_), .B2(new_n561_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n548_), .B1(new_n584_), .B2(new_n568_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT93), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n570_), .A2(new_n563_), .A3(new_n548_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n462_), .B1(KEYINPUT95), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n453_), .A2(new_n454_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n428_), .B1(new_n591_), .B2(KEYINPUT96), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(KEYINPUT96), .B2(new_n591_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n455_), .A2(new_n456_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n427_), .B1(new_n594_), .B2(new_n428_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n590_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n520_), .A2(new_n521_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n462_), .A2(KEYINPUT95), .A3(new_n589_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n583_), .A2(new_n588_), .A3(new_n562_), .A4(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n524_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n573_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n469_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(new_n422_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n574_), .A2(new_n600_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G169gat), .B(G197gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(KEYINPUT76), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n304_), .A2(new_n253_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n261_), .A2(new_n305_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT75), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT75), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n261_), .A2(new_n615_), .A3(new_n305_), .ZN(new_n616_));
  AOI211_X1 g415(.A(new_n610_), .B(new_n612_), .C1(new_n614_), .C2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n304_), .A2(new_n253_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n610_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(new_n611_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n609_), .B1(new_n617_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n614_), .A2(new_n616_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n610_), .A2(new_n612_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n620_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n624_), .B1(KEYINPUT76), .B2(new_n608_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n605_), .A2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n359_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n469_), .A2(G1gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(KEYINPUT104), .A3(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n359_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n631_), .A2(KEYINPUT38), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT106), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n282_), .B(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n605_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n358_), .A2(new_n627_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n317_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT105), .Z(new_n642_));
  AND2_X1   g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n469_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT38), .B1(new_n631_), .B2(new_n634_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(KEYINPUT107), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n648_), .B(KEYINPUT38), .C1(new_n631_), .C2(new_n634_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n635_), .B(new_n645_), .C1(new_n647_), .C2(new_n649_), .ZN(G1324gat));
  NAND3_X1  g449(.A1(new_n629_), .A2(new_n601_), .A3(new_n296_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n643_), .A2(new_n601_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT108), .B(KEYINPUT39), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n652_), .A2(G8gat), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n652_), .B2(G8gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n651_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(G1325gat));
  INV_X1    g457(.A(G15gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n643_), .B2(new_n423_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT41), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n629_), .A2(new_n659_), .A3(new_n423_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1326gat));
  INV_X1    g462(.A(G22gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n664_), .B1(new_n643_), .B2(new_n573_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT42), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n629_), .A2(new_n664_), .A3(new_n573_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1327gat));
  INV_X1    g467(.A(new_n286_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n542_), .A2(new_n573_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n600_), .A3(new_n422_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n602_), .A2(new_n604_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n669_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(KEYINPUT109), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n677_), .B1(new_n605_), .B2(new_n669_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n676_), .A2(new_n678_), .A3(new_n319_), .A4(new_n640_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n318_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n682_), .A2(KEYINPUT44), .A3(new_n640_), .A4(new_n678_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n681_), .A2(G29gat), .A3(new_n603_), .A4(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(G29gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n282_), .A2(new_n319_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(new_n358_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n628_), .A2(KEYINPUT110), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n671_), .A2(new_n672_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n626_), .A3(new_n687_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n688_), .A2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n685_), .B1(new_n693_), .B2(new_n469_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n684_), .A2(new_n694_), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n681_), .A2(new_n601_), .A3(new_n683_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G36gat), .ZN(new_n697_));
  NOR2_X1   g496(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n524_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(G36gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n688_), .A2(new_n692_), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT45), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n688_), .A2(new_n692_), .A3(new_n703_), .A4(new_n700_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n698_), .B1(new_n702_), .B2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT112), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n697_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n697_), .B2(new_n705_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1329gat));
  INV_X1    g508(.A(G43gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n422_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n681_), .A2(new_n683_), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT113), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT113), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n681_), .A2(new_n714_), .A3(new_n683_), .A4(new_n711_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n710_), .B1(new_n693_), .B2(new_n422_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n713_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT47), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n713_), .A2(new_n719_), .A3(new_n715_), .A4(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1330gat));
  NAND4_X1  g520(.A1(new_n681_), .A2(G50gat), .A3(new_n573_), .A4(new_n683_), .ZN(new_n722_));
  INV_X1    g521(.A(G50gat), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n586_), .A2(new_n587_), .B1(new_n561_), .B2(new_n560_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n693_), .B2(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n722_), .A2(new_n725_), .ZN(G1331gat));
  AND2_X1   g525(.A1(new_n355_), .A2(new_n357_), .ZN(new_n727_));
  NOR4_X1   g526(.A1(new_n322_), .A2(new_n605_), .A3(new_n626_), .A4(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(G57gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n729_), .A3(new_n603_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n727_), .A2(new_n626_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n639_), .A2(new_n318_), .A3(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n469_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(G1332gat));
  OAI21_X1  g533(.A(G64gat), .B1(new_n732_), .B2(new_n699_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT48), .ZN(new_n736_));
  INV_X1    g535(.A(G64gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n728_), .A2(new_n737_), .A3(new_n601_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1333gat));
  OAI21_X1  g538(.A(G71gat), .B1(new_n732_), .B2(new_n422_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT49), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n728_), .A2(new_n363_), .A3(new_n423_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1334gat));
  OAI21_X1  g542(.A(G78gat), .B1(new_n732_), .B2(new_n724_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT50), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n724_), .A2(G78gat), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT114), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n728_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n745_), .A2(new_n748_), .ZN(G1335gat));
  NAND3_X1  g548(.A1(new_n682_), .A2(new_n678_), .A3(new_n731_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750_), .B2(new_n469_), .ZN(new_n751_));
  NOR4_X1   g550(.A1(new_n605_), .A2(new_n626_), .A3(new_n727_), .A4(new_n686_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n752_), .A2(new_n207_), .A3(new_n603_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT115), .ZN(G1336gat));
  OAI21_X1  g554(.A(G92gat), .B1(new_n750_), .B2(new_n699_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n752_), .A2(new_n208_), .A3(new_n601_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT116), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n750_), .B2(new_n422_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n752_), .A2(new_n423_), .A3(new_n335_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g562(.A1(new_n752_), .A2(new_n231_), .A3(new_n573_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n682_), .A2(new_n573_), .A3(new_n678_), .A4(new_n731_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(G106gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(G106gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g569(.A1(new_n469_), .A2(new_n422_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n699_), .A2(new_n724_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT121), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT121), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n699_), .A2(new_n771_), .A3(new_n724_), .A4(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n282_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n353_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n626_), .A2(new_n778_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n329_), .A2(new_n330_), .A3(new_n348_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n349_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n327_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n347_), .A2(new_n328_), .A3(new_n349_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(KEYINPUT55), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n327_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n784_), .A2(KEYINPUT118), .A3(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT118), .B1(new_n784_), .B2(new_n786_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n326_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n783_), .A2(KEYINPUT55), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n793_), .A2(new_n350_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n786_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n792_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n784_), .A2(KEYINPUT118), .A3(new_n786_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n326_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n779_), .B1(new_n791_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n354_), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n610_), .A2(new_n611_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n622_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n608_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n619_), .B2(new_n612_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(KEYINPUT119), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n802_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n806_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n808_), .A2(new_n811_), .B1(new_n608_), .B2(new_n624_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n801_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n777_), .B1(new_n800_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n812_), .A2(new_n778_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n326_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n326_), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n790_), .B(new_n819_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n817_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n817_), .B(KEYINPUT58), .C1(new_n818_), .C2(new_n820_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n286_), .A3(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT57), .B(new_n777_), .C1(new_n800_), .C2(new_n813_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n816_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n317_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n816_), .A2(new_n825_), .A3(KEYINPUT120), .A4(new_n826_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n319_), .A2(new_n626_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n727_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n834_), .B1(new_n727_), .B2(new_n833_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n669_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT54), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n727_), .A2(new_n833_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT117), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n286_), .B1(new_n841_), .B2(new_n835_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n839_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n776_), .B1(new_n832_), .B2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(G113gat), .B1(new_n846_), .B2(new_n626_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n846_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT59), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n773_), .A2(KEYINPUT122), .A3(new_n775_), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT122), .B1(new_n773_), .B2(new_n775_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n850_), .A2(new_n851_), .A3(KEYINPUT59), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n842_), .B(KEYINPUT54), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n827_), .A2(new_n319_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n852_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n849_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n626_), .A2(G113gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT123), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n847_), .B1(new_n857_), .B2(new_n859_), .ZN(G1340gat));
  OAI21_X1  g659(.A(G120gat), .B1(new_n856_), .B2(new_n727_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT60), .ZN(new_n862_));
  AOI21_X1  g661(.A(G120gat), .B1(new_n358_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT124), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n862_), .B2(G120gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n863_), .B2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n861_), .B1(new_n848_), .B2(new_n867_), .ZN(G1341gat));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n317_), .B(new_n855_), .C1(new_n846_), .C2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G127gat), .ZN(new_n871_));
  INV_X1    g670(.A(G127gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n846_), .A2(new_n872_), .A3(new_n318_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT125), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT125), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n871_), .A2(new_n876_), .A3(new_n873_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1342gat));
  OAI21_X1  g677(.A(G134gat), .B1(new_n856_), .B2(new_n669_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n637_), .A2(G134gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n848_), .B2(new_n880_), .ZN(G1343gat));
  AOI21_X1  g680(.A(new_n724_), .B1(new_n832_), .B2(new_n845_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n601_), .A2(new_n423_), .A3(new_n469_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n882_), .A2(KEYINPUT126), .A3(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT126), .B1(new_n882_), .B2(new_n883_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n626_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G141gat), .ZN(new_n888_));
  INV_X1    g687(.A(G141gat), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n889_), .B(new_n626_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1344gat));
  OAI21_X1  g690(.A(new_n358_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G148gat), .ZN(new_n893_));
  INV_X1    g692(.A(G148gat), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n894_), .B(new_n358_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(G1345gat));
  OAI21_X1  g695(.A(new_n318_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT61), .B(G155gat), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n898_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n318_), .B(new_n900_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(G1346gat));
  INV_X1    g701(.A(G162gat), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n903_), .B(new_n638_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n886_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n669_), .B1(new_n905_), .B2(new_n884_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n904_), .B1(new_n906_), .B2(new_n903_), .ZN(G1347gat));
  NOR2_X1   g706(.A1(new_n853_), .A2(new_n854_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n699_), .A2(new_n603_), .A3(new_n422_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n724_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n626_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(G169gat), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n912_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n916_));
  INV_X1    g715(.A(new_n497_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n915_), .B(new_n916_), .C1(new_n917_), .C2(new_n912_), .ZN(G1348gat));
  AOI21_X1  g717(.A(G176gat), .B1(new_n911_), .B2(new_n358_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n573_), .B1(new_n832_), .B2(new_n845_), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n909_), .A2(G176gat), .A3(new_n358_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n920_), .B2(new_n921_), .ZN(G1349gat));
  INV_X1    g721(.A(new_n911_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n923_), .A2(new_n386_), .A3(new_n830_), .ZN(new_n924_));
  INV_X1    g723(.A(G183gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n920_), .A2(new_n318_), .A3(new_n909_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n924_), .B1(new_n925_), .B2(new_n926_), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n923_), .B2(new_n669_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n911_), .A2(new_n500_), .A3(new_n638_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1351gat));
  NAND2_X1  g729(.A1(new_n832_), .A2(new_n845_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n573_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n601_), .A2(new_n469_), .A3(new_n422_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n626_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n358_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT63), .B(G211gat), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n932_), .A2(new_n830_), .A3(new_n933_), .ZN(new_n941_));
  MUX2_X1   g740(.A(new_n939_), .B(new_n940_), .S(new_n941_), .Z(G1354gat));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943_));
  INV_X1    g742(.A(G218gat), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n944_), .B1(new_n934_), .B2(new_n286_), .ZN(new_n945_));
  NOR4_X1   g744(.A1(new_n932_), .A2(G218gat), .A3(new_n637_), .A4(new_n933_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n943_), .B1(new_n945_), .B2(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n637_), .A2(G218gat), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n934_), .A2(new_n948_), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n932_), .A2(new_n669_), .A3(new_n933_), .ZN(new_n950_));
  OAI211_X1 g749(.A(new_n949_), .B(KEYINPUT127), .C1(new_n944_), .C2(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n947_), .A2(new_n951_), .ZN(G1355gat));
endmodule


