//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n867_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT94), .B(G197gat), .Z(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(G204gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT21), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(new_n203_), .B2(G204gat), .ZN(new_n208_));
  OAI221_X1 g007(.A(new_n202_), .B1(new_n204_), .B2(new_n206_), .C1(KEYINPUT21), .C2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n202_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(KEYINPUT21), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(KEYINPUT1), .ZN(new_n214_));
  OR2_X1    g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(KEYINPUT1), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT89), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n218_), .B1(new_n217_), .B2(new_n216_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT90), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n214_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(new_n220_), .B2(new_n219_), .ZN(new_n222_));
  INV_X1    g021(.A(G141gat), .ZN(new_n223_));
  INV_X1    g022(.A(G148gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT88), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n223_), .A2(new_n224_), .A3(KEYINPUT88), .ZN(new_n228_));
  AOI22_X1  g027(.A1(new_n227_), .A2(new_n228_), .B1(G141gat), .B2(G148gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n222_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n225_), .A2(KEYINPUT3), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT91), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n234_), .B(new_n235_), .C1(KEYINPUT3), .C2(new_n225_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n213_), .B(new_n215_), .C1(new_n232_), .C2(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n230_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n212_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G228gat), .A2(G233gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n241_), .B(KEYINPUT93), .Z(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G78gat), .B(G106gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT95), .ZN(new_n246_));
  INV_X1    g045(.A(new_n212_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n230_), .A2(new_n237_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n248_), .B2(KEYINPUT29), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n242_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n244_), .A2(new_n246_), .A3(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n252_));
  NOR3_X1   g051(.A1(new_n248_), .A2(KEYINPUT29), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G22gat), .B(G50gat), .Z(new_n255_));
  OAI21_X1  g054(.A(new_n252_), .B1(new_n248_), .B2(KEYINPUT29), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n255_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n256_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(new_n253_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n251_), .A2(new_n257_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n245_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n262_), .B1(new_n244_), .B2(new_n250_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT96), .B1(new_n261_), .B2(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n260_), .A2(new_n257_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT96), .ZN(new_n266_));
  INV_X1    g065(.A(new_n250_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n249_), .A2(new_n242_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n245_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n265_), .A2(new_n266_), .A3(new_n269_), .A4(new_n251_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n246_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n271_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n251_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n265_), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n264_), .A2(new_n270_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT19), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT97), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT98), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n280_), .A2(KEYINPUT98), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT22), .B(G169gat), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n281_), .A2(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT23), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(G183gat), .A3(G190gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT84), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n287_), .B1(G183gat), .B2(G190gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n293_), .A2(KEYINPUT99), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(KEYINPUT99), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n286_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n288_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n297_), .A2(new_n290_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G190gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT25), .B(G183gat), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NOR3_X1   g100(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n302_), .B1(new_n304_), .B2(new_n280_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n212_), .B1(new_n296_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT20), .ZN(new_n308_));
  NOR2_X1   g107(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(G169gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(new_n298_), .B2(new_n292_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT83), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT26), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n312_), .B1(new_n313_), .B2(G190gat), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n300_), .B(new_n314_), .C1(new_n299_), .C2(new_n312_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n305_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n311_), .B1(new_n291_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n308_), .B1(new_n247_), .B2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n279_), .B1(new_n307_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT20), .B1(new_n247_), .B2(new_n318_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n296_), .A2(new_n306_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(new_n323_), .B2(new_n247_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n277_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT18), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  NAND3_X1  g129(.A1(new_n321_), .A2(new_n326_), .A3(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n331_), .A2(KEYINPUT27), .ZN(new_n332_));
  INV_X1    g131(.A(new_n330_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n324_), .A2(new_n325_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n307_), .A2(new_n279_), .A3(new_n319_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  AOI211_X1 g135(.A(new_n277_), .B(new_n322_), .C1(new_n323_), .C2(new_n247_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n333_), .B1(new_n337_), .B2(new_n320_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n331_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT27), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n332_), .A2(new_n336_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G71gat), .B(G99gat), .ZN(new_n342_));
  INV_X1    g141(.A(G43gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT31), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(G15gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n317_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G127gat), .B(G134gat), .Z(new_n352_));
  XOR2_X1   g151(.A(G113gat), .B(G120gat), .Z(new_n353_));
  XOR2_X1   g152(.A(new_n352_), .B(new_n353_), .Z(new_n354_));
  XOR2_X1   g153(.A(new_n354_), .B(KEYINPUT86), .Z(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n351_), .A2(new_n355_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n346_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n358_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(new_n345_), .A3(new_n356_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(KEYINPUT4), .B1(new_n248_), .B2(new_n355_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n354_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n230_), .A2(new_n364_), .A3(new_n237_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n355_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n365_), .B1(new_n238_), .B2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n363_), .B1(new_n367_), .B2(KEYINPUT4), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n369_), .B(KEYINPUT100), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n370_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G1gat), .B(G29gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G57gat), .B(G85gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  NAND2_X1  g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n371_), .A2(new_n381_), .A3(new_n373_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n362_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n275_), .A2(new_n341_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT105), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT102), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n367_), .A2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(KEYINPUT102), .B(new_n365_), .C1(new_n238_), .C2(new_n366_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n370_), .A3(new_n389_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n390_), .B(new_n381_), .C1(new_n370_), .C2(new_n368_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(new_n331_), .A3(new_n338_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT33), .B1(new_n374_), .B2(new_n379_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT33), .ZN(new_n394_));
  AOI211_X1 g193(.A(new_n394_), .B(new_n381_), .C1(new_n371_), .C2(new_n373_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n392_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n371_), .A2(new_n381_), .A3(new_n373_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n381_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n330_), .A2(KEYINPUT32), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n321_), .A2(new_n326_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT103), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT103), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n321_), .A2(new_n326_), .A3(new_n403_), .A4(new_n400_), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT32), .B(new_n330_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n399_), .A2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n275_), .B1(new_n396_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT104), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n275_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(new_n399_), .A3(new_n341_), .ZN(new_n412_));
  OAI211_X1 g211(.A(KEYINPUT104), .B(new_n275_), .C1(new_n396_), .C2(new_n407_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n362_), .B(KEYINPUT87), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n386_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G29gat), .B(G36gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT76), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G43gat), .B(G50gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n418_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G1gat), .B(G8gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G15gat), .B(G22gat), .ZN(new_n423_));
  INV_X1    g222(.A(G1gat), .ZN(new_n424_));
  INV_X1    g223(.A(G8gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT14), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n423_), .B1(new_n426_), .B2(KEYINPUT79), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n426_), .A2(KEYINPUT79), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n422_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  OR3_X1    g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n422_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n421_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT81), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n418_), .B(new_n419_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n429_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT81), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n433_), .A2(new_n437_), .B1(new_n435_), .B2(new_n434_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G229gat), .A2(G233gat), .ZN(new_n439_));
  OR2_X1    g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(KEYINPUT82), .Z(new_n441_));
  NAND2_X1  g240(.A1(new_n434_), .A2(KEYINPUT15), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT15), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n421_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n444_), .A3(new_n435_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n431_), .A2(new_n432_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n436_), .A2(KEYINPUT81), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n441_), .B(new_n445_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n440_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G113gat), .B(G141gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G169gat), .B(G197gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n450_), .B(new_n451_), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n449_), .B(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(G230gat), .A2(G233gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT64), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(G99gat), .B2(G106gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G99gat), .A2(G106gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(KEYINPUT6), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n456_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(KEYINPUT6), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n457_), .A2(G99gat), .A3(G106gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(KEYINPUT64), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G85gat), .ZN(new_n466_));
  INV_X1    g265(.A(G92gat), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n466_), .A2(new_n467_), .A3(KEYINPUT9), .ZN(new_n468_));
  XOR2_X1   g267(.A(G85gat), .B(G92gat), .Z(new_n469_));
  AOI21_X1  g268(.A(new_n468_), .B1(new_n469_), .B2(KEYINPUT9), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT10), .B(G99gat), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n465_), .B(new_n470_), .C1(G106gat), .C2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT8), .ZN(new_n473_));
  INV_X1    g272(.A(G99gat), .ZN(new_n474_));
  INV_X1    g273(.A(G106gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT65), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n474_), .B(new_n475_), .C1(new_n476_), .C2(KEYINPUT7), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n478_), .B(KEYINPUT65), .C1(G99gat), .C2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT67), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n477_), .A2(new_n479_), .A3(KEYINPUT67), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT66), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n462_), .A2(new_n463_), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT66), .B1(new_n458_), .B2(new_n460_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n482_), .A2(new_n483_), .A3(new_n485_), .A4(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n473_), .B1(new_n487_), .B2(new_n469_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n469_), .A2(new_n473_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(new_n465_), .B2(new_n480_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n472_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT68), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G57gat), .B(G64gat), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G71gat), .B(G78gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(KEYINPUT11), .B2(new_n494_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n496_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT68), .B(new_n472_), .C1(new_n488_), .C2(new_n490_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n493_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT69), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT69), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n493_), .A2(new_n504_), .A3(new_n500_), .A4(new_n501_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(KEYINPUT70), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n500_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n469_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n486_), .A2(new_n485_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n477_), .A2(new_n479_), .A3(KEYINPUT67), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT67), .B1(new_n477_), .B2(new_n479_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n508_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n465_), .A2(new_n480_), .ZN(new_n514_));
  OAI22_X1  g313(.A1(new_n513_), .A2(new_n473_), .B1(new_n514_), .B2(new_n489_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT68), .B1(new_n515_), .B2(new_n472_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n501_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n507_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n506_), .A2(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT70), .B1(new_n503_), .B2(new_n505_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n455_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n491_), .A2(KEYINPUT12), .A3(new_n507_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n516_), .A2(new_n517_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n455_), .B1(new_n523_), .B2(new_n500_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT72), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n518_), .B2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n500_), .B1(new_n493_), .B2(new_n501_), .ZN(new_n529_));
  NOR3_X1   g328(.A1(new_n529_), .A2(KEYINPUT72), .A3(new_n526_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n522_), .B(new_n524_), .C1(new_n528_), .C2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT74), .ZN(new_n533_));
  XOR2_X1   g332(.A(KEYINPUT73), .B(KEYINPUT5), .Z(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G120gat), .B(G148gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n521_), .A2(new_n531_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n521_), .B2(new_n531_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT13), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT13), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT37), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT35), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(KEYINPUT77), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT77), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n523_), .A2(new_n421_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n442_), .A2(new_n444_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n558_), .A2(new_n491_), .B1(new_n551_), .B2(new_n550_), .ZN(new_n559_));
  AOI211_X1 g358(.A(new_n554_), .B(new_n556_), .C1(new_n557_), .C2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n557_), .A2(new_n555_), .A3(new_n559_), .A4(new_n552_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G134gat), .B(G162gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT36), .Z(new_n566_));
  NAND3_X1  g365(.A1(new_n561_), .A2(new_n562_), .A3(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n565_), .A2(KEYINPUT36), .ZN(new_n568_));
  INV_X1    g367(.A(new_n562_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n568_), .B1(new_n560_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n547_), .B1(new_n571_), .B2(KEYINPUT78), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT16), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n435_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(new_n500_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT80), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n576_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT17), .B1(new_n579_), .B2(new_n576_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(KEYINPUT17), .B(new_n576_), .C1(new_n579_), .C2(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT78), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n567_), .A2(new_n586_), .A3(KEYINPUT37), .A4(new_n570_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n572_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR4_X1   g388(.A1(new_n416_), .A2(new_n454_), .A3(new_n546_), .A4(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n399_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n424_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT38), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n571_), .B(KEYINPUT106), .Z(new_n595_));
  NOR2_X1   g394(.A1(new_n416_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n585_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n546_), .A2(new_n454_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(G1gat), .B1(new_n599_), .B2(new_n399_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n592_), .A2(new_n593_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n594_), .A2(new_n600_), .A3(new_n601_), .ZN(G1324gat));
  INV_X1    g401(.A(new_n341_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n590_), .A2(new_n425_), .A3(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G8gat), .B1(new_n599_), .B2(new_n341_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n605_), .A2(KEYINPUT39), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(KEYINPUT39), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n604_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g408(.A(G15gat), .B1(new_n599_), .B2(new_n415_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT41), .Z(new_n611_));
  INV_X1    g410(.A(G15gat), .ZN(new_n612_));
  INV_X1    g411(.A(new_n415_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n590_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(G1326gat));
  OAI21_X1  g414(.A(G22gat), .B1(new_n599_), .B2(new_n275_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT42), .ZN(new_n617_));
  INV_X1    g416(.A(G22gat), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n590_), .A2(new_n618_), .A3(new_n411_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(G1327gat));
  NOR2_X1   g419(.A1(new_n416_), .A2(new_n454_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n546_), .A2(new_n585_), .A3(new_n571_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(G29gat), .B1(new_n623_), .B2(new_n591_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT43), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n572_), .A2(new_n587_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n413_), .A2(new_n412_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n398_), .A2(KEYINPUT33), .ZN(new_n628_));
  INV_X1    g427(.A(new_n339_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n391_), .ZN(new_n630_));
  OAI22_X1  g429(.A1(new_n630_), .A2(new_n393_), .B1(new_n399_), .B2(new_n406_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT104), .B1(new_n631_), .B2(new_n275_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n415_), .B1(new_n627_), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n384_), .B(KEYINPUT105), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n626_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT107), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n625_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(KEYINPUT107), .B(KEYINPUT43), .C1(new_n416_), .C2(new_n626_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n546_), .A2(new_n454_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n597_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT44), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644_));
  AOI211_X1 g443(.A(new_n644_), .B(new_n641_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n591_), .A2(G29gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n624_), .B1(new_n646_), .B2(new_n647_), .ZN(G1328gat));
  NAND2_X1  g447(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT109), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT46), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(G36gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n646_), .B2(new_n603_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n341_), .A2(G36gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n621_), .A2(new_n622_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT108), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT108), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n621_), .A2(new_n658_), .A3(new_n622_), .A4(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT45), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n649_), .B(new_n652_), .C1(new_n654_), .C2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n643_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n639_), .A2(KEYINPUT44), .A3(new_n642_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n603_), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G36gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n660_), .B(KEYINPUT45), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n650_), .A4(new_n651_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n663_), .A2(new_n669_), .ZN(G1329gat));
  AOI21_X1  g469(.A(G43gat), .B1(new_n623_), .B2(new_n613_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n362_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(new_n343_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n671_), .B1(new_n646_), .B2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g474(.A(G50gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n623_), .A2(new_n676_), .A3(new_n411_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n646_), .A2(KEYINPUT110), .A3(new_n411_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G50gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT110), .B1(new_n646_), .B2(new_n411_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n677_), .B1(new_n679_), .B2(new_n680_), .ZN(G1331gat));
  NAND2_X1  g480(.A1(new_n633_), .A2(new_n634_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n546_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n453_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(new_n589_), .ZN(new_n686_));
  INV_X1    g485(.A(G57gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n591_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n596_), .A2(new_n585_), .A3(new_n684_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(new_n591_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n688_), .B1(new_n690_), .B2(new_n687_), .ZN(G1332gat));
  INV_X1    g490(.A(G64gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n689_), .B2(new_n603_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT48), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n686_), .A2(new_n692_), .A3(new_n603_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1333gat));
  INV_X1    g495(.A(G71gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n689_), .B2(new_n613_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT49), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n686_), .A2(new_n697_), .A3(new_n613_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1334gat));
  INV_X1    g500(.A(G78gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n689_), .B2(new_n411_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT50), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n686_), .A2(new_n702_), .A3(new_n411_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1335gat));
  INV_X1    g505(.A(new_n639_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n684_), .A2(new_n597_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G85gat), .B1(new_n710_), .B2(new_n399_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n685_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n571_), .A2(new_n585_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n466_), .A3(new_n591_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n711_), .A2(new_n716_), .ZN(G1336gat));
  OAI21_X1  g516(.A(G92gat), .B1(new_n710_), .B2(new_n341_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n715_), .A2(new_n467_), .A3(new_n603_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1337gat));
  NOR3_X1   g519(.A1(new_n714_), .A2(new_n672_), .A3(new_n471_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n709_), .A2(new_n613_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(G99gat), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(G1338gat));
  NAND4_X1  g524(.A1(new_n712_), .A2(new_n475_), .A3(new_n411_), .A4(new_n713_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT112), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n728_));
  INV_X1    g527(.A(new_n708_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n639_), .A2(new_n411_), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n730_), .B2(G106gat), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(G106gat), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT114), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n730_), .A2(new_n728_), .A3(G106gat), .ZN(new_n736_));
  INV_X1    g535(.A(new_n732_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n735_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n733_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT53), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT53), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n733_), .A2(new_n738_), .A3(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1339gat));
  NAND3_X1  g542(.A1(new_n518_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT72), .B1(new_n529_), .B2(new_n526_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n503_), .A2(new_n505_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n522_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n455_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n531_), .A2(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n746_), .A2(KEYINPUT55), .A3(new_n522_), .A4(new_n524_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n749_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n537_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT56), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(new_n756_), .A3(new_n537_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n448_), .B(new_n452_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n441_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n759_), .B(new_n445_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n452_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n760_), .B(new_n761_), .C1(new_n438_), .C2(new_n759_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n758_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT116), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT116), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n758_), .A2(new_n762_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n539_), .A2(new_n767_), .A3(KEYINPUT118), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT118), .B1(new_n539_), .B2(new_n767_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n755_), .B(new_n757_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT58), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT119), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n626_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n755_), .A2(new_n757_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT119), .ZN(new_n776_));
  INV_X1    g575(.A(new_n770_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n768_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n775_), .A2(new_n776_), .A3(KEYINPUT58), .A4(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n773_), .A2(new_n774_), .A3(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n781_));
  INV_X1    g580(.A(new_n767_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n542_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n453_), .A2(new_n539_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n754_), .A2(KEYINPUT115), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(new_n756_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n753_), .B2(new_n537_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT56), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n783_), .B1(new_n786_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n571_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n781_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n781_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n453_), .B(new_n539_), .C1(new_n788_), .C2(KEYINPUT56), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n785_), .A2(new_n756_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n571_), .B(new_n793_), .C1(new_n796_), .C2(new_n783_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n780_), .A2(new_n792_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n597_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n588_), .A2(new_n454_), .A3(new_n545_), .A4(new_n543_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n799_), .A2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n275_), .A2(new_n591_), .A3(new_n341_), .A4(new_n362_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT120), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(KEYINPUT59), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT59), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n802_), .B1(new_n798_), .B2(new_n597_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n806_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n807_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n453_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n809_), .A2(new_n810_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n454_), .A2(G113gat), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n813_), .A2(G113gat), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT121), .ZN(G1340gat));
  INV_X1    g616(.A(G120gat), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n683_), .B2(KEYINPUT60), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n814_), .B(new_n819_), .C1(KEYINPUT60), .C2(new_n818_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n683_), .B1(new_n807_), .B2(new_n811_), .ZN(new_n821_));
  OAI21_X1  g620(.A(G120gat), .B1(new_n821_), .B2(KEYINPUT122), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT122), .ZN(new_n823_));
  AOI211_X1 g622(.A(new_n823_), .B(new_n683_), .C1(new_n807_), .C2(new_n811_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n820_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT123), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT123), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n827_), .B(new_n820_), .C1(new_n822_), .C2(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1341gat));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n814_), .A2(new_n830_), .A3(new_n585_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n597_), .B1(new_n807_), .B2(new_n811_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n830_), .ZN(G1342gat));
  INV_X1    g632(.A(G134gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n814_), .A2(new_n834_), .A3(new_n595_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n626_), .B1(new_n807_), .B2(new_n811_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n834_), .ZN(G1343gat));
  INV_X1    g636(.A(KEYINPUT124), .ZN(new_n838_));
  NOR4_X1   g637(.A1(new_n613_), .A2(new_n603_), .A3(new_n275_), .A4(new_n399_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n804_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n804_), .B2(new_n839_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n454_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(new_n223_), .ZN(G1344gat));
  NOR2_X1   g643(.A1(new_n842_), .A2(new_n683_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(new_n224_), .ZN(G1345gat));
  INV_X1    g645(.A(new_n842_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n585_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT61), .B(G155gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1346gat));
  OAI21_X1  g649(.A(G162gat), .B1(new_n842_), .B2(new_n626_), .ZN(new_n851_));
  INV_X1    g650(.A(G162gat), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n595_), .A2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n851_), .B1(new_n842_), .B2(new_n853_), .ZN(G1347gat));
  NOR2_X1   g653(.A1(new_n809_), .A2(new_n591_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n411_), .A2(new_n415_), .A3(new_n341_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n857_), .A2(new_n453_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT62), .ZN(new_n859_));
  INV_X1    g658(.A(G169gat), .ZN(new_n860_));
  OR3_X1    g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n859_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n858_), .A2(new_n283_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(G1348gat));
  NAND2_X1  g663(.A1(new_n857_), .A2(new_n546_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g665(.A1(new_n857_), .A2(new_n585_), .ZN(new_n867_));
  MUX2_X1   g666(.A(new_n300_), .B(G183gat), .S(new_n867_), .Z(G1350gat));
  NAND3_X1  g667(.A1(new_n857_), .A2(new_n299_), .A3(new_n595_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n626_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n857_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(G190gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n869_), .B1(new_n871_), .B2(new_n872_), .ZN(G1351gat));
  AND4_X1   g672(.A1(new_n415_), .A2(new_n855_), .A3(new_n411_), .A4(new_n603_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n453_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g675(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT125), .B(G204gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n874_), .A2(new_n546_), .ZN(new_n879_));
  MUX2_X1   g678(.A(new_n877_), .B(new_n878_), .S(new_n879_), .Z(G1353gat));
  NOR2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT126), .ZN(new_n882_));
  NAND2_X1  g681(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n874_), .A2(new_n585_), .A3(new_n882_), .A4(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n881_), .A2(KEYINPUT126), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1354gat));
  AOI21_X1  g685(.A(G218gat), .B1(new_n874_), .B2(new_n595_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n870_), .A2(G218gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT127), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n887_), .B1(new_n874_), .B2(new_n889_), .ZN(G1355gat));
endmodule


