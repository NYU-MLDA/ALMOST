//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n939_, new_n941_, new_n942_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n985_, new_n986_, new_n987_, new_n989_, new_n990_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n998_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1007_, new_n1008_;
  INV_X1    g000(.A(KEYINPUT104), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G134gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G127gat), .ZN(new_n206_));
  INV_X1    g005(.A(G127gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G134gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(KEYINPUT85), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n206_), .A2(new_n208_), .A3(KEYINPUT85), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G113gat), .B(G120gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n212_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n211_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n214_), .B1(new_n215_), .B2(new_n209_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT87), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G141gat), .ZN(new_n222_));
  INV_X1    g021(.A(G148gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AND2_X1   g023(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n221_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n219_), .A2(new_n220_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n226_), .A2(new_n227_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n233_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT86), .B1(new_n232_), .B2(new_n236_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G155gat), .A2(G162gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT86), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(KEYINPUT1), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n238_), .A3(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G141gat), .B(G148gat), .Z(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n235_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n218_), .A2(new_n245_), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n231_), .A2(new_n234_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n217_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(KEYINPUT4), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n218_), .A2(new_n245_), .A3(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n251_), .A2(KEYINPUT97), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(KEYINPUT97), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n204_), .B(new_n249_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n246_), .A2(new_n248_), .A3(new_n203_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G1gat), .B(G29gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(G85gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT0), .B(G57gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n260_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n254_), .A2(new_n255_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(KEYINPUT102), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT102), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n256_), .A2(new_n265_), .A3(new_n260_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G64gat), .B(G92gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT96), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G8gat), .B(G36gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT24), .ZN(new_n275_));
  INV_X1    g074(.A(G169gat), .ZN(new_n276_));
  INV_X1    g075(.A(G176gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n278_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT25), .B(G183gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G190gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT83), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(KEYINPUT83), .A2(G183gat), .A3(G190gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(KEYINPUT23), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT82), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n290_), .A2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT23), .B1(new_n288_), .B2(new_n289_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n294_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n298_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT22), .B(G169gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n280_), .B1(new_n302_), .B2(new_n277_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n285_), .A2(new_n297_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT90), .ZN(new_n305_));
  INV_X1    g104(.A(G197gat), .ZN(new_n306_));
  INV_X1    g105(.A(G204gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G197gat), .A2(G204gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n305_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G218gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(G211gat), .ZN(new_n312_));
  INV_X1    g111(.A(G211gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(G218gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n312_), .A2(new_n314_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT21), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(G197gat), .A2(G204gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G197gat), .A2(G204gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT90), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G211gat), .B(G218gat), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT21), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n274_), .B1(new_n304_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT84), .ZN(new_n327_));
  AOI21_X1  g126(.A(G176gat), .B1(new_n327_), .B2(KEYINPUT22), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(new_n276_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n280_), .A2(new_n281_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT25), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n332_), .B1(new_n333_), .B2(G183gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n284_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G183gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT25), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(G183gat), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n332_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(KEYINPUT81), .B(new_n331_), .C1(new_n335_), .C2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n278_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n289_), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT83), .B1(G183gat), .B2(G190gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n292_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n295_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n286_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n341_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n340_), .A2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n331_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n330_), .B1(new_n349_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT91), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n318_), .A2(new_n354_), .A3(new_n324_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT21), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n321_), .A2(new_n322_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n308_), .A2(new_n309_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n315_), .A2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n356_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT91), .B1(new_n360_), .B2(new_n323_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n326_), .B1(new_n353_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G226gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT19), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT20), .B1(new_n304_), .B2(new_n325_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n367_), .B1(new_n362_), .B2(new_n353_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n365_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n366_), .A2(KEYINPUT101), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n329_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n297_), .A2(new_n298_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n340_), .A2(new_n348_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n284_), .B(new_n334_), .C1(new_n283_), .C2(new_n332_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT81), .B1(new_n375_), .B2(new_n331_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n373_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(new_n355_), .A3(new_n361_), .ZN(new_n378_));
  AOI211_X1 g177(.A(KEYINPUT101), .B(new_n369_), .C1(new_n378_), .C2(new_n326_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n273_), .B1(new_n370_), .B2(new_n380_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n326_), .B(new_n369_), .C1(new_n353_), .C2(new_n362_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT94), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n377_), .B1(new_n355_), .B2(new_n361_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n365_), .B1(new_n384_), .B2(new_n367_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT94), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n378_), .A2(new_n386_), .A3(new_n369_), .A4(new_n326_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n383_), .A2(new_n385_), .A3(new_n273_), .A4(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT27), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT103), .B1(new_n381_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT27), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n352_), .A2(new_n340_), .A3(new_n348_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n354_), .B1(new_n318_), .B2(new_n324_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n360_), .A2(KEYINPUT91), .A3(new_n323_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n392_), .B(new_n373_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n285_), .A2(new_n297_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n301_), .A2(new_n303_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n357_), .A2(new_n359_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n323_), .B1(new_n399_), .B2(KEYINPUT21), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n274_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n369_), .B1(new_n395_), .B2(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n378_), .A2(new_n369_), .A3(new_n326_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n402_), .B1(new_n403_), .B2(new_n386_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n273_), .B1(new_n404_), .B2(new_n383_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n388_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n391_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n273_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n395_), .A2(new_n369_), .A3(new_n401_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n369_), .B1(new_n378_), .B2(new_n326_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT101), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n408_), .B1(new_n412_), .B2(new_n379_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT103), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(KEYINPUT27), .A4(new_n388_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n390_), .A2(new_n407_), .A3(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G22gat), .B(G50gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G78gat), .B(G106gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n417_), .B(new_n418_), .Z(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT29), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n235_), .B2(new_n244_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G228gat), .A2(G233gat), .ZN(new_n423_));
  XOR2_X1   g222(.A(new_n423_), .B(KEYINPUT89), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(new_n355_), .A3(new_n361_), .ZN(new_n427_));
  OAI211_X1 g226(.A(KEYINPUT92), .B(new_n425_), .C1(new_n422_), .C2(new_n325_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n400_), .B1(new_n247_), .B2(new_n421_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT92), .B1(new_n430_), .B2(new_n425_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n427_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT93), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT93), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n434_), .B(new_n427_), .C1(new_n429_), .C2(new_n431_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n247_), .A2(new_n421_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n433_), .A2(new_n435_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n439_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n420_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n435_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n425_), .B1(new_n422_), .B2(new_n325_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT92), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n428_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n434_), .B1(new_n447_), .B2(new_n427_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n438_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n433_), .A2(new_n435_), .A3(new_n439_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n419_), .A3(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(G43gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n377_), .B(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n454_), .A2(new_n217_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n217_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G227gat), .A2(G233gat), .ZN(new_n457_));
  INV_X1    g256(.A(G15gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT30), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT31), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OR3_X1    g261(.A1(new_n455_), .A2(new_n456_), .A3(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n462_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n442_), .A2(new_n451_), .A3(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n465_), .B1(new_n442_), .B2(new_n451_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n267_), .B(new_n416_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n273_), .A2(KEYINPUT32), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n412_), .B2(new_n379_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n404_), .A2(new_n383_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n470_), .B1(new_n471_), .B2(new_n469_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n408_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n388_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n203_), .B(new_n249_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT100), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n251_), .B(KEYINPUT97), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT100), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(new_n203_), .A4(new_n249_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n246_), .A2(new_n248_), .A3(new_n204_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n480_), .A2(KEYINPUT99), .A3(new_n260_), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT99), .B1(new_n480_), .B2(new_n260_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n476_), .A2(new_n479_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT98), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n485_), .A2(KEYINPUT33), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n263_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n254_), .A2(new_n255_), .A3(new_n262_), .A4(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n490_));
  OAI22_X1  g289(.A1(new_n267_), .A2(new_n472_), .B1(new_n474_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n442_), .A2(new_n451_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n465_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n468_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G113gat), .B(G141gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G169gat), .B(G197gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n495_), .B(new_n496_), .Z(new_n497_));
  XNOR2_X1  g296(.A(G29gat), .B(G36gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT70), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G43gat), .B(G50gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT70), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n498_), .B(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(new_n500_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT14), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT74), .B(G1gat), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n507_), .B1(new_n508_), .B2(G8gat), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT75), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G1gat), .B(G8gat), .Z(new_n514_));
  AND2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n513_), .A2(new_n514_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n506_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n513_), .A2(new_n514_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n506_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n513_), .A2(new_n514_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT15), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n526_), .B1(new_n502_), .B2(new_n505_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n504_), .A2(new_n500_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n499_), .A2(new_n501_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(KEYINPUT15), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n518_), .A2(new_n531_), .A3(new_n520_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n517_), .A2(new_n532_), .A3(new_n523_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n525_), .A2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n497_), .B1(new_n534_), .B2(KEYINPUT78), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT78), .ZN(new_n536_));
  INV_X1    g335(.A(new_n497_), .ZN(new_n537_));
  AOI211_X1 g336(.A(new_n536_), .B(new_n537_), .C1(new_n525_), .C2(new_n533_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n535_), .A2(new_n538_), .A3(KEYINPUT79), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT79), .ZN(new_n540_));
  INV_X1    g339(.A(new_n533_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n523_), .B1(new_n517_), .B2(new_n521_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT78), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n537_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n534_), .A2(KEYINPUT78), .A3(new_n497_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n540_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n539_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n202_), .B1(new_n494_), .B2(new_n548_), .ZN(new_n549_));
  AOI211_X1 g348(.A(KEYINPUT104), .B(new_n547_), .C1(new_n468_), .C2(new_n493_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n518_), .A2(new_n520_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n554_));
  XOR2_X1   g353(.A(G71gat), .B(G78gat), .Z(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n554_), .A2(new_n555_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n556_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT76), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n560_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n552_), .B(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G127gat), .B(G155gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G183gat), .B(G211gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n564_), .A2(KEYINPUT17), .A3(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(KEYINPUT17), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n564_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT64), .ZN(new_n575_));
  OAI211_X1 g374(.A(G85gat), .B(G92gat), .C1(new_n575_), .C2(KEYINPUT9), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT65), .ZN(new_n577_));
  AND2_X1   g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT65), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n578_), .B(new_n579_), .C1(new_n575_), .C2(KEYINPUT9), .ZN(new_n580_));
  NOR2_X1   g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT9), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n581_), .A2(KEYINPUT64), .A3(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n577_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n585_));
  NOR2_X1   g384(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(G106gat), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT6), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT6), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(G99gat), .A3(G106gat), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n587_), .A2(new_n588_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n584_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n583_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT66), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n577_), .A2(new_n580_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n583_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT66), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n599_), .A2(new_n600_), .A3(new_n584_), .A4(new_n593_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n578_), .A2(new_n581_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(KEYINPUT8), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n590_), .A2(new_n592_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT7), .ZN(new_n606_));
  INV_X1    g405(.A(G99gat), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(new_n607_), .A3(new_n588_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n604_), .B1(new_n605_), .B2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT67), .B1(new_n590_), .B2(new_n592_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(new_n610_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n590_), .A2(new_n592_), .A3(KEYINPUT67), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n603_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT8), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n611_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n602_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n560_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n560_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n602_), .A2(new_n618_), .A3(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(KEYINPUT12), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n621_), .B1(new_n602_), .B2(new_n618_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT12), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT68), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT68), .ZN(new_n630_));
  INV_X1    g429(.A(new_n628_), .ZN(new_n631_));
  AOI211_X1 g430(.A(new_n630_), .B(new_n631_), .C1(new_n623_), .C2(new_n626_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n602_), .A2(new_n618_), .A3(new_n621_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n631_), .B1(new_n634_), .B2(new_n624_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT5), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n637_), .B(new_n638_), .Z(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n633_), .A2(new_n635_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n639_), .B(KEYINPUT69), .Z(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT13), .B1(new_n642_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n645_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT13), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(new_n648_), .A3(new_n641_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT37), .ZN(new_n652_));
  NAND2_X1  g451(.A1(G232gat), .A2(G233gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT34), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(KEYINPUT35), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n531_), .B2(new_n619_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT71), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n614_), .A2(new_n612_), .A3(new_n610_), .ZN(new_n658_));
  OAI21_X1  g457(.A(KEYINPUT8), .B1(new_n658_), .B2(new_n603_), .ZN(new_n659_));
  AOI22_X1  g458(.A1(new_n596_), .A2(new_n601_), .B1(new_n659_), .B2(new_n611_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n657_), .B1(new_n660_), .B2(new_n506_), .ZN(new_n661_));
  AND4_X1   g460(.A1(new_n657_), .A2(new_n602_), .A3(new_n618_), .A4(new_n506_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n656_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n654_), .A2(KEYINPUT35), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n656_), .B(new_n664_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(KEYINPUT73), .A3(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(G190gat), .B(G218gat), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT72), .ZN(new_n670_));
  XOR2_X1   g469(.A(G134gat), .B(G162gat), .Z(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(KEYINPUT36), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n668_), .A2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n666_), .A2(KEYINPUT73), .A3(new_n667_), .A4(new_n674_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n673_), .A2(KEYINPUT36), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n652_), .B1(new_n678_), .B2(new_n681_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT37), .B(new_n680_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NOR4_X1   g484(.A1(new_n551_), .A2(new_n574_), .A3(new_n651_), .A4(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n267_), .B(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(new_n508_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT38), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n680_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n494_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT106), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n535_), .A2(new_n538_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n651_), .A2(new_n574_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n694_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n694_), .A2(KEYINPUT107), .A3(new_n697_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n267_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(G1gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n691_), .B1(new_n702_), .B2(new_n703_), .ZN(G1324gat));
  INV_X1    g503(.A(new_n416_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n694_), .A2(new_n705_), .A3(new_n697_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G8gat), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(KEYINPUT108), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT39), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n706_), .B2(G8gat), .ZN(new_n711_));
  OR3_X1    g510(.A1(new_n708_), .A2(new_n709_), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n709_), .ZN(new_n713_));
  INV_X1    g512(.A(G8gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n686_), .A2(new_n714_), .A3(new_n705_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n712_), .A2(KEYINPUT40), .A3(new_n713_), .A4(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT40), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n708_), .A2(new_n711_), .A3(new_n709_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n713_), .A2(new_n715_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n716_), .A2(new_n720_), .ZN(G1325gat));
  INV_X1    g520(.A(new_n465_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n686_), .A2(new_n458_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n700_), .A2(new_n701_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n458_), .B1(new_n724_), .B2(new_n722_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(KEYINPUT41), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(KEYINPUT41), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(G1326gat));
  INV_X1    g527(.A(G22gat), .ZN(new_n729_));
  INV_X1    g528(.A(new_n492_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n686_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n492_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n732_), .A2(new_n729_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n732_), .A2(KEYINPUT42), .A3(new_n729_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n731_), .B1(new_n735_), .B2(new_n736_), .ZN(G1327gat));
  NOR2_X1   g536(.A1(new_n692_), .A2(new_n573_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n738_), .A2(KEYINPUT110), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(KEYINPUT110), .ZN(new_n740_));
  AOI22_X1  g539(.A1(new_n739_), .A2(new_n740_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n741_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n741_), .B(KEYINPUT111), .C1(new_n549_), .C2(new_n550_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n267_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G29gat), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n650_), .A2(new_n574_), .A3(new_n695_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(KEYINPUT109), .B1(new_n682_), .B2(new_n683_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT43), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n752_), .A2(new_n685_), .A3(new_n494_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n684_), .B1(new_n468_), .B2(new_n493_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n754_), .A2(new_n752_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n750_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n494_), .A2(new_n685_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(KEYINPUT43), .A3(new_n751_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n754_), .A2(new_n752_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT44), .B1(new_n762_), .B2(new_n750_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n758_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n688_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n765_), .A2(G29gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n748_), .B1(new_n764_), .B2(new_n766_), .ZN(G1328gat));
  NOR2_X1   g566(.A1(KEYINPUT114), .A2(KEYINPUT46), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n416_), .A2(G36gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n744_), .A2(new_n745_), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT113), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n744_), .A2(new_n772_), .A3(new_n745_), .A4(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n771_), .A2(KEYINPUT45), .A3(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n756_), .A2(new_n757_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n762_), .A2(KEYINPUT44), .A3(new_n750_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n705_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n781_), .A2(KEYINPUT112), .A3(G36gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT112), .B1(new_n781_), .B2(G36gat), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n768_), .B1(new_n778_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n781_), .A2(G36gat), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n781_), .A2(KEYINPUT112), .A3(G36gat), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n768_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n776_), .A4(new_n777_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n785_), .A2(new_n792_), .ZN(G1329gat));
  NAND3_X1  g592(.A1(new_n764_), .A2(G43gat), .A3(new_n722_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n746_), .A2(new_n722_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(G43gat), .ZN(new_n796_));
  XOR2_X1   g595(.A(KEYINPUT115), .B(KEYINPUT47), .Z(new_n797_));
  XNOR2_X1  g596(.A(new_n796_), .B(new_n797_), .ZN(G1330gat));
  NOR2_X1   g597(.A1(new_n492_), .A2(G50gat), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT116), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n746_), .A2(new_n800_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n758_), .A2(new_n763_), .A3(new_n492_), .ZN(new_n802_));
  INV_X1    g601(.A(G50gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(G1331gat));
  AND3_X1   g603(.A1(new_n651_), .A2(new_n494_), .A3(new_n696_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n805_), .A2(new_n573_), .A3(new_n684_), .ZN(new_n806_));
  INV_X1    g605(.A(G57gat), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n765_), .ZN(new_n808_));
  AND4_X1   g607(.A1(new_n694_), .A2(new_n573_), .A3(new_n651_), .A4(new_n547_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n809_), .A2(new_n747_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n810_), .B2(new_n807_), .ZN(G1332gat));
  INV_X1    g610(.A(G64gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n809_), .B2(new_n705_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT48), .Z(new_n814_));
  NAND3_X1  g613(.A1(new_n806_), .A2(new_n812_), .A3(new_n705_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(G1333gat));
  INV_X1    g615(.A(G71gat), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(new_n809_), .B2(new_n722_), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(KEYINPUT49), .Z(new_n819_));
  NAND3_X1  g618(.A1(new_n806_), .A2(new_n817_), .A3(new_n722_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1334gat));
  INV_X1    g620(.A(G78gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n809_), .B2(new_n730_), .ZN(new_n823_));
  XOR2_X1   g622(.A(new_n823_), .B(KEYINPUT50), .Z(new_n824_));
  NAND3_X1  g623(.A1(new_n806_), .A2(new_n822_), .A3(new_n730_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1335gat));
  NAND2_X1  g625(.A1(new_n739_), .A2(new_n740_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n805_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(G85gat), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n765_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n650_), .A2(new_n573_), .A3(new_n695_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n762_), .A2(new_n831_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n832_), .A2(new_n747_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n830_), .B1(new_n833_), .B2(new_n829_), .ZN(G1336gat));
  AOI21_X1  g633(.A(G92gat), .B1(new_n828_), .B2(new_n705_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT117), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n705_), .A2(G92gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n832_), .B2(new_n837_), .ZN(G1337gat));
  NAND3_X1  g637(.A1(new_n828_), .A2(new_n587_), .A3(new_n722_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(KEYINPUT118), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n607_), .B1(new_n832_), .B2(new_n722_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1338gat));
  NAND3_X1  g643(.A1(new_n828_), .A2(new_n588_), .A3(new_n730_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n832_), .A2(new_n730_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(G106gat), .ZN(new_n848_));
  AOI211_X1 g647(.A(KEYINPUT52), .B(new_n588_), .C1(new_n832_), .C2(new_n730_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n845_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g650(.A(G113gat), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n765_), .A2(new_n416_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n853_), .A2(new_n730_), .A3(new_n465_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n523_), .B1(new_n552_), .B2(new_n506_), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n532_), .A2(new_n856_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n857_), .A2(new_n497_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n534_), .A2(new_n497_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n642_), .B2(new_n645_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n695_), .A2(new_n641_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT56), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n623_), .A2(new_n631_), .A3(new_n626_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n634_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n626_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n628_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n864_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n633_), .B2(new_n868_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n863_), .B1(new_n870_), .B2(new_n644_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n867_), .A2(new_n630_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n631_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT68), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(new_n868_), .A3(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n864_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(KEYINPUT55), .B2(new_n873_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n644_), .B1(new_n875_), .B2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT56), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n862_), .B1(new_n871_), .B2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n861_), .B1(new_n880_), .B2(KEYINPUT119), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n695_), .A2(new_n641_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n878_), .A2(KEYINPUT56), .ZN(new_n883_));
  AOI211_X1 g682(.A(new_n863_), .B(new_n644_), .C1(new_n875_), .C2(new_n877_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n882_), .B(KEYINPUT119), .C1(new_n883_), .C2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n692_), .B1(new_n881_), .B2(new_n886_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(KEYINPUT121), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(new_n885_), .A3(new_n861_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n692_), .A2(KEYINPUT57), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n860_), .A2(new_n641_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n871_), .B2(new_n879_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n898_), .A2(KEYINPUT58), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n684_), .B1(new_n898_), .B2(KEYINPUT58), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n895_), .A2(new_n896_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n888_), .B1(new_n895_), .B2(new_n692_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n574_), .B1(new_n891_), .B2(new_n904_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n650_), .A2(new_n573_), .A3(new_n547_), .A4(new_n684_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n855_), .B1(new_n905_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n852_), .B1(new_n911_), .B2(new_n696_), .ZN(new_n912_));
  AOI21_X1  g711(.A(KEYINPUT59), .B1(new_n854_), .B2(KEYINPUT122), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n573_), .B1(new_n890_), .B2(new_n901_), .ZN(new_n914_));
  OAI221_X1 g713(.A(new_n913_), .B1(KEYINPUT122), .B2(new_n854_), .C1(new_n914_), .C2(new_n908_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n547_), .A2(new_n852_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n915_), .B(new_n916_), .C1(new_n910_), .C2(new_n917_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n912_), .A2(new_n918_), .ZN(G1340gat));
  XNOR2_X1  g718(.A(KEYINPUT123), .B(G120gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n920_), .B1(new_n650_), .B2(KEYINPUT60), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n910_), .B(new_n921_), .C1(KEYINPUT60), .C2(new_n920_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n915_), .A2(new_n651_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n911_), .B2(KEYINPUT59), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n924_), .B2(new_n920_), .ZN(G1341gat));
  OAI21_X1  g724(.A(new_n207_), .B1(new_n911_), .B2(new_n574_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n574_), .A2(new_n207_), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n915_), .B(new_n927_), .C1(new_n910_), .C2(new_n917_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1342gat));
  OAI21_X1  g728(.A(new_n205_), .B1(new_n911_), .B2(new_n692_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n684_), .A2(new_n205_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n915_), .B(new_n931_), .C1(new_n910_), .C2(new_n917_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1343gat));
  NAND2_X1  g732(.A1(new_n905_), .A2(new_n909_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n765_), .A2(new_n416_), .A3(new_n466_), .ZN(new_n935_));
  XOR2_X1   g734(.A(new_n935_), .B(KEYINPUT124), .Z(new_n936_));
  NAND3_X1  g735(.A1(new_n934_), .A2(new_n695_), .A3(new_n936_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g737(.A1(new_n934_), .A2(new_n651_), .A3(new_n936_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g739(.A1(new_n934_), .A2(new_n573_), .A3(new_n936_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT61), .B(G155gat), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n941_), .B(new_n942_), .ZN(G1346gat));
  INV_X1    g742(.A(G162gat), .ZN(new_n944_));
  INV_X1    g743(.A(new_n692_), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n934_), .A2(new_n944_), .A3(new_n945_), .A4(new_n936_), .ZN(new_n946_));
  AND3_X1   g745(.A1(new_n934_), .A2(new_n685_), .A3(new_n936_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n947_), .B2(new_n944_), .ZN(G1347gat));
  NAND2_X1  g747(.A1(new_n899_), .A2(new_n900_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n896_), .B1(new_n881_), .B2(new_n886_), .ZN(new_n950_));
  INV_X1    g749(.A(new_n861_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n951_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n945_), .B1(new_n952_), .B2(new_n885_), .ZN(new_n953_));
  OAI211_X1 g752(.A(new_n949_), .B(new_n950_), .C1(new_n953_), .C2(new_n888_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n908_), .B1(new_n954_), .B2(new_n574_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n955_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n765_), .A2(new_n416_), .A3(new_n465_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n695_), .A2(new_n302_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  NAND4_X1  g758(.A1(new_n956_), .A2(new_n492_), .A3(new_n957_), .A4(new_n959_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n957_), .A2(new_n962_), .A3(new_n695_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n963_), .A2(new_n492_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n962_), .B1(new_n957_), .B2(new_n695_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  OAI211_X1 g766(.A(new_n961_), .B(G169gat), .C1(new_n955_), .C2(new_n967_), .ZN(new_n968_));
  INV_X1    g767(.A(new_n968_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n966_), .B1(new_n914_), .B2(new_n908_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n961_), .B1(new_n970_), .B2(G169gat), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n960_), .B1(new_n969_), .B2(new_n971_), .ZN(new_n972_));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n972_), .A2(new_n973_), .ZN(new_n974_));
  OAI211_X1 g773(.A(KEYINPUT126), .B(new_n960_), .C1(new_n969_), .C2(new_n971_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n974_), .A2(new_n975_), .ZN(G1348gat));
  OAI211_X1 g775(.A(new_n492_), .B(new_n957_), .C1(new_n914_), .C2(new_n908_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n277_), .B1(new_n977_), .B2(new_n650_), .ZN(new_n978_));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979_));
  OR2_X1    g778(.A1(new_n978_), .A2(new_n979_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n978_), .A2(new_n979_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n730_), .B1(new_n905_), .B2(new_n909_), .ZN(new_n982_));
  AND3_X1   g781(.A1(new_n957_), .A2(G176gat), .A3(new_n651_), .ZN(new_n983_));
  AOI22_X1  g782(.A1(new_n980_), .A2(new_n981_), .B1(new_n982_), .B2(new_n983_), .ZN(G1349gat));
  NAND2_X1  g783(.A1(new_n957_), .A2(new_n573_), .ZN(new_n985_));
  NOR4_X1   g784(.A1(new_n955_), .A2(new_n283_), .A3(new_n730_), .A4(new_n985_), .ZN(new_n986_));
  NAND3_X1  g785(.A1(new_n982_), .A2(new_n573_), .A3(new_n957_), .ZN(new_n987_));
  AOI21_X1  g786(.A(new_n986_), .B1(new_n987_), .B2(new_n336_), .ZN(G1350gat));
  OAI21_X1  g787(.A(G190gat), .B1(new_n977_), .B2(new_n684_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n945_), .A2(new_n284_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n989_), .B1(new_n977_), .B2(new_n990_), .ZN(G1351gat));
  NOR4_X1   g790(.A1(new_n416_), .A2(new_n747_), .A3(new_n492_), .A4(new_n722_), .ZN(new_n992_));
  AND2_X1   g791(.A1(new_n934_), .A2(new_n992_), .ZN(new_n993_));
  AOI21_X1  g792(.A(G197gat), .B1(new_n993_), .B2(new_n695_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n934_), .A2(new_n992_), .ZN(new_n995_));
  NOR3_X1   g794(.A1(new_n995_), .A2(new_n306_), .A3(new_n696_), .ZN(new_n996_));
  NOR2_X1   g795(.A1(new_n994_), .A2(new_n996_), .ZN(G1352gat));
  NAND3_X1  g796(.A1(new_n934_), .A2(new_n651_), .A3(new_n992_), .ZN(new_n998_));
  XNOR2_X1  g797(.A(new_n998_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g798(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1000_));
  INV_X1    g799(.A(new_n1000_), .ZN(new_n1001_));
  AOI21_X1  g800(.A(new_n574_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1002_));
  AOI21_X1  g801(.A(new_n1001_), .B1(new_n993_), .B2(new_n1002_), .ZN(new_n1003_));
  INV_X1    g802(.A(new_n1002_), .ZN(new_n1004_));
  NOR3_X1   g803(.A1(new_n995_), .A2(new_n1000_), .A3(new_n1004_), .ZN(new_n1005_));
  NOR2_X1   g804(.A1(new_n1003_), .A2(new_n1005_), .ZN(G1354gat));
  NAND3_X1  g805(.A1(new_n993_), .A2(new_n311_), .A3(new_n945_), .ZN(new_n1007_));
  OAI21_X1  g806(.A(G218gat), .B1(new_n995_), .B2(new_n684_), .ZN(new_n1008_));
  NAND2_X1  g807(.A1(new_n1007_), .A2(new_n1008_), .ZN(G1355gat));
endmodule


