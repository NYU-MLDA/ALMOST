//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G134gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n203_), .B(G162gat), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT10), .B(G99gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT64), .ZN(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(G85gat), .B(G92gat), .Z(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT9), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT6), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n214_), .B(new_n216_), .C1(KEYINPUT9), .C2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n212_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  OR3_X1    g020(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n216_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n213_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT8), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n224_), .B(KEYINPUT8), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(KEYINPUT66), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n220_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G29gat), .B(G36gat), .ZN(new_n232_));
  INV_X1    g031(.A(G43gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(G50gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT15), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n231_), .A2(KEYINPUT68), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n229_), .A2(KEYINPUT66), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n226_), .A2(new_n227_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n219_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n235_), .B(KEYINPUT15), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n239_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n226_), .A2(new_n219_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n235_), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n238_), .A2(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G232gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT34), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT35), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n249_), .A2(KEYINPUT35), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n247_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n250_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n206_), .B(new_n208_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n238_), .A2(new_n244_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n226_), .A2(new_n219_), .A3(new_n235_), .ZN(new_n256_));
  OAI211_X1 g055(.A(KEYINPUT35), .B(new_n249_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n247_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n207_), .B(KEYINPUT69), .Z(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n254_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n254_), .A2(KEYINPUT70), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n262_), .B1(new_n263_), .B2(KEYINPUT37), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT37), .ZN(new_n265_));
  AOI211_X1 g064(.A(KEYINPUT71), .B(new_n265_), .C1(new_n254_), .C2(KEYINPUT70), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n261_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n207_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n268_), .B1(new_n269_), .B2(new_n206_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT71), .B1(new_n270_), .B2(new_n265_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n263_), .A2(new_n262_), .A3(KEYINPUT37), .ZN(new_n272_));
  INV_X1    g071(.A(new_n261_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n267_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G57gat), .B(G64gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT11), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT65), .B(G71gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G78gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(KEYINPUT11), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n280_), .B1(new_n282_), .B2(new_n279_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n245_), .A2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n283_), .B1(new_n226_), .B2(new_n219_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(G230gat), .A2(G233gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n231_), .A2(KEYINPUT12), .A3(new_n283_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT12), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n285_), .A3(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n289_), .B1(new_n293_), .B2(new_n288_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G120gat), .B(G148gat), .ZN(new_n295_));
  INV_X1    g094(.A(G204gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT5), .ZN(new_n298_));
  INV_X1    g097(.A(G176gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT67), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n294_), .B(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n303_), .A2(KEYINPUT13), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(KEYINPUT13), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G127gat), .B(G155gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G183gat), .B(G211gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT72), .B(G22gat), .ZN(new_n312_));
  INV_X1    g111(.A(G15gat), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G1gat), .ZN(new_n315_));
  INV_X1    g114(.A(G8gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT14), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(new_n313_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n314_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G1gat), .B(G8gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G231gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(new_n283_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n311_), .B1(new_n324_), .B2(KEYINPUT74), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT17), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n324_), .B2(new_n311_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n327_), .B1(new_n329_), .B2(new_n325_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n275_), .A2(new_n306_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G127gat), .B(G134gat), .ZN(new_n334_));
  INV_X1    g133(.A(G113gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G120gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G15gat), .B(G43gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(G183gat), .A3(G190gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT23), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n342_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n344_), .B1(new_n348_), .B2(new_n343_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n349_), .B1(G183gat), .B2(G190gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT22), .B(G169gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n352_), .B1(new_n353_), .B2(new_n299_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT25), .B(G183gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G190gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G169gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n299_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n359_), .A2(KEYINPUT24), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(KEYINPUT24), .A3(new_n351_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n357_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n350_), .A2(new_n354_), .B1(new_n347_), .B2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n340_), .B(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G71gat), .B(G99gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G227gat), .A2(G233gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT30), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n368_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n365_), .B(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n372_), .B(KEYINPUT82), .Z(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT84), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT83), .B1(G141gat), .B2(G148gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT2), .ZN(new_n381_));
  OAI22_X1  g180(.A1(new_n378_), .A2(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383_));
  OAI211_X1 g182(.A(KEYINPUT84), .B(KEYINPUT2), .C1(new_n383_), .C2(KEYINPUT83), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n377_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n385_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT85), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT1), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n383_), .B1(KEYINPUT1), .B2(new_n386_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n392_), .B(new_n393_), .C1(G141gat), .C2(G148gat), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT85), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n385_), .A2(new_n395_), .A3(new_n388_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n390_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n398_));
  OR3_X1    g197(.A1(new_n397_), .A2(KEYINPUT29), .A3(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G22gat), .B(G50gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n398_), .B1(new_n397_), .B2(KEYINPUT29), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n401_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G78gat), .B(G106gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n407_), .B(KEYINPUT92), .Z(new_n408_));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(G211gat), .A2(G218gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(G211gat), .A2(G218gat), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT88), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(G211gat), .ZN(new_n414_));
  INV_X1    g213(.A(G218gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT88), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G211gat), .A2(G218gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n413_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G197gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT87), .B1(new_n421_), .B2(G204gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n296_), .A3(G197gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(G204gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n420_), .A2(KEYINPUT89), .A3(KEYINPUT21), .A4(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT89), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n413_), .A2(new_n419_), .A3(KEYINPUT21), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n422_), .A2(new_n424_), .B1(new_n421_), .B2(G204gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n428_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT21), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n296_), .A2(G197gat), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(new_n426_), .B2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n436_), .B1(new_n431_), .B2(new_n434_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n413_), .A2(new_n419_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n433_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT90), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n428_), .A2(new_n432_), .B1(new_n438_), .B2(new_n437_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT90), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n410_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n397_), .A2(KEYINPUT29), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n440_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(KEYINPUT91), .A3(new_n410_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT91), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n442_), .B1(new_n397_), .B2(KEYINPUT29), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n449_), .B1(new_n450_), .B2(new_n409_), .ZN(new_n451_));
  AOI221_X4 g250(.A(new_n408_), .B1(new_n445_), .B2(new_n446_), .C1(new_n448_), .C2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n408_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n448_), .A2(new_n451_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n445_), .A2(new_n446_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n453_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n406_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT91), .B1(new_n447_), .B2(new_n410_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n450_), .A2(new_n449_), .A3(new_n409_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n455_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n408_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n404_), .A2(new_n405_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n454_), .A2(new_n453_), .A3(new_n455_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n457_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT0), .B(G57gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(G85gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(G1gat), .B(G29gat), .Z(new_n469_));
  XOR2_X1   g268(.A(new_n468_), .B(new_n469_), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT94), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n397_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n338_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n338_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n475_), .B1(new_n397_), .B2(new_n472_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G225gat), .A2(G233gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(KEYINPUT4), .A3(new_n476_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT4), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n475_), .A2(new_n482_), .A3(new_n397_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n478_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n471_), .B1(new_n480_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT95), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(KEYINPUT33), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(KEYINPUT33), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n471_), .B(new_n488_), .C1(new_n480_), .C2(new_n484_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n364_), .ZN(new_n491_));
  AOI221_X4 g290(.A(KEYINPUT90), .B1(new_n437_), .B2(new_n438_), .C1(new_n428_), .C2(new_n432_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n443_), .B1(new_n433_), .B2(new_n439_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G226gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT19), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT20), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n347_), .B1(G183gat), .B2(G190gat), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n363_), .A2(new_n349_), .B1(new_n354_), .B2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n498_), .B1(new_n442_), .B2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n494_), .A2(new_n497_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT93), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n441_), .A2(new_n364_), .A3(new_n444_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT20), .B1(new_n442_), .B2(new_n500_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n496_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT18), .B(G64gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(G92gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G8gat), .B(G36gat), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n511_), .B(new_n512_), .Z(new_n513_));
  NAND4_X1  g312(.A1(new_n494_), .A2(KEYINPUT93), .A3(new_n497_), .A4(new_n501_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n504_), .A2(new_n509_), .A3(new_n513_), .A4(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n504_), .A2(new_n509_), .A3(new_n514_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n513_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n477_), .A2(new_n479_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n481_), .A2(new_n478_), .A3(new_n483_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(new_n470_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n490_), .A2(new_n515_), .A3(new_n518_), .A4(new_n521_), .ZN(new_n522_));
  OR3_X1    g321(.A1(new_n480_), .A2(new_n484_), .A3(new_n471_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n485_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n513_), .A2(KEYINPUT32), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT96), .B1(new_n516_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n505_), .A2(new_n497_), .A3(new_n507_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n494_), .A2(new_n501_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n527_), .A2(KEYINPUT97), .B1(new_n528_), .B2(new_n496_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n528_), .A2(KEYINPUT97), .A3(new_n496_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n525_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  OR3_X1    g330(.A1(new_n516_), .A2(KEYINPUT96), .A3(new_n525_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n524_), .A2(new_n526_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n466_), .B1(new_n522_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n518_), .A2(new_n515_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT27), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n517_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(KEYINPUT27), .A3(new_n515_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n540_), .A2(new_n524_), .A3(new_n465_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n373_), .B1(new_n534_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT99), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n537_), .A2(new_n465_), .A3(new_n539_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT98), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n537_), .A2(new_n465_), .A3(KEYINPUT98), .A4(new_n539_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n524_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n372_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n543_), .B1(new_n548_), .B2(new_n552_), .ZN(new_n553_));
  AOI211_X1 g352(.A(KEYINPUT99), .B(new_n551_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n542_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n321_), .B(new_n235_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT76), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G229gat), .A2(G233gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n237_), .A2(new_n321_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT77), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n321_), .A2(new_n235_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT77), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n237_), .A2(new_n565_), .A3(new_n321_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n563_), .A2(new_n559_), .A3(new_n564_), .A4(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n561_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(G197gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT78), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(new_n358_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT79), .B1(new_n568_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT79), .ZN(new_n574_));
  INV_X1    g373(.A(new_n572_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n561_), .A2(new_n574_), .A3(new_n567_), .A4(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n568_), .A2(new_n572_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n580_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n333_), .A2(new_n555_), .A3(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(new_n315_), .A3(new_n524_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT38), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n306_), .A2(new_n330_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n579_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT100), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n555_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n586_), .A2(KEYINPUT100), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n588_), .A2(new_n273_), .A3(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n590_), .A2(new_n524_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n584_), .B1(new_n315_), .B2(new_n591_), .ZN(G1324gat));
  NAND3_X1  g391(.A1(new_n582_), .A2(new_n316_), .A3(new_n540_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n590_), .A2(new_n540_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(G8gat), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n595_), .A2(KEYINPUT39), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(KEYINPUT39), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n593_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g398(.A(new_n373_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n313_), .B1(new_n590_), .B2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT41), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n582_), .A2(new_n313_), .A3(new_n600_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(G1326gat));
  INV_X1    g403(.A(G22gat), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n582_), .A2(new_n605_), .A3(new_n466_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n590_), .A2(new_n466_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(G22gat), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n608_), .A2(KEYINPUT42), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(KEYINPUT42), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n606_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT101), .Z(G1327gat));
  AND2_X1   g411(.A1(new_n555_), .A2(new_n273_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n330_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n306_), .A2(new_n580_), .A3(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(G29gat), .B1(new_n616_), .B2(new_n524_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT43), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n555_), .A2(new_n618_), .A3(new_n275_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n555_), .B2(new_n275_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n615_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT44), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(KEYINPUT44), .B(new_n615_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(new_n549_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n617_), .B1(new_n626_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g426(.A1(new_n623_), .A2(new_n540_), .A3(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(G36gat), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT102), .ZN(new_n630_));
  INV_X1    g429(.A(G36gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n616_), .A2(new_n631_), .A3(new_n540_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT45), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(new_n634_), .A3(G36gat), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n630_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n636_), .A2(new_n637_), .A3(KEYINPUT46), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT46), .B1(new_n636_), .B2(new_n637_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1329gat));
  INV_X1    g439(.A(new_n616_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n233_), .B1(new_n641_), .B2(new_n373_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n550_), .A2(G43gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n642_), .B1(new_n625_), .B2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n646_), .B1(new_n625_), .B2(new_n465_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n623_), .A2(KEYINPUT104), .A3(new_n466_), .A4(new_n624_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(G50gat), .A3(new_n648_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n465_), .A2(G50gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n641_), .B2(new_n650_), .ZN(G1331gat));
  INV_X1    g450(.A(new_n306_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(new_n579_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n555_), .A2(new_n614_), .A3(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(new_n261_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(G57gat), .A3(new_n524_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT105), .ZN(new_n657_));
  INV_X1    g456(.A(new_n275_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n654_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(G57gat), .B1(new_n659_), .B2(new_n524_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n657_), .A2(new_n660_), .ZN(G1332gat));
  NAND2_X1  g460(.A1(new_n655_), .A2(new_n540_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G64gat), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT106), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n662_), .A2(new_n665_), .A3(G64gat), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT48), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n664_), .A2(KEYINPUT48), .A3(new_n666_), .ZN(new_n670_));
  INV_X1    g469(.A(G64gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n659_), .A2(new_n671_), .A3(new_n540_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(new_n670_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n669_), .A2(new_n670_), .A3(KEYINPUT107), .A4(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1333gat));
  INV_X1    g476(.A(G71gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n655_), .B2(new_n600_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT49), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n659_), .A2(new_n678_), .A3(new_n600_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1334gat));
  INV_X1    g481(.A(G78gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n655_), .B2(new_n466_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT109), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n684_), .B(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n659_), .A2(new_n683_), .A3(new_n466_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT110), .ZN(G1335gat));
  NAND3_X1  g489(.A1(new_n613_), .A2(new_n330_), .A3(new_n653_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT111), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G85gat), .B1(new_n693_), .B2(new_n524_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n619_), .A2(new_n620_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n653_), .A2(new_n330_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT112), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT113), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(new_n524_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n694_), .B1(new_n700_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g500(.A(G92gat), .B1(new_n693_), .B2(new_n540_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n540_), .A2(G92gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n699_), .B2(new_n703_), .ZN(G1337gat));
  INV_X1    g503(.A(G99gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n699_), .B2(new_n600_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n693_), .A2(new_n210_), .A3(new_n550_), .ZN(new_n707_));
  OR3_X1    g506(.A1(new_n706_), .A2(KEYINPUT51), .A3(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT51), .B1(new_n706_), .B2(new_n707_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1338gat));
  XNOR2_X1  g509(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n695_), .A2(new_n466_), .A3(new_n697_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT114), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT114), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n695_), .A2(new_n714_), .A3(new_n466_), .A4(new_n697_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n713_), .A2(G106gat), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT52), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n713_), .A2(new_n718_), .A3(G106gat), .A4(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n693_), .A2(new_n211_), .A3(new_n466_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n711_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n711_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n721_), .ZN(new_n724_));
  AOI211_X1 g523(.A(new_n723_), .B(new_n724_), .C1(new_n717_), .C2(new_n719_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n722_), .A2(new_n725_), .ZN(G1339gat));
  NAND4_X1  g525(.A1(new_n267_), .A2(new_n585_), .A3(new_n580_), .A4(new_n274_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT54), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT57), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT55), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n293_), .B2(new_n288_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n293_), .A2(new_n288_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n293_), .A2(new_n730_), .A3(new_n288_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n301_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT56), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT56), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n737_), .B(new_n301_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n294_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n300_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n736_), .A2(new_n579_), .A3(new_n738_), .A4(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n303_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n558_), .A2(new_n559_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n563_), .A2(new_n560_), .A3(new_n564_), .A4(new_n566_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(new_n572_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n742_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n741_), .A2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n729_), .B1(new_n748_), .B2(new_n261_), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT57), .B(new_n273_), .C1(new_n741_), .C2(new_n747_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n736_), .A2(new_n746_), .A3(new_n738_), .A4(new_n740_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT58), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n735_), .A2(KEYINPUT56), .B1(new_n739_), .B2(new_n300_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n755_), .A2(KEYINPUT58), .A3(new_n746_), .A4(new_n738_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n274_), .B2(new_n267_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n330_), .B1(new_n751_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n728_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n548_), .A2(new_n524_), .A3(new_n550_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n761_), .A2(KEYINPUT59), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n764_), .B1(new_n751_), .B2(new_n758_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n748_), .A2(new_n261_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT57), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n748_), .A2(new_n729_), .A3(new_n261_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n275_), .A2(new_n754_), .A3(new_n756_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(KEYINPUT116), .A3(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n765_), .A2(new_n330_), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n761_), .B1(new_n772_), .B2(new_n728_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT59), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n763_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G113gat), .B1(new_n775_), .B2(new_n580_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n773_), .A2(KEYINPUT117), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n778_));
  AOI211_X1 g577(.A(new_n778_), .B(new_n761_), .C1(new_n772_), .C2(new_n728_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n335_), .B(new_n579_), .C1(new_n777_), .C2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n776_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n776_), .B2(new_n780_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1340gat));
  OR2_X1    g583(.A1(new_n777_), .A2(new_n779_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n337_), .B1(new_n652_), .B2(KEYINPUT60), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n785_), .B(new_n786_), .C1(KEYINPUT60), .C2(new_n337_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n775_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n306_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n787_), .B1(new_n337_), .B2(new_n790_), .ZN(G1341gat));
  AOI21_X1  g590(.A(G127gat), .B1(new_n785_), .B2(new_n614_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n788_), .A2(G127gat), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n614_), .B2(new_n794_), .ZN(G1342gat));
  AOI21_X1  g594(.A(G134gat), .B1(new_n785_), .B2(new_n273_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT119), .B(G134gat), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n658_), .A2(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT120), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n796_), .B1(new_n788_), .B2(new_n799_), .ZN(G1343gat));
  AOI21_X1  g599(.A(new_n600_), .B1(new_n772_), .B2(new_n728_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n540_), .ZN(new_n802_));
  AND4_X1   g601(.A1(new_n524_), .A2(new_n801_), .A3(new_n466_), .A4(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n579_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n306_), .ZN(new_n806_));
  XOR2_X1   g605(.A(KEYINPUT121), .B(G148gat), .Z(new_n807_));
  XNOR2_X1  g606(.A(new_n806_), .B(new_n807_), .ZN(G1345gat));
  NAND2_X1  g607(.A1(new_n803_), .A2(new_n614_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(KEYINPUT61), .B(G155gat), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n809_), .B(new_n810_), .ZN(G1346gat));
  AOI21_X1  g610(.A(G162gat), .B1(new_n803_), .B2(new_n273_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n275_), .A2(G162gat), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT122), .Z(new_n814_));
  AOI21_X1  g613(.A(new_n812_), .B1(new_n803_), .B2(new_n814_), .ZN(G1347gat));
  NOR4_X1   g614(.A1(new_n373_), .A2(new_n802_), .A3(new_n524_), .A4(new_n466_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n760_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n579_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(G169gat), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT123), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT62), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n821_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n818_), .A2(G169gat), .A3(new_n823_), .A4(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n353_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n822_), .B(new_n825_), .C1(new_n826_), .C2(new_n818_), .ZN(G1348gat));
  AOI21_X1  g626(.A(G176gat), .B1(new_n817_), .B2(new_n306_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n299_), .B(new_n652_), .C1(new_n772_), .C2(new_n728_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n816_), .ZN(G1349gat));
  NAND2_X1  g629(.A1(new_n817_), .A2(new_n614_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(G183gat), .ZN(new_n832_));
  INV_X1    g631(.A(new_n355_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n831_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT124), .ZN(G1350gat));
  INV_X1    g634(.A(new_n817_), .ZN(new_n836_));
  OAI21_X1  g635(.A(G190gat), .B1(new_n836_), .B2(new_n658_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n817_), .A2(new_n273_), .A3(new_n356_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(G1351gat));
  XNOR2_X1  g638(.A(KEYINPUT126), .B(G197gat), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n802_), .A2(new_n524_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n801_), .A2(new_n466_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT125), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n801_), .A2(KEYINPUT125), .A3(new_n466_), .A4(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n840_), .B1(new_n846_), .B2(new_n579_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n840_), .ZN(new_n848_));
  AOI211_X1 g647(.A(new_n580_), .B(new_n848_), .C1(new_n844_), .C2(new_n845_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n849_), .ZN(G1352gat));
  AOI21_X1  g649(.A(G204gat), .B1(new_n846_), .B2(new_n306_), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n296_), .B(new_n652_), .C1(new_n844_), .C2(new_n845_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1353gat));
  OR2_X1    g652(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n846_), .B2(new_n614_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT63), .B(G211gat), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n330_), .B(new_n856_), .C1(new_n844_), .C2(new_n845_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1354gat));
  XOR2_X1   g657(.A(KEYINPUT127), .B(G218gat), .Z(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n846_), .B2(new_n273_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n859_), .ZN(new_n861_));
  AOI211_X1 g660(.A(new_n658_), .B(new_n861_), .C1(new_n844_), .C2(new_n845_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1355gat));
endmodule


