//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G1gat), .B(G8gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT68), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT69), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n206_), .A2(KEYINPUT68), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT69), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n206_), .A2(KEYINPUT68), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n208_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G15gat), .A2(G22gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G15gat), .A2(G22gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G1gat), .A2(G8gat), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n215_), .A2(new_n216_), .B1(KEYINPUT14), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n213_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n208_), .A2(new_n212_), .A3(new_n218_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n205_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT72), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n220_), .A2(new_n225_), .A3(new_n221_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT73), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n220_), .A2(new_n221_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n223_), .B1(new_n230_), .B2(new_n204_), .ZN(new_n231_));
  AOI211_X1 g030(.A(KEYINPUT72), .B(new_n205_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n232_));
  OAI22_X1  g031(.A1(new_n231_), .A2(new_n232_), .B1(new_n204_), .B2(new_n230_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n228_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G113gat), .B(G141gat), .Z(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT75), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G169gat), .B(G197gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n238_), .B(new_n239_), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(KEYINPUT74), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n236_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n236_), .A2(new_n242_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT76), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT76), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT96), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT95), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT23), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n254_), .A2(KEYINPUT80), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(KEYINPUT80), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n253_), .A2(KEYINPUT23), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(G183gat), .B2(G190gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT81), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n260_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT22), .B(G169gat), .ZN(new_n263_));
  INV_X1    g062(.A(G176gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT79), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n261_), .A2(new_n262_), .A3(new_n266_), .A4(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT25), .B(G183gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G190gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(G169gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n264_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(KEYINPUT24), .A3(new_n267_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT77), .B1(new_n253_), .B2(KEYINPUT23), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(new_n254_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT24), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(new_n272_), .A3(new_n264_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n275_), .B1(new_n280_), .B2(KEYINPUT78), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(KEYINPUT78), .B2(new_n280_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n268_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G197gat), .B(G204gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT88), .ZN(new_n285_));
  INV_X1    g084(.A(G204gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G197gat), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n285_), .B(KEYINPUT21), .C1(KEYINPUT88), .C2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G211gat), .B(G218gat), .Z(new_n289_));
  INV_X1    g088(.A(KEYINPUT21), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n289_), .B1(new_n290_), .B2(new_n284_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n284_), .A2(new_n290_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n288_), .A2(new_n291_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n283_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT20), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n293_), .B(KEYINPUT89), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n277_), .B1(G183gat), .B2(G190gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n258_), .A2(new_n279_), .A3(new_n271_), .A4(new_n274_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n296_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n295_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G226gat), .A2(G233gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT19), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n268_), .A2(new_n282_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n293_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n305_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n299_), .A2(new_n300_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n296_), .B1(new_n310_), .B2(new_n294_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n308_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n252_), .B1(new_n306_), .B2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT95), .B1(new_n303_), .B2(new_n305_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G8gat), .B(G36gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(G64gat), .B(G92gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT32), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n251_), .B1(new_n316_), .B2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G127gat), .B(G134gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G113gat), .B(G120gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n333_), .B(KEYINPUT3), .Z(new_n334_));
  NAND2_X1  g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n335_), .B(KEYINPUT2), .Z(new_n336_));
  OAI211_X1 g135(.A(new_n330_), .B(new_n332_), .C1(new_n334_), .C2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n331_), .B1(KEYINPUT1), .B2(new_n330_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(KEYINPUT1), .B2(new_n330_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n333_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(new_n335_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n329_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT4), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT4), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n329_), .A2(new_n346_), .A3(new_n342_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G1gat), .B(G29gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G57gat), .B(G85gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n344_), .A2(new_n349_), .ZN(new_n357_));
  OR3_X1    g156(.A1(new_n350_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n356_), .B1(new_n350_), .B2(new_n357_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n315_), .A2(KEYINPUT96), .A3(KEYINPUT32), .A4(new_n322_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n308_), .A2(new_n311_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n362_), .A2(new_n309_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT91), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT90), .B1(new_n310_), .B2(new_n294_), .ZN(new_n365_));
  OR3_X1    g164(.A1(new_n310_), .A2(KEYINPUT90), .A3(new_n294_), .ZN(new_n366_));
  AOI211_X1 g165(.A(new_n296_), .B(new_n305_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n364_), .B1(new_n367_), .B2(new_n295_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n364_), .A3(new_n295_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n363_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n323_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n324_), .A2(new_n360_), .A3(new_n361_), .A4(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n359_), .B(KEYINPUT33), .ZN(new_n374_));
  INV_X1    g173(.A(new_n370_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(new_n368_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n321_), .B1(new_n376_), .B2(new_n363_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n371_), .A2(new_n322_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n356_), .B1(new_n344_), .B2(new_n349_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n380_), .B(KEYINPUT94), .Z(new_n381_));
  NAND4_X1  g180(.A1(new_n374_), .A2(new_n377_), .A3(new_n378_), .A4(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n373_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G228gat), .A2(G233gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n384_), .B(KEYINPUT87), .Z(new_n385_));
  AND2_X1   g184(.A1(new_n342_), .A2(KEYINPUT29), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n385_), .B1(new_n386_), .B2(new_n293_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n386_), .A2(new_n385_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(new_n297_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n342_), .A2(KEYINPUT29), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G22gat), .B(G50gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n389_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G78gat), .B(G106gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n393_), .B(new_n396_), .Z(new_n397_));
  XNOR2_X1  g196(.A(G71gat), .B(G99gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(G43gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n329_), .B(KEYINPUT31), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G227gat), .A2(G233gat), .ZN(new_n404_));
  INV_X1    g203(.A(G15gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n283_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n283_), .A2(new_n406_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  OR3_X1    g209(.A1(new_n407_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n410_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n403_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(new_n403_), .A3(new_n412_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n399_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n415_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n399_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n417_), .A2(new_n413_), .A3(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n383_), .A2(new_n397_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n416_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n419_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n397_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n397_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n377_), .A2(new_n378_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT27), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n315_), .A2(new_n321_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n429_), .B1(new_n371_), .B2(new_n322_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n428_), .A2(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n360_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n427_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n250_), .B1(new_n421_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT37), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT64), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n437_), .A2(KEYINPUT9), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(KEYINPUT9), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(G85gat), .ZN(new_n441_));
  INV_X1    g240(.A(G92gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(KEYINPUT9), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G85gat), .A2(G92gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n440_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n438_), .A2(new_n444_), .A3(new_n443_), .A4(new_n439_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G99gat), .A2(G106gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT6), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT6), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(G99gat), .A3(G106gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  OR2_X1    g251(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n453_));
  INV_X1    g252(.A(G106gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n446_), .A2(new_n447_), .A3(new_n452_), .A4(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G85gat), .B(G92gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AOI211_X1 g261(.A(KEYINPUT8), .B(new_n458_), .C1(new_n462_), .C2(new_n452_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT8), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT7), .ZN(new_n465_));
  INV_X1    g264(.A(G99gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n454_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n450_), .B1(G99gat), .B2(G106gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n448_), .A2(KEYINPUT6), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n459_), .B(new_n467_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n458_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n464_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n457_), .B1(new_n463_), .B2(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n225_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G232gat), .A2(G233gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT34), .ZN(new_n476_));
  OAI22_X1  g275(.A1(new_n473_), .A2(new_n205_), .B1(KEYINPUT35), .B2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(KEYINPUT35), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT66), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n479_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G190gat), .B(G218gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G134gat), .B(G162gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n486_), .A2(KEYINPUT36), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n483_), .B(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n480_), .A2(new_n482_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(KEYINPUT36), .A3(new_n486_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n436_), .B1(new_n492_), .B2(KEYINPUT67), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT67), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n494_), .A3(KEYINPUT37), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G231gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n230_), .B(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(KEYINPUT65), .B(G71gat), .Z(new_n499_));
  INV_X1    g298(.A(G78gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT65), .B(G71gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(G78gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G57gat), .B(G64gat), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n501_), .A2(new_n503_), .B1(KEYINPUT11), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT11), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n504_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n501_), .A2(new_n503_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n505_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n498_), .B(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G127gat), .B(G155gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT70), .B(KEYINPUT16), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G183gat), .B(G211gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT17), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n512_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n512_), .A2(KEYINPUT17), .A3(new_n517_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT71), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n521_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n519_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(G230gat), .ZN(new_n526_));
  INV_X1    g325(.A(G233gat), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n470_), .A2(new_n471_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT8), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n470_), .A2(new_n464_), .A3(new_n471_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n456_), .A2(new_n452_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n445_), .B2(new_n440_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n530_), .A2(new_n531_), .B1(new_n533_), .B2(new_n447_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n528_), .B1(new_n534_), .B2(new_n511_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT12), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n537_));
  INV_X1    g336(.A(new_n503_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n502_), .A2(G78gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n540_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n473_), .A2(new_n536_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n536_), .B1(new_n473_), .B2(new_n541_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n535_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n534_), .A2(new_n511_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n473_), .A2(new_n541_), .ZN(new_n547_));
  AOI211_X1 g346(.A(new_n526_), .B(new_n527_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G120gat), .B(G148gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT5), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G176gat), .B(G204gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  NOR3_X1   g351(.A1(new_n545_), .A2(new_n548_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n552_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n557_), .A2(KEYINPUT13), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(KEYINPUT13), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n496_), .A2(new_n525_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n435_), .A2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n360_), .B(KEYINPUT97), .Z(new_n563_));
  NOR3_X1   g362(.A1(new_n562_), .A2(G1gat), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT38), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT98), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT38), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n491_), .B1(new_n421_), .B2(new_n434_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n560_), .A2(new_n246_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT99), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n570_), .A2(new_n525_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n360_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n567_), .B1(new_n574_), .B2(G1gat), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n566_), .B1(new_n575_), .B2(new_n564_), .ZN(G1324gat));
  NOR3_X1   g375(.A1(new_n562_), .A2(G8gat), .A3(new_n432_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT100), .ZN(new_n578_));
  OAI21_X1  g377(.A(G8gat), .B1(new_n572_), .B2(new_n432_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT39), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n580_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n578_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n583_), .B(new_n585_), .ZN(G1325gat));
  OAI21_X1  g385(.A(G15gat), .B1(new_n572_), .B2(new_n420_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n588_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n562_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n420_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n405_), .A3(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n589_), .A2(new_n590_), .A3(new_n593_), .ZN(G1326gat));
  OAI21_X1  g393(.A(G22gat), .B1(new_n572_), .B2(new_n397_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n595_), .A2(KEYINPUT42), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(KEYINPUT42), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n397_), .A2(G22gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT103), .Z(new_n599_));
  OAI22_X1  g398(.A1(new_n596_), .A2(new_n597_), .B1(new_n562_), .B2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT104), .Z(G1327gat));
  NAND2_X1  g400(.A1(new_n525_), .A2(new_n491_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(new_n560_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n435_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(G29gat), .B1(new_n605_), .B2(new_n360_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n570_), .A2(new_n524_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT43), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n421_), .A2(new_n434_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(new_n496_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n496_), .ZN(new_n611_));
  AOI211_X1 g410(.A(KEYINPUT43), .B(new_n611_), .C1(new_n421_), .C2(new_n434_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n607_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT44), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  OAI211_X1 g414(.A(KEYINPUT44), .B(new_n607_), .C1(new_n610_), .C2(new_n612_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n563_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n618_), .A2(G29gat), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n606_), .B1(new_n617_), .B2(new_n619_), .ZN(G1328gat));
  NOR2_X1   g419(.A1(new_n432_), .A2(G36gat), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n435_), .A2(new_n603_), .A3(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT45), .Z(new_n623_));
  INV_X1    g422(.A(new_n432_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n615_), .A2(new_n624_), .A3(new_n616_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n623_), .B1(new_n625_), .B2(G36gat), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT105), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT46), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n626_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n627_), .A2(new_n628_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n626_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n629_), .A2(new_n632_), .ZN(G1329gat));
  INV_X1    g432(.A(G43gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n420_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n615_), .A2(new_n616_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT106), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT106), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n615_), .A2(new_n638_), .A3(new_n616_), .A4(new_n635_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n634_), .B1(new_n604_), .B2(new_n420_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n637_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT47), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT47), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n637_), .A2(new_n643_), .A3(new_n639_), .A4(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1330gat));
  AOI21_X1  g444(.A(G50gat), .B1(new_n605_), .B2(new_n424_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n424_), .A2(G50gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n617_), .B2(new_n647_), .ZN(G1331gat));
  AOI21_X1  g447(.A(new_n245_), .B1(new_n421_), .B2(new_n434_), .ZN(new_n649_));
  AND4_X1   g448(.A1(new_n524_), .A2(new_n649_), .A3(new_n560_), .A4(new_n611_), .ZN(new_n650_));
  INV_X1    g449(.A(G57gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n618_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n568_), .A2(new_n524_), .A3(new_n560_), .A4(new_n250_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT107), .Z(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(new_n360_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n652_), .B1(new_n655_), .B2(new_n651_), .ZN(G1332gat));
  INV_X1    g455(.A(G64gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n650_), .A2(new_n657_), .A3(new_n624_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT48), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n654_), .A2(new_n624_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(G64gat), .ZN(new_n661_));
  AOI211_X1 g460(.A(KEYINPUT48), .B(new_n657_), .C1(new_n654_), .C2(new_n624_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n658_), .B1(new_n661_), .B2(new_n662_), .ZN(G1333gat));
  INV_X1    g462(.A(G71gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n650_), .A2(new_n664_), .A3(new_n592_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT49), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n654_), .A2(new_n592_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n667_), .B2(G71gat), .ZN(new_n668_));
  AOI211_X1 g467(.A(KEYINPUT49), .B(new_n664_), .C1(new_n654_), .C2(new_n592_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(G1334gat));
  NAND3_X1  g469(.A1(new_n650_), .A2(new_n500_), .A3(new_n424_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT50), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n654_), .A2(new_n424_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n673_), .B2(G78gat), .ZN(new_n674_));
  AOI211_X1 g473(.A(KEYINPUT50), .B(new_n500_), .C1(new_n654_), .C2(new_n424_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(G1335gat));
  INV_X1    g475(.A(new_n560_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n602_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n649_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n680_), .A2(new_n441_), .A3(new_n618_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n677_), .A2(new_n524_), .A3(new_n245_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT109), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n609_), .A2(new_n496_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT43), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n609_), .A2(new_n608_), .A3(new_n496_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT108), .ZN(new_n688_));
  OR3_X1    g487(.A1(new_n610_), .A2(new_n612_), .A3(KEYINPUT108), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n683_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(new_n360_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n681_), .B1(new_n691_), .B2(new_n441_), .ZN(G1336gat));
  NAND3_X1  g491(.A1(new_n680_), .A2(new_n442_), .A3(new_n624_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n690_), .A2(new_n624_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(new_n442_), .ZN(G1337gat));
  NAND2_X1  g494(.A1(new_n453_), .A2(new_n455_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n679_), .A2(new_n420_), .A3(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n690_), .A2(new_n592_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n698_), .B(new_n699_), .C1(new_n700_), .C2(new_n466_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n699_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n466_), .B1(new_n690_), .B2(new_n592_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(new_n697_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(G1338gat));
  NOR2_X1   g504(.A1(new_n683_), .A2(new_n397_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n454_), .B1(new_n687_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT52), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n680_), .A2(new_n454_), .A3(new_n424_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT53), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT53), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n713_), .A3(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1339gat));
  NOR2_X1   g514(.A1(new_n496_), .A2(new_n560_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n250_), .A2(KEYINPUT111), .A3(new_n524_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n247_), .A2(new_n524_), .A3(new_n249_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n716_), .A2(new_n717_), .A3(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n716_), .A2(new_n717_), .A3(new_n720_), .A4(new_n722_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n224_), .A2(new_n227_), .A3(new_n234_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n233_), .A2(new_n228_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n241_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n240_), .B1(new_n229_), .B2(new_n235_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n556_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n546_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n544_), .A2(KEYINPUT55), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT55), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n535_), .B(new_n736_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n737_));
  AOI221_X4 g536(.A(new_n733_), .B1(new_n734_), .B2(new_n528_), .C1(new_n735_), .C2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n735_), .A2(new_n737_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n734_), .A2(new_n528_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT113), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n552_), .B1(new_n738_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT56), .ZN(new_n745_));
  OAI211_X1 g544(.A(KEYINPUT114), .B(new_n552_), .C1(new_n738_), .C2(new_n741_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n744_), .A2(KEYINPUT115), .A3(new_n745_), .A4(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n553_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  OAI211_X1 g548(.A(KEYINPUT56), .B(new_n552_), .C1(new_n738_), .C2(new_n741_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT56), .B1(new_n742_), .B2(new_n743_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n746_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n732_), .B1(new_n749_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT57), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n491_), .A2(new_n756_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n755_), .A2(KEYINPUT118), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT118), .B1(new_n755_), .B2(new_n757_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n755_), .A2(new_n492_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n554_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n742_), .A2(new_n745_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n750_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT117), .B1(new_n764_), .B2(KEYINPUT116), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT117), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(KEYINPUT58), .ZN(new_n768_));
  OAI22_X1  g567(.A1(new_n765_), .A2(KEYINPUT58), .B1(new_n764_), .B2(new_n768_), .ZN(new_n769_));
  AOI22_X1  g568(.A1(new_n761_), .A2(new_n756_), .B1(new_n769_), .B2(new_n496_), .ZN(new_n770_));
  AOI211_X1 g569(.A(KEYINPUT120), .B(new_n524_), .C1(new_n760_), .C2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT120), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n761_), .A2(new_n756_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n755_), .A2(new_n757_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n769_), .A2(new_n496_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n755_), .A2(KEYINPUT118), .A3(new_n757_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n773_), .A2(new_n776_), .A3(new_n777_), .A4(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n772_), .B1(new_n779_), .B2(new_n525_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n727_), .B1(new_n771_), .B2(new_n780_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n624_), .A2(new_n426_), .A3(new_n563_), .ZN(new_n782_));
  XOR2_X1   g581(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n524_), .B1(new_n760_), .B2(new_n770_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n785_), .A2(new_n726_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n782_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT59), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n784_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(G113gat), .B1(new_n789_), .B2(new_n250_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n786_), .A2(new_n787_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n246_), .A2(G113gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n790_), .B1(new_n792_), .B2(new_n793_), .ZN(G1340gat));
  INV_X1    g593(.A(KEYINPUT122), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n789_), .B2(new_n677_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n784_), .A2(KEYINPUT122), .A3(new_n560_), .A4(new_n788_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(G120gat), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT60), .ZN(new_n799_));
  AOI21_X1  g598(.A(G120gat), .B1(new_n560_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT121), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT121), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n799_), .B2(G120gat), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n791_), .B(new_n801_), .C1(new_n800_), .C2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n798_), .A2(new_n804_), .ZN(G1341gat));
  OAI21_X1  g604(.A(G127gat), .B1(new_n789_), .B2(new_n525_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n525_), .A2(G127gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n792_), .B2(new_n807_), .ZN(G1342gat));
  NAND2_X1  g607(.A1(new_n496_), .A2(G134gat), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT123), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n784_), .A2(new_n788_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(G134gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n792_), .B2(new_n492_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT124), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n811_), .A2(new_n813_), .A3(KEYINPUT124), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(G1343gat));
  INV_X1    g617(.A(new_n786_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n624_), .A2(new_n425_), .A3(new_n563_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n245_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n560_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g625(.A1(new_n821_), .A2(new_n525_), .ZN(new_n827_));
  XOR2_X1   g626(.A(KEYINPUT61), .B(G155gat), .Z(new_n828_));
  XNOR2_X1  g627(.A(new_n827_), .B(new_n828_), .ZN(G1346gat));
  OAI21_X1  g628(.A(G162gat), .B1(new_n821_), .B2(new_n611_), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n492_), .A2(G162gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n821_), .B2(new_n831_), .ZN(G1347gat));
  INV_X1    g631(.A(KEYINPUT125), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n618_), .A2(new_n432_), .A3(new_n420_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n397_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n781_), .A2(new_n245_), .A3(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n781_), .A2(new_n263_), .A3(new_n245_), .A4(new_n836_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT62), .B1(new_n837_), .B2(G169gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n833_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n837_), .A2(G169gat), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT62), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n845_), .A2(KEYINPUT125), .A3(new_n839_), .A4(new_n838_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(G1348gat));
  NAND3_X1  g646(.A1(new_n781_), .A2(new_n560_), .A3(new_n836_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n786_), .A2(new_n424_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n834_), .A2(G176gat), .A3(new_n560_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n848_), .A2(new_n264_), .B1(new_n849_), .B2(new_n850_), .ZN(G1349gat));
  INV_X1    g650(.A(KEYINPUT126), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n781_), .A2(new_n836_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n525_), .A2(new_n269_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n852_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n849_), .A2(new_n524_), .A3(new_n834_), .ZN(new_n857_));
  INV_X1    g656(.A(G183gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n781_), .A2(KEYINPUT126), .A3(new_n836_), .A4(new_n854_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n856_), .A2(new_n859_), .A3(new_n860_), .ZN(G1350gat));
  OAI21_X1  g660(.A(G190gat), .B1(new_n853_), .B2(new_n611_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n491_), .A2(new_n270_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n853_), .B2(new_n863_), .ZN(G1351gat));
  NAND3_X1  g663(.A1(new_n420_), .A2(new_n433_), .A3(new_n424_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT127), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n624_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n866_), .B2(new_n865_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n819_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n245_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g671(.A1(new_n869_), .A2(new_n677_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n286_), .ZN(G1353gat));
  NAND2_X1  g673(.A1(new_n870_), .A2(new_n524_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n876_));
  AND2_X1   g675(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n875_), .B2(new_n876_), .ZN(G1354gat));
  OAI21_X1  g678(.A(G218gat), .B1(new_n869_), .B2(new_n611_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n492_), .A2(G218gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n869_), .B2(new_n881_), .ZN(G1355gat));
endmodule


