//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_;
  XNOR2_X1  g000(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n202_));
  XOR2_X1   g001(.A(G22gat), .B(G50gat), .Z(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G141gat), .ZN(new_n205_));
  INV_X1    g004(.A(G148gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT3), .ZN(new_n208_));
  OR3_X1    g007(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n208_), .A2(new_n209_), .A3(new_n212_), .A4(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT84), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(KEYINPUT84), .A3(new_n216_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n214_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n216_), .A2(KEYINPUT1), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n215_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n216_), .A2(KEYINPUT1), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n210_), .B(new_n207_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT85), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n221_), .A2(KEYINPUT85), .A3(new_n225_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT29), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n204_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n230_), .A2(new_n231_), .A3(new_n204_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n202_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n234_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n202_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n232_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G211gat), .B(G218gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT21), .B1(new_n240_), .B2(KEYINPUT89), .ZN(new_n241_));
  XOR2_X1   g040(.A(G197gat), .B(G204gat), .Z(new_n242_));
  OAI211_X1 g041(.A(new_n241_), .B(new_n242_), .C1(KEYINPUT21), .C2(new_n240_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n244_), .B(KEYINPUT21), .C1(KEYINPUT89), .C2(new_n240_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G228gat), .ZN(new_n248_));
  INV_X1    g047(.A(G233gat), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n249_), .A2(KEYINPUT88), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(KEYINPUT88), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n248_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n247_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n228_), .A2(KEYINPUT29), .A3(new_n229_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n221_), .A2(new_n225_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n246_), .B1(new_n255_), .B2(new_n231_), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n253_), .A2(new_n254_), .B1(new_n256_), .B2(new_n252_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G78gat), .B(G106gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT90), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT91), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n239_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n257_), .B(new_n260_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT87), .B1(new_n235_), .B2(new_n238_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n237_), .B1(new_n236_), .B2(new_n232_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n233_), .A2(new_n202_), .A3(new_n234_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT87), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n263_), .B1(new_n264_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT27), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G226gat), .A2(G233gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT20), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT23), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(G183gat), .B2(G190gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT22), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G169gat), .ZN(new_n285_));
  INV_X1    g084(.A(G169gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT22), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G176gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n283_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n281_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT26), .B(G190gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT25), .B(G183gat), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n294_), .A2(KEYINPUT93), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(KEYINPUT93), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n293_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT79), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n300_), .A2(KEYINPUT24), .A3(new_n282_), .A4(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT24), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n280_), .A3(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n291_), .B1(new_n297_), .B2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n278_), .B1(new_n306_), .B2(new_n246_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT78), .B(G183gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n280_), .B1(new_n309_), .B2(G190gat), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n285_), .A2(KEYINPUT80), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n285_), .A2(KEYINPUT80), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n311_), .A2(new_n289_), .A3(new_n312_), .A4(new_n287_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n313_), .A3(new_n282_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT25), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n308_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n292_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n298_), .B(new_n299_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n303_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n318_), .A2(new_n280_), .A3(new_n320_), .A4(new_n302_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n247_), .A2(new_n314_), .A3(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n277_), .B1(new_n307_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT20), .B1(new_n306_), .B2(new_n246_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n321_), .A2(new_n314_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n326_));
  OR3_X1    g125(.A1(new_n325_), .A2(new_n326_), .A3(new_n276_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT18), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n324_), .A2(new_n327_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n325_), .A2(new_n326_), .A3(new_n276_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n331_), .B1(new_n335_), .B2(new_n323_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n273_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n276_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n307_), .A2(new_n322_), .A3(new_n277_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n331_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n333_), .A2(new_n342_), .A3(KEYINPUT27), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n338_), .A2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n272_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT96), .B(G85gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT0), .B(G57gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G127gat), .B(G134gat), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n351_), .A2(KEYINPUT83), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(KEYINPUT83), .ZN(new_n353_));
  XOR2_X1   g152(.A(G113gat), .B(G120gat), .Z(new_n354_));
  OR3_X1    g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n354_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n228_), .A2(new_n357_), .A3(new_n229_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n255_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(KEYINPUT4), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(KEYINPUT94), .Z(new_n362_));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n228_), .A2(new_n357_), .A3(new_n363_), .A4(new_n229_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n360_), .A2(KEYINPUT95), .A3(new_n362_), .A4(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n362_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n358_), .A2(new_n359_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n364_), .A2(new_n362_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT95), .B1(new_n369_), .B2(new_n360_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n350_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT95), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n358_), .A2(KEYINPUT4), .A3(new_n359_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n364_), .A2(new_n362_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n350_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(new_n367_), .A4(new_n365_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n371_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n321_), .A2(new_n314_), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n380_), .B(KEYINPUT30), .Z(new_n381_));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n357_), .B(KEYINPUT31), .Z(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT82), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n383_), .B(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n381_), .A2(new_n382_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G71gat), .B(G99gat), .ZN(new_n388_));
  INV_X1    g187(.A(G43gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G227gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(G15gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n390_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n387_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n386_), .B(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n345_), .A2(new_n379_), .A3(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n338_), .A2(new_n377_), .A3(new_n371_), .A4(new_n343_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n271_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n332_), .A2(KEYINPUT32), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(new_n335_), .B2(new_n323_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n399_), .B2(new_n341_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n378_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT98), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n358_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n364_), .A2(new_n366_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n350_), .B(new_n405_), .C1(new_n373_), .C2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n333_), .A2(new_n407_), .A3(new_n336_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n409_), .B2(new_n377_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n368_), .A2(new_n370_), .A3(new_n350_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(KEYINPUT97), .A3(KEYINPUT33), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT97), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n377_), .B2(new_n409_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n410_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n378_), .A2(KEYINPUT98), .A3(new_n401_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n404_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n398_), .B1(new_n417_), .B2(new_n271_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n396_), .B1(new_n418_), .B2(new_n395_), .ZN(new_n419_));
  INV_X1    g218(.A(G1gat), .ZN(new_n420_));
  INV_X1    g219(.A(G8gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT14), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT71), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(KEYINPUT71), .B(KEYINPUT14), .C1(new_n420_), .C2(new_n421_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G15gat), .B(G22gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT72), .ZN(new_n428_));
  XOR2_X1   g227(.A(G1gat), .B(G8gat), .Z(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G29gat), .B(G36gat), .Z(new_n431_));
  XOR2_X1   g230(.A(G43gat), .B(G50gat), .Z(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT69), .B(KEYINPUT15), .Z(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n430_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n429_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n428_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n428_), .A2(new_n437_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n433_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G229gat), .A2(G233gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n436_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n433_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n430_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n441_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n442_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT74), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT74), .ZN(new_n449_));
  AOI211_X1 g248(.A(new_n449_), .B(new_n442_), .C1(new_n445_), .C2(new_n441_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n443_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G113gat), .B(G141gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT76), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G169gat), .B(G197gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n453_), .B(new_n454_), .Z(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n456_), .A2(KEYINPUT75), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n451_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n440_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n444_), .B1(new_n459_), .B2(new_n438_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n439_), .A2(new_n440_), .A3(new_n433_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n449_), .B1(new_n462_), .B2(new_n442_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n446_), .A2(KEYINPUT74), .A3(new_n447_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n457_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n443_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n458_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT77), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n419_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT66), .B(G92gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT9), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(G85gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT6), .ZN(new_n476_));
  OR2_X1    g275(.A1(G85gat), .A2(G92gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G85gat), .A2(G92gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT9), .A3(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n474_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT64), .ZN(new_n482_));
  AND2_X1   g281(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n482_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT10), .ZN(new_n486_));
  INV_X1    g285(.A(G99gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(KEYINPUT64), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(G106gat), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT65), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT65), .ZN(new_n494_));
  AOI211_X1 g293(.A(new_n494_), .B(G106gat), .C1(new_n485_), .C2(new_n490_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n481_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT67), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n481_), .B(KEYINPUT67), .C1(new_n493_), .C2(new_n495_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n477_), .A2(new_n478_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(G99gat), .A2(G106gat), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT7), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n475_), .B(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n500_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT8), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT8), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n508_), .B(new_n500_), .C1(new_n503_), .C2(new_n505_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n498_), .A2(new_n499_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n435_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT34), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n514_), .A2(KEYINPUT35), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n512_), .B(new_n515_), .C1(new_n511_), .C2(new_n444_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(KEYINPUT35), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT68), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n516_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G190gat), .B(G218gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT70), .ZN(new_n521_));
  XOR2_X1   g320(.A(G134gat), .B(G162gat), .Z(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n519_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n519_), .A2(new_n524_), .A3(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT37), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n526_), .A2(KEYINPUT37), .A3(new_n527_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G57gat), .B(G64gat), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n533_), .A2(KEYINPUT11), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(KEYINPUT11), .ZN(new_n535_));
  XOR2_X1   g334(.A(G71gat), .B(G78gat), .Z(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n535_), .A2(new_n536_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G231gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n430_), .B(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G127gat), .B(G155gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G183gat), .B(G211gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT17), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n547_), .A2(KEYINPUT17), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n542_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n542_), .A2(new_n548_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554_));
  INV_X1    g353(.A(new_n539_), .ZN(new_n555_));
  NOR3_X1   g354(.A1(new_n483_), .A2(new_n484_), .A3(new_n482_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT64), .B1(new_n488_), .B2(new_n489_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n492_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n494_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n491_), .A2(KEYINPUT65), .A3(new_n492_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n480_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n510_), .B1(new_n561_), .B2(KEYINPUT67), .ZN(new_n562_));
  INV_X1    g361(.A(new_n499_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n555_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n498_), .A2(new_n499_), .A3(new_n510_), .A4(new_n539_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n554_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(KEYINPUT12), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT12), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n511_), .A2(new_n568_), .A3(new_n555_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n565_), .A2(new_n554_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n566_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G120gat), .B(G148gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT5), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G176gat), .B(G204gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n572_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n572_), .A2(new_n577_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT13), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n578_), .A2(KEYINPUT13), .A3(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n532_), .A2(new_n553_), .A3(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n471_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(new_n420_), .A3(new_n378_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT102), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n587_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n588_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  XNOR2_X1  g391(.A(new_n528_), .B(KEYINPUT100), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n419_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n468_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n584_), .A2(new_n595_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n594_), .A2(new_n552_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n420_), .B1(new_n597_), .B2(new_n378_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT101), .Z(new_n599_));
  NAND2_X1  g398(.A1(new_n592_), .A2(new_n599_), .ZN(G1324gat));
  NAND2_X1  g399(.A1(new_n597_), .A2(new_n344_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n601_), .A2(KEYINPUT104), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(KEYINPUT104), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(G8gat), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n602_), .A2(KEYINPUT39), .A3(G8gat), .A4(new_n603_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n586_), .A2(new_n421_), .A3(new_n344_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT103), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n606_), .A2(new_n607_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT40), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n606_), .A2(KEYINPUT40), .A3(new_n607_), .A4(new_n609_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(G1325gat));
  INV_X1    g413(.A(G15gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n597_), .B2(new_n395_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT105), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n617_), .A2(KEYINPUT41), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(KEYINPUT41), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n586_), .A2(new_n615_), .A3(new_n395_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .ZN(G1326gat));
  INV_X1    g420(.A(G22gat), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n597_), .B2(new_n272_), .ZN(new_n623_));
  XOR2_X1   g422(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n586_), .A2(new_n622_), .A3(new_n272_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1327gat));
  XOR2_X1   g426(.A(new_n528_), .B(KEYINPUT100), .Z(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n553_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(new_n584_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n471_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n631_), .A2(G29gat), .A3(new_n379_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n596_), .A2(new_n553_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n419_), .A2(new_n532_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT43), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n419_), .A2(new_n636_), .A3(new_n532_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n633_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT107), .B1(new_n638_), .B2(KEYINPUT44), .ZN(new_n639_));
  INV_X1    g438(.A(new_n633_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n419_), .A2(new_n636_), .A3(new_n532_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n636_), .B1(new_n419_), .B2(new_n532_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n640_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT107), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n639_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n638_), .A2(KEYINPUT44), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(new_n378_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n632_), .B1(new_n649_), .B2(G29gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT108), .ZN(G1328gat));
  INV_X1    g450(.A(new_n631_), .ZN(new_n652_));
  INV_X1    g451(.A(G36gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n653_), .A3(new_n344_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT45), .ZN(new_n655_));
  INV_X1    g454(.A(new_n344_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n638_), .B2(KEYINPUT44), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT109), .B(new_n653_), .C1(new_n647_), .C2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT109), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n638_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n644_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n657_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n659_), .B1(new_n662_), .B2(G36gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n655_), .B1(new_n658_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(KEYINPUT46), .B(new_n655_), .C1(new_n658_), .C2(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1329gat));
  INV_X1    g467(.A(new_n395_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n389_), .B1(new_n631_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n647_), .A2(new_n648_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n395_), .A2(G43gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g473(.A(G50gat), .B1(new_n652_), .B2(new_n272_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n671_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n272_), .A2(G50gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n675_), .B1(new_n676_), .B2(new_n677_), .ZN(G1331gat));
  AND2_X1   g477(.A1(new_n419_), .A2(new_n595_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n532_), .A2(new_n553_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(new_n584_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(G57gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n682_), .A3(new_n378_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n594_), .A2(new_n552_), .A3(new_n584_), .A4(new_n469_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G57gat), .B1(new_n684_), .B2(new_n379_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1332gat));
  OAI21_X1  g485(.A(G64gat), .B1(new_n684_), .B2(new_n656_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT48), .ZN(new_n688_));
  INV_X1    g487(.A(G64gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n681_), .A2(new_n689_), .A3(new_n344_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1333gat));
  OAI21_X1  g490(.A(G71gat), .B1(new_n684_), .B2(new_n669_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(G71gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n681_), .A2(new_n695_), .A3(new_n395_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1334gat));
  OAI21_X1  g496(.A(G78gat), .B1(new_n684_), .B2(new_n271_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT50), .ZN(new_n699_));
  INV_X1    g498(.A(G78gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n681_), .A2(new_n700_), .A3(new_n272_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1335gat));
  AND4_X1   g501(.A1(new_n628_), .A2(new_n679_), .A3(new_n553_), .A4(new_n584_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G85gat), .B1(new_n703_), .B2(new_n378_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT111), .Z(new_n705_));
  INV_X1    g504(.A(new_n584_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n706_), .A2(new_n552_), .A3(new_n468_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n641_), .A2(new_n642_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n709_), .A2(KEYINPUT112), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(KEYINPUT112), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n708_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n378_), .A2(G85gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n705_), .B1(new_n712_), .B2(new_n713_), .ZN(G1336gat));
  AOI21_X1  g513(.A(G92gat), .B1(new_n703_), .B2(new_n344_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n344_), .A2(new_n472_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n712_), .B2(new_n716_), .ZN(G1337gat));
  OR2_X1    g516(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n487_), .B1(new_n712_), .B2(new_n395_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n703_), .A2(new_n395_), .A3(new_n491_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(G1338gat));
  NAND2_X1  g523(.A1(new_n707_), .A2(new_n272_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G106gat), .B1(new_n709_), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT52), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n703_), .A2(new_n492_), .A3(new_n272_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g529(.A(KEYINPUT54), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n680_), .A2(new_n731_), .A3(new_n706_), .A4(new_n469_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n585_), .A2(new_n469_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT54), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n585_), .A2(KEYINPUT114), .A3(new_n731_), .A4(new_n469_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n734_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n451_), .A2(new_n455_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n462_), .A2(new_n447_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n436_), .A2(new_n441_), .A3(new_n447_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n456_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n580_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n466_), .B1(new_n465_), .B2(new_n443_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n443_), .ZN(new_n747_));
  AOI211_X1 g546(.A(new_n457_), .B(new_n747_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n579_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n496_), .A2(new_n497_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT12), .B(new_n539_), .C1(new_n750_), .C2(new_n499_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n568_), .B1(new_n511_), .B2(new_n555_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n565_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n554_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n571_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT55), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(new_n571_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n758_));
  AOI221_X4 g557(.A(KEYINPUT115), .B1(new_n753_), .B2(new_n754_), .C1(new_n756_), .C2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n756_), .A2(new_n758_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n753_), .A2(new_n754_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n576_), .B1(new_n759_), .B2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n749_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n757_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n758_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n762_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT115), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n761_), .A2(new_n760_), .A3(new_n762_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n577_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n765_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n745_), .B1(new_n767_), .B2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT117), .B1(new_n775_), .B2(new_n628_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n458_), .A2(new_n467_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n773_), .B2(new_n765_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n764_), .A2(new_n766_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n744_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n593_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n776_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT58), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n743_), .A2(new_n579_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(new_n764_), .B2(KEYINPUT56), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n773_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n773_), .A2(new_n788_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n764_), .A2(KEYINPUT56), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(KEYINPUT58), .A4(new_n786_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n532_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT118), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n790_), .A2(new_n796_), .A3(new_n532_), .A4(new_n793_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n780_), .A2(KEYINPUT57), .A3(new_n593_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n784_), .A2(new_n795_), .A3(new_n797_), .A4(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n738_), .B1(new_n799_), .B2(new_n553_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n669_), .A2(new_n379_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n345_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT59), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(G113gat), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n469_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n784_), .A2(new_n794_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n784_), .A2(KEYINPUT119), .A3(new_n794_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n798_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n738_), .B1(new_n810_), .B2(new_n553_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n802_), .A2(KEYINPUT59), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n803_), .B(new_n805_), .C1(new_n811_), .C2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n799_), .A2(new_n553_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n738_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n345_), .A3(new_n801_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n804_), .B1(new_n818_), .B2(new_n595_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n814_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n814_), .A2(KEYINPUT120), .A3(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1340gat));
  INV_X1    g623(.A(new_n818_), .ZN(new_n825_));
  INV_X1    g624(.A(G120gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n706_), .B2(KEYINPUT60), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n825_), .B(new_n827_), .C1(KEYINPUT60), .C2(new_n826_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n584_), .B(new_n803_), .C1(new_n811_), .C2(new_n813_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n828_), .B1(new_n830_), .B2(new_n826_), .ZN(G1341gat));
  INV_X1    g630(.A(G127gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n825_), .A2(new_n832_), .A3(new_n552_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n552_), .B(new_n803_), .C1(new_n811_), .C2(new_n813_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n835_), .B2(new_n832_), .ZN(G1342gat));
  AOI21_X1  g635(.A(G134gat), .B1(new_n825_), .B2(new_n628_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n811_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n838_), .A2(new_n812_), .B1(KEYINPUT59), .B2(new_n818_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n532_), .A2(G134gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT121), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n837_), .B1(new_n839_), .B2(new_n841_), .ZN(G1343gat));
  NOR2_X1   g641(.A1(new_n395_), .A2(new_n271_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n800_), .A2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n379_), .A2(new_n344_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT122), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  AND4_X1   g646(.A1(KEYINPUT122), .A2(new_n817_), .A3(new_n843_), .A4(new_n846_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n468_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G141gat), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n205_), .B(new_n468_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1344gat));
  OAI21_X1  g651(.A(new_n584_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(G148gat), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n206_), .B(new_n584_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1345gat));
  OAI21_X1  g655(.A(new_n552_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT61), .B(G155gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT123), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n857_), .A2(new_n860_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n552_), .B(new_n859_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1346gat));
  OR2_X1    g662(.A1(new_n847_), .A2(new_n848_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n532_), .A2(G162gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT124), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n628_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n867_));
  INV_X1    g666(.A(G162gat), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n864_), .A2(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(G1347gat));
  NAND2_X1  g668(.A1(new_n379_), .A2(new_n344_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n669_), .A2(new_n272_), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n798_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n552_), .B1(new_n873_), .B2(new_n809_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n468_), .B(new_n871_), .C1(new_n874_), .C2(new_n738_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G169gat), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n875_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n879_));
  INV_X1    g678(.A(new_n288_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n878_), .B(new_n879_), .C1(new_n880_), .C2(new_n875_), .ZN(G1348gat));
  NAND3_X1  g680(.A1(new_n838_), .A2(new_n584_), .A3(new_n871_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n817_), .A2(new_n871_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n706_), .A2(new_n289_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n882_), .A2(new_n289_), .B1(new_n883_), .B2(new_n884_), .ZN(G1349gat));
  AOI21_X1  g684(.A(new_n309_), .B1(new_n883_), .B2(new_n552_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n838_), .A2(new_n871_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n552_), .A2(new_n296_), .A3(new_n295_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n886_), .B1(new_n888_), .B2(new_n889_), .ZN(G1350gat));
  INV_X1    g689(.A(new_n532_), .ZN(new_n891_));
  OAI21_X1  g690(.A(G190gat), .B1(new_n887_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n628_), .A2(new_n292_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n887_), .B2(new_n893_), .ZN(G1351gat));
  NOR3_X1   g693(.A1(new_n800_), .A2(new_n844_), .A3(new_n870_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n468_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n584_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n899_));
  XOR2_X1   g698(.A(new_n899_), .B(KEYINPUT126), .Z(new_n900_));
  XOR2_X1   g699(.A(new_n898_), .B(new_n900_), .Z(G1353gat));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n902_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n895_), .A2(new_n552_), .A3(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n902_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n906_));
  XOR2_X1   g705(.A(new_n905_), .B(new_n906_), .Z(G1354gat));
  INV_X1    g706(.A(G218gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n895_), .A2(new_n908_), .A3(new_n628_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n895_), .A2(new_n532_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n908_), .ZN(G1355gat));
endmodule


