//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n571_, new_n572_, new_n573_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT23), .ZN(new_n206_));
  OR2_X1    g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT24), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(KEYINPUT24), .A3(new_n209_), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n204_), .A2(new_n206_), .A3(new_n208_), .A4(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT79), .B(G176gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT22), .B(G169gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(new_n209_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n216_), .A2(KEYINPUT88), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n206_), .B1(G183gat), .B2(G190gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(new_n216_), .B2(KEYINPUT88), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n211_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G197gat), .B(G204gat), .Z(new_n221_));
  OR2_X1    g020(.A1(new_n221_), .A2(KEYINPUT21), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(KEYINPUT21), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G211gat), .B(G218gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n225_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n215_), .A2(KEYINPUT80), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n218_), .B1(new_n215_), .B2(KEYINPUT80), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n211_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT81), .ZN(new_n231_));
  OAI211_X1 g030(.A(KEYINPUT20), .B(new_n227_), .C1(new_n231_), .C2(new_n226_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT89), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G226gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT19), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n232_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT20), .B1(new_n220_), .B2(new_n226_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n237_), .B1(new_n231_), .B2(new_n226_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n235_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n232_), .A2(new_n235_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT89), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G8gat), .B(G36gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT18), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G64gat), .B(G92gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n241_), .A2(new_n248_), .A3(new_n243_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT27), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n238_), .A2(new_n239_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(new_n235_), .B2(new_n232_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n256_), .B2(new_n249_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n251_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT2), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(G141gat), .A2(G148gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT84), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n263_), .B1(KEYINPUT3), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(KEYINPUT3), .B2(new_n265_), .ZN(new_n267_));
  XOR2_X1   g066(.A(G155gat), .B(G162gat), .Z(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n264_), .B(KEYINPUT83), .ZN(new_n272_));
  NAND3_X1  g071(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n261_), .A4(new_n273_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G113gat), .B(G120gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(G127gat), .B(G134gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n269_), .A2(new_n274_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT90), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G225gat), .A2(G233gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT90), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n280_), .A2(new_n288_), .A3(KEYINPUT4), .A4(new_n282_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n281_), .A2(new_n284_), .A3(new_n278_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n285_), .A2(new_n287_), .A3(new_n289_), .A4(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n280_), .A2(new_n286_), .A3(new_n282_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT91), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G1gat), .B(G29gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(G85gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT0), .B(G57gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n296_), .B(new_n297_), .Z(new_n298_));
  NAND3_X1  g097(.A1(new_n291_), .A2(new_n294_), .A3(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT97), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(KEYINPUT97), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n275_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G22gat), .B(G50gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n307_), .B(KEYINPUT28), .ZN(new_n312_));
  INV_X1    g111(.A(new_n310_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n314_), .A3(KEYINPUT87), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G78gat), .B(G106gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(KEYINPUT86), .Z(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n226_), .B1(new_n275_), .B2(new_n306_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G228gat), .A2(G233gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n320_), .B(KEYINPUT85), .Z(new_n321_));
  NOR2_X1   g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(KEYINPUT85), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(new_n319_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n315_), .A2(new_n318_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n318_), .B1(new_n315_), .B2(new_n324_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n311_), .A2(new_n314_), .ZN(new_n328_));
  OAI22_X1  g127(.A1(new_n326_), .A2(new_n327_), .B1(KEYINPUT87), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n327_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n328_), .A2(KEYINPUT87), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(new_n325_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n260_), .A2(new_n305_), .A3(new_n334_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n291_), .A2(new_n294_), .A3(KEYINPUT33), .A4(new_n298_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT92), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n285_), .A2(new_n286_), .A3(new_n289_), .A4(new_n290_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n298_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n338_), .B(new_n339_), .C1(new_n286_), .C2(new_n283_), .ZN(new_n340_));
  AND4_X1   g139(.A1(new_n337_), .A2(new_n340_), .A3(new_n251_), .A4(new_n250_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT93), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT33), .B1(new_n299_), .B2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(new_n342_), .B2(new_n299_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT94), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n343_), .B(KEYINPUT94), .C1(new_n342_), .C2(new_n299_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n248_), .A2(KEYINPUT32), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n302_), .A2(new_n303_), .B1(new_n350_), .B2(new_n256_), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n349_), .B(KEYINPUT95), .Z(new_n352_));
  NAND3_X1  g151(.A1(new_n241_), .A2(new_n243_), .A3(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n353_), .B(KEYINPUT96), .Z(new_n354_));
  AOI22_X1  g153(.A1(new_n341_), .A2(new_n348_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n335_), .B1(new_n355_), .B2(new_n334_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G71gat), .B(G99gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G43gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n231_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(new_n278_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G227gat), .A2(G233gat), .ZN(new_n361_));
  INV_X1    g160(.A(G15gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT30), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT31), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n360_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT82), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n260_), .A2(new_n305_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT98), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n260_), .A2(KEYINPUT98), .A3(new_n369_), .A4(new_n305_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n356_), .A2(new_n368_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G229gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G29gat), .B(G36gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G43gat), .B(G50gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT15), .ZN(new_n380_));
  INV_X1    g179(.A(G1gat), .ZN(new_n381_));
  INV_X1    g180(.A(G8gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G1gat), .A2(G8gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(G15gat), .A2(G22gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(G15gat), .A2(G22gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT14), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(G1gat), .B2(G8gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n385_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G15gat), .B(G22gat), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n392_), .A2(new_n389_), .A3(new_n384_), .A4(new_n383_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n380_), .A2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n377_), .A2(new_n378_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n377_), .A2(new_n378_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n391_), .B(new_n393_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT75), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n379_), .A2(KEYINPUT75), .A3(new_n391_), .A4(new_n393_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n376_), .B1(new_n395_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT76), .ZN(new_n404_));
  INV_X1    g203(.A(new_n379_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n394_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n402_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n403_), .B1(new_n409_), .B2(new_n376_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G113gat), .B(G141gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT77), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G169gat), .B(G197gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT78), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n402_), .A2(new_n406_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT76), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n402_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n376_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n395_), .A2(new_n402_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n375_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n414_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n416_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  AOI211_X1 g224(.A(KEYINPUT78), .B(new_n414_), .C1(new_n420_), .C2(new_n422_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n415_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G232gat), .A2(G233gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n429_), .B(KEYINPUT34), .Z(new_n430_));
  INV_X1    g229(.A(KEYINPUT35), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT7), .ZN(new_n433_));
  INV_X1    g232(.A(G99gat), .ZN(new_n434_));
  INV_X1    g233(.A(G106gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G99gat), .A2(G106gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT6), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(G99gat), .A3(G106gat), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT65), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT65), .B1(new_n440_), .B2(new_n442_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n438_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(G85gat), .A2(G92gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G85gat), .A2(G92gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n448_), .A2(KEYINPUT8), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n440_), .A2(new_n442_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n436_), .A2(new_n437_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n445_), .A2(new_n449_), .B1(new_n453_), .B2(KEYINPUT8), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n443_), .A2(new_n444_), .ZN(new_n455_));
  OR2_X1    g254(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n456_));
  NAND2_X1  g255(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n456_), .A2(G85gat), .A3(G92gat), .A4(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n446_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n447_), .ZN(new_n459_));
  OR2_X1    g258(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n435_), .A3(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n455_), .A2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT66), .B1(new_n454_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n440_), .A2(new_n442_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT65), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT65), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n452_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n449_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n448_), .B1(new_n438_), .B2(new_n466_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT8), .ZN(new_n473_));
  OAI22_X1  g272(.A1(new_n470_), .A2(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT66), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n455_), .A2(new_n463_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n465_), .A2(new_n380_), .A3(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(new_n379_), .A3(new_n476_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n430_), .A2(new_n431_), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n480_), .B(KEYINPUT69), .Z(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n481_), .A3(KEYINPUT70), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT70), .B1(new_n479_), .B2(new_n481_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n432_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n432_), .B(KEYINPUT71), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n478_), .A2(new_n479_), .A3(new_n481_), .A4(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT36), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G190gat), .B(G218gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(G134gat), .B(G162gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  NOR2_X1   g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n485_), .A2(new_n487_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n493_), .A3(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n497_), .B(KEYINPUT37), .Z(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n501_));
  XOR2_X1   g300(.A(G71gat), .B(G78gat), .Z(new_n502_));
  OR2_X1    g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n502_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n503_), .B(KEYINPUT12), .C1(new_n504_), .C2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n465_), .A2(new_n477_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT67), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n465_), .A2(new_n477_), .A3(KEYINPUT67), .A4(new_n507_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G230gat), .A2(G233gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n514_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n474_), .A2(new_n476_), .A3(new_n514_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(KEYINPUT12), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n512_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n513_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n516_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n521_), .B2(new_n515_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G120gat), .B(G148gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT5), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G176gat), .B(G204gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n525_), .B(new_n526_), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT68), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n523_), .B(new_n528_), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n529_), .A2(KEYINPUT13), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(KEYINPUT13), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G231gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n394_), .B(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(new_n514_), .Z(new_n535_));
  XOR2_X1   g334(.A(G127gat), .B(G155gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(G183gat), .B(G211gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n535_), .A2(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n543_), .B(KEYINPUT73), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n540_), .B(new_n541_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n544_), .B1(new_n535_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT74), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n499_), .A2(new_n532_), .A3(new_n547_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n374_), .A2(new_n428_), .A3(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(new_n381_), .A3(new_n304_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT38), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n547_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n497_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n374_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n532_), .A2(new_n427_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT99), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(G1gat), .B1(new_n558_), .B2(new_n305_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n550_), .A2(new_n551_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n552_), .A2(new_n559_), .A3(new_n560_), .ZN(G1324gat));
  NAND3_X1  g360(.A1(new_n555_), .A2(new_n259_), .A3(new_n557_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(G8gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT39), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n549_), .A2(new_n382_), .A3(new_n259_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT100), .Z(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n564_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(G1325gat));
  OAI21_X1  g369(.A(G15gat), .B1(new_n558_), .B2(new_n368_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT41), .Z(new_n572_));
  NAND3_X1  g371(.A1(new_n549_), .A2(new_n362_), .A3(new_n367_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(G1326gat));
  OAI21_X1  g373(.A(G22gat), .B1(new_n558_), .B2(new_n333_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT42), .ZN(new_n576_));
  INV_X1    g375(.A(G22gat), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n549_), .A2(new_n577_), .A3(new_n334_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(G1327gat));
  NOR2_X1   g378(.A1(new_n374_), .A2(new_n428_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n553_), .A2(new_n554_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n532_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(G29gat), .B1(new_n585_), .B2(new_n304_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT103), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n499_), .A2(KEYINPUT43), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n341_), .A2(new_n348_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n354_), .A2(new_n351_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n333_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n367_), .B1(new_n591_), .B2(new_n335_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n372_), .A2(new_n373_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n587_), .B(new_n588_), .C1(new_n592_), .C2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n498_), .B(KEYINPUT102), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT43), .B1(new_n374_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n588_), .ZN(new_n598_));
  OAI21_X1  g397(.A(KEYINPUT103), .B1(new_n374_), .B2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n595_), .A2(new_n597_), .A3(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n557_), .A2(new_n553_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n600_), .A2(KEYINPUT44), .A3(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT44), .B1(new_n600_), .B2(new_n601_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n304_), .A2(G29gat), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n586_), .B1(new_n604_), .B2(new_n605_), .ZN(G1328gat));
  NOR2_X1   g405(.A1(new_n260_), .A2(G36gat), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n580_), .A2(new_n583_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT104), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT104), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n580_), .A2(new_n610_), .A3(new_n583_), .A4(new_n607_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n609_), .A2(KEYINPUT45), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT45), .B1(new_n609_), .B2(new_n611_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n602_), .A2(new_n603_), .A3(new_n260_), .ZN(new_n615_));
  INV_X1    g414(.A(G36gat), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n614_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT46), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n614_), .B(KEYINPUT46), .C1(new_n615_), .C2(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1329gat));
  NAND2_X1  g420(.A1(new_n600_), .A2(new_n601_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT44), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n600_), .A2(KEYINPUT44), .A3(new_n601_), .ZN(new_n625_));
  INV_X1    g424(.A(G43gat), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n366_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n626_), .B1(new_n584_), .B2(new_n368_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(G1330gat));
  AOI21_X1  g431(.A(G50gat), .B1(new_n585_), .B2(new_n334_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n334_), .A2(G50gat), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n633_), .B1(new_n604_), .B2(new_n634_), .ZN(G1331gat));
  NAND3_X1  g434(.A1(new_n555_), .A2(new_n428_), .A3(new_n582_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G57gat), .B1(new_n636_), .B2(new_n305_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n374_), .A2(new_n427_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n638_), .A2(new_n582_), .A3(new_n547_), .A4(new_n499_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n305_), .A2(G57gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n637_), .B1(new_n639_), .B2(new_n640_), .ZN(G1332gat));
  OAI21_X1  g440(.A(G64gat), .B1(new_n636_), .B2(new_n260_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT48), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n260_), .A2(G64gat), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n643_), .B1(new_n639_), .B2(new_n644_), .ZN(G1333gat));
  OAI21_X1  g444(.A(G71gat), .B1(new_n636_), .B2(new_n368_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT49), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n368_), .A2(G71gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n639_), .B2(new_n648_), .ZN(G1334gat));
  OAI21_X1  g448(.A(G78gat), .B1(new_n636_), .B2(new_n333_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT50), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n333_), .A2(G78gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n651_), .B1(new_n639_), .B2(new_n652_), .ZN(G1335gat));
  NOR4_X1   g452(.A1(new_n374_), .A2(new_n427_), .A3(new_n532_), .A4(new_n581_), .ZN(new_n654_));
  INV_X1    g453(.A(G85gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n304_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n532_), .A2(new_n427_), .A3(new_n547_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n600_), .A2(new_n304_), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n656_), .B1(new_n658_), .B2(new_n655_), .ZN(G1336gat));
  AOI21_X1  g458(.A(G92gat), .B1(new_n654_), .B2(new_n259_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT106), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n600_), .A2(G92gat), .A3(new_n259_), .A4(new_n657_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1337gat));
  INV_X1    g462(.A(new_n366_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n654_), .A2(new_n664_), .A3(new_n460_), .A4(new_n461_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n600_), .A2(new_n367_), .A3(new_n657_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(new_n434_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g467(.A1(new_n654_), .A2(new_n435_), .A3(new_n334_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n600_), .A2(new_n334_), .A3(new_n657_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT52), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(G106gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n670_), .B2(G106gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT53), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT53), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n676_), .B(new_n669_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1339gat));
  XOR2_X1   g477(.A(KEYINPUT111), .B(KEYINPUT57), .Z(new_n679_));
  INV_X1    g478(.A(new_n527_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n519_), .A2(new_n522_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n427_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n512_), .A2(new_n518_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(KEYINPUT109), .A3(new_n520_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n517_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(new_n513_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n512_), .A2(KEYINPUT55), .A3(new_n513_), .A4(new_n518_), .ZN(new_n691_));
  AOI211_X1 g490(.A(new_n520_), .B(new_n517_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT108), .B(KEYINPUT55), .Z(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  OAI211_X1 g493(.A(KEYINPUT56), .B(new_n527_), .C1(new_n690_), .C2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n693_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n519_), .A2(new_n696_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n686_), .A2(new_n697_), .A3(new_n689_), .A4(new_n691_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT56), .B1(new_n698_), .B2(new_n527_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n699_), .B2(KEYINPUT110), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n527_), .B1(new_n690_), .B2(new_n694_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT56), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n701_), .A2(KEYINPUT110), .A3(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n684_), .B1(new_n700_), .B2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n409_), .A2(new_n376_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n414_), .B1(new_n421_), .B2(new_n375_), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n425_), .A2(new_n426_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n529_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n704_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n679_), .B1(new_n710_), .B2(new_n554_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT115), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT58), .ZN(new_n713_));
  INV_X1    g512(.A(new_n681_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n707_), .A2(new_n714_), .A3(KEYINPUT112), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT112), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n705_), .A2(new_n706_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT78), .B1(new_n410_), .B2(new_n414_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n423_), .A2(new_n416_), .A3(new_n424_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n716_), .B1(new_n720_), .B2(new_n681_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n715_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT113), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n695_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n701_), .A2(new_n702_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n701_), .A2(new_n723_), .A3(new_n702_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n722_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n713_), .B1(new_n728_), .B2(KEYINPUT114), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT114), .ZN(new_n730_));
  AOI211_X1 g529(.A(new_n730_), .B(new_n722_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n712_), .B(new_n498_), .C1(new_n729_), .C2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n728_), .A2(KEYINPUT58), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n715_), .A2(new_n721_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n699_), .B1(new_n723_), .B2(new_n695_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n727_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n730_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n728_), .A2(KEYINPUT114), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n713_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n712_), .B1(new_n741_), .B2(new_n498_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n711_), .B1(new_n734_), .B2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n709_), .A2(KEYINPUT57), .A3(new_n497_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT116), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n709_), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n497_), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n743_), .A2(KEYINPUT117), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT117), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n749_), .B(new_n711_), .C1(new_n734_), .C2(new_n742_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n547_), .B1(new_n748_), .B2(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n499_), .A2(new_n428_), .A3(new_n532_), .A4(new_n547_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT54), .Z(new_n753_));
  NOR2_X1   g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n260_), .A2(new_n304_), .A3(new_n369_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT59), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n746_), .A2(new_n747_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n758_), .B(new_n711_), .C1(new_n734_), .C2(new_n742_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n553_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n753_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n755_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  OAI22_X1  g563(.A1(new_n754_), .A2(new_n757_), .B1(new_n764_), .B2(new_n756_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G113gat), .B1(new_n765_), .B2(new_n428_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n428_), .A2(G113gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n763_), .B2(new_n767_), .ZN(G1340gat));
  OAI21_X1  g567(.A(G120gat), .B1(new_n765_), .B2(new_n532_), .ZN(new_n769_));
  INV_X1    g568(.A(G120gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n770_), .B1(new_n532_), .B2(KEYINPUT60), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(KEYINPUT60), .B2(new_n770_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n769_), .B1(new_n763_), .B2(new_n772_), .ZN(G1341gat));
  OAI21_X1  g572(.A(G127gat), .B1(new_n765_), .B2(new_n553_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n553_), .A2(G127gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n763_), .B2(new_n775_), .ZN(G1342gat));
  AOI21_X1  g575(.A(G134gat), .B1(new_n764_), .B2(new_n554_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n765_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(KEYINPUT118), .B(G134gat), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n499_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n777_), .B1(new_n778_), .B2(new_n780_), .ZN(G1343gat));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n367_), .A2(new_n333_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(new_n304_), .A3(new_n260_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n762_), .A2(new_n782_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n753_), .B1(new_n759_), .B2(new_n553_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT119), .B1(new_n787_), .B2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n427_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n582_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g592(.A(KEYINPUT120), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n789_), .B2(new_n547_), .ZN(new_n795_));
  AOI211_X1 g594(.A(KEYINPUT120), .B(new_n553_), .C1(new_n786_), .C2(new_n788_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT61), .B(G155gat), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n795_), .A2(new_n796_), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n782_), .B1(new_n762_), .B2(new_n785_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n787_), .A2(KEYINPUT119), .A3(new_n784_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n547_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT120), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n789_), .A2(new_n794_), .A3(new_n547_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n797_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n799_), .A2(new_n805_), .ZN(G1346gat));
  AOI21_X1  g605(.A(G162gat), .B1(new_n789_), .B2(new_n554_), .ZN(new_n807_));
  INV_X1    g606(.A(G162gat), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n596_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n789_), .B2(new_n809_), .ZN(G1347gat));
  NOR4_X1   g609(.A1(new_n368_), .A2(new_n260_), .A3(new_n304_), .A4(new_n334_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n427_), .B(new_n811_), .C1(new_n751_), .C2(new_n753_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G169gat), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT121), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(new_n815_), .A3(G169gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n814_), .A2(KEYINPUT62), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n213_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n812_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n815_), .B1(new_n812_), .B2(G169gat), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT62), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n817_), .A2(new_n822_), .ZN(G1348gat));
  INV_X1    g622(.A(new_n212_), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n751_), .A2(new_n753_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n825_), .A2(new_n811_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n824_), .B1(new_n826_), .B2(new_n582_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n762_), .A2(new_n811_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(G176gat), .A3(new_n582_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT122), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n827_), .A2(new_n830_), .ZN(G1349gat));
  AND2_X1   g630(.A1(new_n828_), .A2(new_n547_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n832_), .A2(G183gat), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n553_), .A2(new_n202_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n825_), .A2(new_n811_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT123), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n825_), .A2(new_n837_), .A3(new_n811_), .A4(new_n834_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n833_), .A2(new_n836_), .A3(new_n838_), .ZN(G1350gat));
  NAND3_X1  g638(.A1(new_n826_), .A2(new_n203_), .A3(new_n554_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT124), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n498_), .B(new_n811_), .C1(new_n751_), .C2(new_n753_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(G190gat), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n842_), .A2(new_n841_), .A3(G190gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n840_), .B1(new_n843_), .B2(new_n844_), .ZN(G1351gat));
  NAND2_X1  g644(.A1(new_n783_), .A2(new_n305_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n259_), .B1(new_n846_), .B2(KEYINPUT125), .ZN(new_n847_));
  AOI211_X1 g646(.A(new_n847_), .B(new_n787_), .C1(KEYINPUT125), .C2(new_n846_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n427_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT126), .B(G197gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n849_), .B2(new_n852_), .ZN(G1352gat));
  INV_X1    g652(.A(G204gat), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n848_), .B(new_n582_), .C1(KEYINPUT127), .C2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(KEYINPUT127), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1353gat));
  NAND2_X1  g656(.A1(new_n848_), .A2(new_n547_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n859_));
  AND2_X1   g658(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n858_), .B2(new_n859_), .ZN(G1354gat));
  INV_X1    g661(.A(G218gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n848_), .A2(new_n863_), .A3(new_n554_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n848_), .A2(new_n498_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n863_), .ZN(G1355gat));
endmodule


