//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n955_, new_n956_, new_n957_, new_n959_, new_n960_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n975_;
  OR2_X1    g000(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(KEYINPUT9), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n205_), .A2(new_n208_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n206_), .A2(new_n207_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR3_X1   g017(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  AOI211_X1 g019(.A(KEYINPUT8), .B(new_n216_), .C1(new_n220_), .C2(new_n213_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT8), .ZN(new_n222_));
  OR3_X1    g021(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n211_), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n223_), .B(new_n217_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n216_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n222_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n215_), .B1(new_n221_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G29gat), .B(G36gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G43gat), .B(G50gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT15), .ZN(new_n235_));
  OAI211_X1 g034(.A(KEYINPUT65), .B(new_n215_), .C1(new_n221_), .C2(new_n228_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n231_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G232gat), .A2(G233gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n238_), .B(KEYINPUT34), .Z(new_n239_));
  INV_X1    g038(.A(KEYINPUT35), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT70), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n240_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT71), .ZN(new_n244_));
  INV_X1    g043(.A(new_n215_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n228_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n226_), .A2(new_n222_), .A3(new_n227_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n245_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n244_), .B1(new_n248_), .B2(new_n234_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n237_), .A2(new_n242_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT72), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT72), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n237_), .A2(new_n249_), .A3(new_n252_), .A4(new_n242_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n237_), .A2(new_n249_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n242_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT75), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G190gat), .B(G218gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G134gat), .B(G162gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n262_), .B(KEYINPUT36), .Z(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT74), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n258_), .A2(new_n259_), .A3(new_n264_), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n251_), .A2(new_n253_), .B1(new_n256_), .B2(new_n255_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n264_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT75), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n242_), .B1(new_n237_), .B2(new_n249_), .ZN(new_n269_));
  NOR3_X1   g068(.A1(new_n269_), .A2(KEYINPUT36), .A3(new_n262_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT73), .B1(new_n254_), .B2(new_n270_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n254_), .A2(new_n270_), .A3(KEYINPUT73), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n265_), .B(new_n268_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT76), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n274_), .A3(KEYINPUT37), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n272_), .A2(new_n271_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT37), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n258_), .A2(new_n263_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n274_), .B1(new_n273_), .B2(KEYINPUT37), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G57gat), .B(G64gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G71gat), .B(G78gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(KEYINPUT11), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(KEYINPUT11), .ZN(new_n286_));
  INV_X1    g085(.A(new_n284_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n283_), .A2(KEYINPUT11), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n285_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G231gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(KEYINPUT77), .B(G1gat), .Z(new_n293_));
  INV_X1    g092(.A(G8gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT14), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G15gat), .B(G22gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n295_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n292_), .B(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G127gat), .B(G155gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT16), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G183gat), .B(G211gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT17), .B1(new_n304_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT78), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n304_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  OAI211_X1 g111(.A(KEYINPUT17), .B(new_n308_), .C1(new_n304_), .C2(new_n310_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n282_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT79), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n316_), .A2(KEYINPUT79), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G230gat), .ZN(new_n321_));
  INV_X1    g120(.A(G233gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n290_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n229_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT64), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n290_), .B(new_n215_), .C1(new_n221_), .C2(new_n228_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n327_), .A2(new_n326_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n323_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n231_), .A2(KEYINPUT12), .A3(new_n324_), .A4(new_n236_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n327_), .A2(KEYINPUT12), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n325_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n323_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n331_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G120gat), .B(G148gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G176gat), .B(G204gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n330_), .A2(new_n335_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT68), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n330_), .A2(new_n335_), .A3(KEYINPUT68), .A4(new_n340_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n340_), .B(KEYINPUT67), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(new_n330_), .B2(new_n335_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n345_), .A2(KEYINPUT69), .A3(new_n348_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(KEYINPUT13), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT13), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT69), .B1(new_n345_), .B2(new_n348_), .ZN(new_n355_));
  AOI211_X1 g154(.A(new_n350_), .B(new_n347_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n354_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n353_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G78gat), .B(G106gat), .ZN(new_n359_));
  INV_X1    g158(.A(G228gat), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n360_), .A2(new_n322_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT21), .ZN(new_n363_));
  AND2_X1   g162(.A1(G197gat), .A2(G204gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(G197gat), .A2(G204gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(G197gat), .ZN(new_n367_));
  INV_X1    g166(.A(G204gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G197gat), .A2(G204gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(KEYINPUT21), .A3(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G211gat), .B(G218gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n366_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(G218gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(G211gat), .ZN(new_n375_));
  INV_X1    g174(.A(G211gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(G218gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n378_), .A2(KEYINPUT21), .A3(new_n369_), .A4(new_n370_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT88), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n373_), .A2(new_n379_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  OR2_X1    g183(.A1(G155gat), .A2(G162gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G141gat), .A2(G148gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT86), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(G141gat), .A3(G148gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT2), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n390_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n395_));
  INV_X1    g194(.A(G141gat), .ZN(new_n396_));
  INV_X1    g195(.A(G148gat), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .A4(KEYINPUT87), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT87), .ZN(new_n399_));
  OAI22_X1  g198(.A1(new_n399_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n398_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n388_), .B1(new_n394_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n396_), .A2(new_n397_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n405_));
  AND4_X1   g204(.A1(new_n390_), .A2(new_n392_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT1), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n385_), .A2(new_n407_), .A3(new_n386_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n403_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT29), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n362_), .B1(new_n384_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n380_), .A2(new_n362_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(KEYINPUT29), .B2(new_n410_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n359_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n359_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n413_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n411_), .A2(new_n417_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n381_), .A2(new_n383_), .B1(new_n410_), .B2(KEYINPUT29), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n416_), .B(new_n418_), .C1(new_n419_), .C2(new_n362_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT89), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n418_), .B1(new_n419_), .B2(new_n362_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n422_), .B1(new_n423_), .B2(new_n359_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n410_), .A2(KEYINPUT29), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G22gat), .B(G50gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT28), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n425_), .B(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n421_), .B1(new_n424_), .B2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n415_), .A2(new_n422_), .A3(new_n428_), .A4(new_n420_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433_));
  OAI21_X1  g232(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G183gat), .A2(G190gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT23), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT23), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(G183gat), .A3(G190gat), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(G183gat), .A2(G190gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n437_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  OR2_X1    g243(.A1(G169gat), .A2(G176gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G169gat), .A2(G176gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(KEYINPUT24), .A3(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G169gat), .A2(G176gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT24), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(KEYINPUT81), .A2(G183gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT25), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT25), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(KEYINPUT81), .A3(G183gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G190gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT26), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT26), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(G190gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n447_), .B(new_n450_), .C1(new_n455_), .C2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n441_), .A2(KEYINPUT82), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT82), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n463_), .A2(new_n440_), .A3(G183gat), .A4(G190gat), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n462_), .A2(new_n464_), .B1(KEYINPUT23), .B2(new_n438_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n444_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT20), .B1(new_n466_), .B2(new_n380_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n373_), .A2(new_n379_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n458_), .A2(G190gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n456_), .A2(KEYINPUT26), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT25), .B(G183gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n457_), .A2(new_n459_), .A3(KEYINPUT91), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n476_));
  NOR2_X1   g275(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n445_), .B(new_n446_), .C1(new_n476_), .C2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n476_), .A2(new_n477_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n479_), .A2(new_n448_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n475_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n437_), .B1(new_n465_), .B2(new_n443_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n468_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G226gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n467_), .A2(new_n483_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT20), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(new_n466_), .B2(new_n380_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n481_), .A2(new_n482_), .A3(new_n468_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n488_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G8gat), .B(G36gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(G64gat), .B(G92gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n487_), .A2(new_n492_), .A3(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n490_), .A2(new_n491_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n486_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n481_), .A2(new_n482_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n380_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n461_), .A2(new_n465_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(new_n444_), .A3(new_n468_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n503_), .A2(KEYINPUT20), .A3(new_n505_), .A4(new_n488_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n497_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n433_), .B1(new_n499_), .B2(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n467_), .A2(new_n483_), .A3(new_n488_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n381_), .A2(new_n383_), .A3(new_n481_), .A4(new_n482_), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT95), .B(KEYINPUT20), .Z(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n466_), .B2(new_n380_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n486_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n497_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n498_), .B1(new_n487_), .B2(new_n492_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT27), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n432_), .A2(new_n508_), .A3(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n398_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n390_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n387_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n390_), .A2(new_n392_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n407_), .B2(new_n388_), .ZN(new_n522_));
  INV_X1    g321(.A(G134gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(G127gat), .ZN(new_n524_));
  INV_X1    g323(.A(G127gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(G134gat), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT85), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n524_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n527_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G113gat), .B(G120gat), .Z(new_n530_));
  NOR3_X1   g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G113gat), .B(G120gat), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n525_), .A2(G134gat), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n523_), .A2(G127gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT85), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n524_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n532_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  OAI22_X1  g336(.A1(new_n520_), .A2(new_n522_), .B1(new_n531_), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n530_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(new_n536_), .A3(new_n532_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n403_), .A2(new_n539_), .A3(new_n409_), .A4(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(KEYINPUT4), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G225gat), .A2(G233gat), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT4), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n540_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n410_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n538_), .A2(new_n541_), .A3(new_n543_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G1gat), .B(G29gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(G85gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT0), .B(G57gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n554_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n548_), .A2(new_n549_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n504_), .A2(KEYINPUT30), .A3(new_n444_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n466_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT84), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n560_), .A2(KEYINPUT84), .A3(new_n562_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G227gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(G15gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT83), .B(G43gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G71gat), .B(G99gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n567_), .A2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT84), .B1(new_n560_), .B2(new_n562_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n546_), .B(KEYINPUT31), .Z(new_n579_));
  NAND3_X1  g378(.A1(new_n575_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n579_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n573_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n581_), .B1(new_n582_), .B2(new_n577_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n559_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT98), .B1(new_n517_), .B2(new_n584_), .ZN(new_n585_));
  AND4_X1   g384(.A1(new_n580_), .A2(new_n583_), .A3(new_n557_), .A4(new_n555_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n507_), .A2(new_n433_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n501_), .A2(new_n506_), .A3(new_n497_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n515_), .A2(new_n589_), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n588_), .A2(new_n514_), .B1(new_n590_), .B2(new_n433_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n586_), .A2(new_n587_), .A3(new_n432_), .A4(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n585_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n580_), .A2(new_n583_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n519_), .A2(new_n398_), .A3(new_n401_), .A4(new_n400_), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n595_), .A2(new_n388_), .B1(new_n408_), .B2(new_n406_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT29), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n373_), .A2(new_n382_), .A3(new_n379_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n382_), .B1(new_n373_), .B2(new_n379_), .ZN(new_n599_));
  OAI22_X1  g398(.A1(new_n596_), .A2(new_n597_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n600_), .A2(new_n361_), .B1(new_n411_), .B2(new_n417_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT89), .B1(new_n601_), .B2(new_n416_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n602_), .A2(new_n428_), .B1(new_n415_), .B2(new_n420_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n431_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT32), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n497_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n501_), .A2(new_n506_), .ZN(new_n609_));
  AOI22_X1  g408(.A1(new_n555_), .A2(new_n557_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n607_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI211_X1 g412(.A(KEYINPUT96), .B(new_n607_), .C1(new_n509_), .C2(new_n513_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n610_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n499_), .A2(new_n507_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n542_), .A2(new_n543_), .A3(new_n547_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT94), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n542_), .A2(new_n620_), .A3(new_n543_), .A4(new_n547_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n538_), .A2(new_n541_), .A3(new_n544_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n622_), .A2(new_n554_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(new_n621_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n557_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n548_), .A2(KEYINPUT33), .A3(new_n549_), .A4(new_n556_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n617_), .A2(new_n624_), .A3(new_n626_), .A4(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n605_), .B1(new_n616_), .B2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n508_), .A2(new_n430_), .A3(new_n431_), .A4(new_n516_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n630_), .A2(new_n558_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n594_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT97), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n634_), .B(new_n594_), .C1(new_n629_), .C2(new_n631_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n593_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n302_), .B(new_n234_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G229gat), .A2(G233gat), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n235_), .A2(new_n301_), .A3(new_n300_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n302_), .A2(new_n234_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n638_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G113gat), .B(G141gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G169gat), .B(G197gat), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n645_), .B(new_n646_), .Z(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n644_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n640_), .A2(new_n643_), .A3(new_n647_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT80), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n649_), .A2(KEYINPUT80), .A3(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT99), .B1(new_n636_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n585_), .A2(new_n592_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n635_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n591_), .A2(new_n605_), .A3(new_n559_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n619_), .A2(new_n621_), .A3(new_n623_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(new_n590_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n626_), .A2(new_n627_), .ZN(new_n663_));
  AOI22_X1  g462(.A1(new_n662_), .A2(new_n663_), .B1(new_n610_), .B2(new_n615_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n660_), .B1(new_n664_), .B2(new_n605_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n634_), .B1(new_n665_), .B2(new_n594_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n658_), .B1(new_n659_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n655_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n358_), .B1(new_n657_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n320_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n320_), .A2(KEYINPUT100), .A3(new_n671_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n558_), .A2(new_n293_), .ZN(new_n677_));
  XOR2_X1   g476(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n678_));
  NAND3_X1  g477(.A1(new_n676_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n276_), .A2(new_n278_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n667_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n353_), .A2(new_n357_), .A3(new_n655_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT102), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n353_), .A2(new_n357_), .A3(new_n686_), .A4(new_n655_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n683_), .A2(new_n314_), .A3(new_n685_), .A4(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G1gat), .B1(new_n688_), .B2(new_n559_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n679_), .A2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n678_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1324gat));
  INV_X1    g491(.A(KEYINPUT40), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n688_), .A2(new_n591_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G8gat), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n697_), .A2(KEYINPUT39), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n694_), .A2(KEYINPUT103), .A3(G8gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n697_), .A2(KEYINPUT39), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  NOR4_X1   g500(.A1(new_n674_), .A2(new_n675_), .A3(G8gat), .A4(new_n591_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n693_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n591_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n676_), .A2(new_n294_), .A3(new_n704_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n705_), .A2(KEYINPUT40), .A3(new_n698_), .A4(new_n700_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(G1325gat));
  OAI21_X1  g506(.A(G15gat), .B1(new_n688_), .B2(new_n594_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT41), .Z(new_n709_));
  INV_X1    g508(.A(G15gat), .ZN(new_n710_));
  INV_X1    g509(.A(new_n594_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n672_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(G1326gat));
  OAI21_X1  g512(.A(G22gat), .B1(new_n688_), .B2(new_n432_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT42), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n432_), .A2(G22gat), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT104), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n672_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1327gat));
  NAND2_X1  g518(.A1(new_n680_), .A2(new_n315_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n671_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G29gat), .B1(new_n721_), .B2(new_n558_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n685_), .A2(new_n315_), .A3(new_n687_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n273_), .A2(KEYINPUT37), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT76), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n279_), .A3(new_n275_), .ZN(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT43), .B1(new_n726_), .B2(new_n636_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n282_), .A2(new_n667_), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n723_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(KEYINPUT44), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n729_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n723_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(KEYINPUT44), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT105), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n730_), .A2(new_n736_), .A3(KEYINPUT44), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n731_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n558_), .A2(G29gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n722_), .B1(new_n738_), .B2(new_n739_), .ZN(G1328gat));
  INV_X1    g539(.A(G36gat), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n735_), .A2(new_n737_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n704_), .B1(new_n730_), .B2(KEYINPUT44), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n741_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n720_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n591_), .A2(G36gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n670_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT45), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n670_), .A2(new_n750_), .A3(new_n746_), .A4(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT106), .B1(new_n745_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n743_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n756_), .B(new_n752_), .C1(new_n757_), .C2(new_n741_), .ZN(new_n758_));
  AND4_X1   g557(.A1(KEYINPUT107), .A2(new_n754_), .A3(new_n755_), .A4(new_n758_), .ZN(new_n759_));
  OAI211_X1 g558(.A(KEYINPUT46), .B(new_n752_), .C1(new_n757_), .C2(new_n741_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n752_), .B1(new_n757_), .B2(new_n741_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT46), .B1(new_n763_), .B2(KEYINPUT106), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n762_), .B1(new_n764_), .B2(new_n758_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n759_), .A2(new_n765_), .ZN(G1329gat));
  AND3_X1   g565(.A1(new_n738_), .A2(G43gat), .A3(new_n711_), .ZN(new_n767_));
  AOI21_X1  g566(.A(G43gat), .B1(new_n721_), .B2(new_n711_), .ZN(new_n768_));
  OR3_X1    g567(.A1(new_n767_), .A2(KEYINPUT47), .A3(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT47), .B1(new_n767_), .B2(new_n768_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1330gat));
  INV_X1    g570(.A(new_n738_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G50gat), .B1(new_n772_), .B2(new_n432_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n432_), .A2(G50gat), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT108), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n721_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(G1331gat));
  NAND4_X1  g576(.A1(new_n683_), .A2(new_n314_), .A3(new_n358_), .A4(new_n656_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G57gat), .B1(new_n778_), .B2(new_n559_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n358_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n636_), .A2(new_n780_), .A3(new_n655_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n559_), .A2(G57gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(G1332gat));
  OAI21_X1  g583(.A(G64gat), .B1(new_n778_), .B2(new_n591_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT48), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n591_), .A2(G64gat), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT109), .Z(new_n788_));
  OAI21_X1  g587(.A(new_n786_), .B1(new_n782_), .B2(new_n788_), .ZN(G1333gat));
  OAI21_X1  g588(.A(G71gat), .B1(new_n778_), .B2(new_n594_), .ZN(new_n790_));
  XOR2_X1   g589(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n791_));
  XNOR2_X1  g590(.A(new_n790_), .B(new_n791_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n594_), .A2(G71gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n782_), .B2(new_n793_), .ZN(G1334gat));
  OAI21_X1  g593(.A(G78gat), .B1(new_n778_), .B2(new_n432_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT50), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n432_), .A2(G78gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n782_), .B2(new_n797_), .ZN(G1335gat));
  INV_X1    g597(.A(new_n732_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n358_), .A2(new_n315_), .A3(new_n656_), .ZN(new_n800_));
  OR2_X1    g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(G85gat), .B1(new_n801_), .B2(new_n559_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n781_), .A2(new_n746_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(G85gat), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n558_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n802_), .A2(new_n807_), .ZN(G1336gat));
  AOI21_X1  g607(.A(G92gat), .B1(new_n805_), .B2(new_n704_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n801_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n704_), .A2(G92gat), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT112), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n809_), .B1(new_n810_), .B2(new_n812_), .ZN(G1337gat));
  OAI21_X1  g612(.A(G99gat), .B1(new_n801_), .B2(new_n594_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT113), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n805_), .A2(new_n202_), .A3(new_n204_), .A4(new_n711_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT51), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n815_), .A2(new_n819_), .A3(new_n816_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(G1338gat));
  OAI21_X1  g620(.A(G106gat), .B1(new_n801_), .B2(new_n432_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT52), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n432_), .A2(G106gat), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT114), .B1(new_n805_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n805_), .A2(KEYINPUT114), .A3(new_n824_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n823_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT53), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n823_), .A2(new_n831_), .A3(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1339gat));
  NAND4_X1  g632(.A1(new_n726_), .A2(new_n314_), .A3(new_n780_), .A4(new_n656_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n834_), .B(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n335_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n335_), .B2(new_n837_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n334_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n840_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT56), .B1(new_n843_), .B2(new_n346_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845_));
  INV_X1    g644(.A(new_n346_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n841_), .A2(new_n842_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n845_), .B(new_n846_), .C1(new_n847_), .C2(new_n840_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n637_), .A2(new_n638_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n641_), .A2(new_n642_), .A3(new_n639_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n648_), .A3(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n650_), .A2(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n844_), .A2(new_n848_), .A3(new_n345_), .A4(new_n852_), .ZN(new_n853_));
  XOR2_X1   g652(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT118), .B1(new_n726_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n853_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n280_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n725_), .A4(new_n855_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n857_), .A2(new_n859_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT119), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n857_), .A2(new_n862_), .A3(new_n865_), .A4(new_n859_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n844_), .A2(new_n655_), .A3(new_n848_), .A4(new_n345_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n852_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n680_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  AND2_X1   g668(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n869_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n864_), .A2(new_n866_), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n836_), .B1(new_n876_), .B2(new_n315_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n517_), .A2(new_n594_), .A3(new_n559_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n877_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(G113gat), .B1(new_n880_), .B2(new_n655_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n836_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n875_), .A2(new_n863_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n314_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n878_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n880_), .B2(new_n885_), .ZN(new_n889_));
  OAI211_X1 g688(.A(KEYINPUT121), .B(KEYINPUT59), .C1(new_n877_), .C2(new_n879_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n887_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n655_), .A2(G113gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n881_), .B1(new_n891_), .B2(new_n892_), .ZN(G1340gat));
  INV_X1    g692(.A(G120gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n894_), .B1(new_n780_), .B2(KEYINPUT60), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n880_), .B(new_n895_), .C1(KEYINPUT60), .C2(new_n894_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n886_), .A2(new_n358_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n898_), .B2(new_n894_), .ZN(G1341gat));
  AOI21_X1  g698(.A(G127gat), .B1(new_n880_), .B2(new_n314_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n315_), .A2(new_n525_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n891_), .B2(new_n901_), .ZN(G1342gat));
  AOI21_X1  g701(.A(new_n874_), .B1(new_n863_), .B2(KEYINPUT119), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n314_), .B1(new_n903_), .B2(new_n866_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n680_), .B(new_n878_), .C1(new_n904_), .C2(new_n836_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n523_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n905_), .A2(KEYINPUT122), .A3(new_n523_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  XOR2_X1   g709(.A(KEYINPUT123), .B(G134gat), .Z(new_n911_));
  NOR2_X1   g710(.A1(new_n726_), .A2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n891_), .B2(new_n912_), .ZN(G1343gat));
  NOR2_X1   g712(.A1(new_n630_), .A2(new_n559_), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n594_), .B(new_n914_), .C1(new_n904_), .C2(new_n836_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n656_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n396_), .ZN(G1344gat));
  NOR2_X1   g716(.A1(new_n915_), .A2(new_n780_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(new_n397_), .ZN(G1345gat));
  NAND2_X1  g718(.A1(new_n876_), .A2(new_n315_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n711_), .B1(new_n920_), .B2(new_n882_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n921_), .A2(KEYINPUT124), .A3(new_n314_), .A4(new_n914_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n923_), .B1(new_n915_), .B2(new_n315_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT61), .B(G155gat), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n922_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n922_), .B2(new_n924_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1346gat));
  OAI21_X1  g727(.A(G162gat), .B1(new_n915_), .B2(new_n726_), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n681_), .A2(G162gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n915_), .B2(new_n930_), .ZN(G1347gat));
  NAND2_X1  g730(.A1(new_n884_), .A2(new_n432_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n584_), .A2(new_n591_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n656_), .A2(new_n935_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT22), .B(G169gat), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n933_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  XOR2_X1   g737(.A(new_n936_), .B(KEYINPUT125), .Z(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(new_n940_));
  OAI21_X1  g739(.A(G169gat), .B1(new_n932_), .B2(new_n940_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n941_), .A2(KEYINPUT62), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(KEYINPUT62), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n938_), .B1(new_n942_), .B2(new_n943_), .ZN(G1348gat));
  NAND3_X1  g743(.A1(new_n884_), .A2(new_n432_), .A3(new_n934_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(G176gat), .B1(new_n946_), .B2(new_n358_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n877_), .A2(new_n605_), .ZN(new_n948_));
  AND3_X1   g747(.A1(new_n358_), .A2(G176gat), .A3(new_n934_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n948_), .A2(KEYINPUT126), .A3(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n948_), .A2(new_n949_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n947_), .B1(new_n950_), .B2(new_n953_), .ZN(G1349gat));
  NOR2_X1   g753(.A1(new_n935_), .A2(new_n315_), .ZN(new_n955_));
  AOI21_X1  g754(.A(G183gat), .B1(new_n948_), .B2(new_n955_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n935_), .A2(new_n315_), .A3(new_n473_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n956_), .B1(new_n933_), .B2(new_n957_), .ZN(G1350gat));
  OAI21_X1  g757(.A(G190gat), .B1(new_n945_), .B2(new_n726_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n680_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n945_), .B2(new_n960_), .ZN(G1351gat));
  NOR3_X1   g760(.A1(new_n591_), .A2(new_n432_), .A3(new_n558_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n921_), .A2(new_n962_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n963_), .A2(new_n656_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n964_), .B(new_n367_), .ZN(G1352gat));
  NOR2_X1   g764(.A1(new_n963_), .A2(new_n780_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(new_n368_), .ZN(G1353gat));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n314_), .B1(new_n968_), .B2(new_n376_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n963_), .A2(new_n969_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n968_), .A2(new_n376_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(KEYINPUT127), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n970_), .B(new_n972_), .ZN(G1354gat));
  OAI21_X1  g772(.A(G218gat), .B1(new_n963_), .B2(new_n726_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n680_), .A2(new_n374_), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n974_), .B1(new_n963_), .B2(new_n975_), .ZN(G1355gat));
endmodule


