//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_;
  XNOR2_X1  g000(.A(KEYINPUT85), .B(G127gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G134gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(G113gat), .B(G120gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G134gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n202_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n204_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n205_), .A2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT89), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT88), .ZN(new_n217_));
  INV_X1    g016(.A(G141gat), .ZN(new_n218_));
  INV_X1    g017(.A(G148gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n216_), .A2(KEYINPUT88), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n217_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(KEYINPUT88), .B(new_n216_), .C1(new_n218_), .C2(new_n219_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n222_), .A2(new_n223_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT87), .ZN(new_n229_));
  OR3_X1    g028(.A1(new_n212_), .A2(new_n229_), .A3(KEYINPUT1), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n229_), .B1(new_n212_), .B2(KEYINPUT1), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n230_), .A2(new_n211_), .A3(new_n231_), .A4(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n220_), .A2(new_n224_), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n215_), .A2(new_n228_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n210_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n210_), .A2(new_n235_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(KEYINPUT4), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G225gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT96), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n236_), .A2(KEYINPUT97), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT97), .B1(new_n236_), .B2(new_n242_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n239_), .B(new_n241_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n237_), .A2(new_n238_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n240_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G85gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G1gat), .B(G29gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT99), .B(G57gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(new_n253_), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n248_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n245_), .A2(new_n247_), .A3(new_n254_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n235_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G22gat), .B(G50gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n261_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n235_), .A2(new_n259_), .A3(new_n264_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n262_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n263_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G78gat), .B(G106gat), .Z(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G228gat), .A2(G233gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT91), .Z(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(KEYINPUT21), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT21), .ZN(new_n276_));
  XOR2_X1   g075(.A(G197gat), .B(G204gat), .Z(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n276_), .A2(new_n277_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(new_n235_), .B2(new_n259_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT92), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  OAI211_X1 g082(.A(KEYINPUT92), .B(new_n280_), .C1(new_n235_), .C2(new_n259_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n273_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n284_), .A2(new_n273_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n270_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n285_), .A2(new_n270_), .A3(new_n286_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n268_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT93), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n285_), .A2(new_n286_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n269_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n287_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(KEYINPUT93), .A3(new_n268_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n289_), .A2(KEYINPUT94), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n298_), .B1(new_n295_), .B2(KEYINPUT94), .ZN(new_n299_));
  INV_X1    g098(.A(new_n268_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n258_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G226gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT19), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT24), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307_));
  MUX2_X1   g106(.A(new_n306_), .B(KEYINPUT24), .S(new_n307_), .Z(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT26), .B(G190gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT25), .B(G183gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(G183gat), .B2(G190gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT83), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AOI211_X1 g114(.A(KEYINPUT83), .B(new_n312_), .C1(G183gat), .C2(G190gat), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G183gat), .ZN(new_n318_));
  INV_X1    g117(.A(G190gat), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n318_), .A2(new_n319_), .A3(KEYINPUT23), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n308_), .B(new_n311_), .C1(new_n317_), .C2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n305_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT22), .B(G169gat), .ZN(new_n323_));
  INV_X1    g122(.A(G176gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n322_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n313_), .A2(KEYINPUT84), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n313_), .A2(KEYINPUT84), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n320_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n325_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n321_), .A2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT20), .B1(new_n331_), .B2(new_n280_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n280_), .ZN(new_n333_));
  OR3_X1    g132(.A1(new_n326_), .A2(new_n327_), .A3(new_n320_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n309_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n310_), .B(KEYINPUT95), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n334_), .B(new_n308_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n315_), .A2(new_n316_), .A3(new_n320_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n325_), .B1(new_n338_), .B2(new_n329_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n333_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n304_), .B1(new_n332_), .B2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT18), .B(G64gat), .ZN(new_n342_));
  INV_X1    g141(.A(G92gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G8gat), .B(G36gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT20), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(new_n331_), .B2(new_n280_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n304_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n337_), .A2(new_n333_), .A3(new_n339_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n341_), .A2(new_n346_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n332_), .A2(new_n340_), .A3(new_n304_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n337_), .A2(new_n339_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT101), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n348_), .B1(new_n357_), .B2(new_n280_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n354_), .B1(new_n358_), .B2(new_n304_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n346_), .B(KEYINPUT102), .ZN(new_n360_));
  OAI211_X1 g159(.A(KEYINPUT27), .B(new_n353_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n346_), .B1(new_n341_), .B2(new_n351_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n352_), .A2(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n363_), .A2(KEYINPUT27), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n302_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n355_), .A2(new_n356_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT101), .B1(new_n337_), .B2(new_n339_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n280_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n348_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n304_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n341_), .A2(KEYINPUT100), .A3(new_n351_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n354_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n346_), .A2(KEYINPUT32), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT100), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n341_), .A2(new_n351_), .A3(new_n378_), .A4(new_n375_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n258_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT33), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n257_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n254_), .B1(new_n246_), .B2(new_n241_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n243_), .A2(new_n244_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n239_), .A2(new_n240_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n245_), .A2(new_n247_), .A3(KEYINPUT33), .A4(new_n254_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n382_), .A2(new_n363_), .A3(new_n386_), .A4(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n380_), .A2(new_n388_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n292_), .A2(new_n296_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n366_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n210_), .B(KEYINPUT31), .Z(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G15gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G71gat), .B(G99gat), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n395_), .B(new_n396_), .Z(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n331_), .A2(KEYINPUT30), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n331_), .A2(KEYINPUT30), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n400_), .A2(G43gat), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G43gat), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n331_), .A2(KEYINPUT30), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(new_n399_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n398_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(G43gat), .B1(new_n400_), .B2(new_n401_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n403_), .A3(new_n399_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n397_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n406_), .A2(KEYINPUT86), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT86), .B1(new_n406_), .B2(new_n409_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n393_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n411_), .A2(new_n393_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n390_), .A2(new_n365_), .A3(new_n414_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n258_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n392_), .A2(new_n415_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G190gat), .B(G218gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(G134gat), .ZN(new_n421_));
  INV_X1    g220(.A(G162gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT36), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NOR3_X1   g227(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT66), .ZN(new_n435_));
  AND2_X1   g234(.A1(G85gat), .A2(G92gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G85gat), .A2(G92gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G85gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n343_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G85gat), .A2(G92gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(KEYINPUT66), .A3(new_n441_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n430_), .A2(new_n434_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT8), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT68), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n438_), .A2(new_n442_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT7), .ZN(new_n447_));
  INV_X1    g246(.A(G99gat), .ZN(new_n448_));
  INV_X1    g247(.A(G106gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G99gat), .A2(G106gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n450_), .A2(new_n453_), .A3(new_n431_), .A4(new_n427_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n446_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT68), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(KEYINPUT8), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n446_), .A2(new_n444_), .A3(new_n454_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT67), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT67), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n446_), .A2(new_n460_), .A3(new_n444_), .A4(new_n454_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n445_), .A2(new_n457_), .A3(new_n459_), .A4(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(KEYINPUT10), .B(G99gat), .Z(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n449_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n440_), .A2(new_n441_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT9), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT64), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT64), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT9), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  OAI22_X1  g269(.A1(new_n465_), .A2(new_n470_), .B1(new_n441_), .B2(new_n467_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n471_), .A2(KEYINPUT65), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(KEYINPUT65), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n464_), .B(new_n434_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n462_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G29gat), .B(G36gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(new_n403_), .ZN(new_n477_));
  INV_X1    g276(.A(G50gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT35), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G232gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT34), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n475_), .A2(new_n479_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT73), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n485_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n462_), .A2(new_n474_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT69), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT69), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n462_), .A2(new_n490_), .A3(new_n474_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n479_), .A2(KEYINPUT15), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n477_), .B(G50gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT15), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT72), .B1(new_n492_), .B2(new_n497_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n462_), .A2(new_n490_), .A3(new_n474_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n490_), .B1(new_n462_), .B2(new_n474_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT72), .B(new_n497_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n486_), .B(new_n487_), .C1(new_n498_), .C2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n483_), .A2(new_n480_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n504_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n506_), .B(new_n484_), .C1(new_n498_), .C2(new_n502_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(KEYINPUT74), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT74), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n497_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT72), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n504_), .B1(new_n512_), .B2(new_n501_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n509_), .B1(new_n513_), .B2(new_n484_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n426_), .B(new_n505_), .C1(new_n508_), .C2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(KEYINPUT74), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n513_), .A2(new_n509_), .A3(new_n484_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n516_), .A2(new_n517_), .B1(new_n504_), .B2(new_n503_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n423_), .B(new_n424_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n515_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT75), .B1(new_n518_), .B2(new_n519_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(KEYINPUT37), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT37), .ZN(new_n523_));
  OAI221_X1 g322(.A(new_n515_), .B1(KEYINPUT75), .B2(new_n523_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G183gat), .B(G211gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G155gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT79), .B(G127gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532_));
  OR3_X1    g331(.A1(new_n531_), .A2(KEYINPUT77), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n532_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(G1gat), .ZN(new_n536_));
  INV_X1    g335(.A(G8gat), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT14), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n538_), .A2(KEYINPUT76), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(KEYINPUT76), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G15gat), .B(G22gat), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G1gat), .B(G8gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n547_));
  XOR2_X1   g346(.A(G71gat), .B(G78gat), .Z(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n547_), .A2(new_n548_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n544_), .B(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n535_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n533_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT80), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n419_), .A2(new_n525_), .A3(new_n559_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n462_), .A2(new_n551_), .A3(new_n474_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n488_), .A2(new_n552_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT12), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n551_), .A2(new_n563_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n564_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n565_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n551_), .B1(new_n462_), .B2(new_n474_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n569_), .B1(new_n561_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G120gat), .B(G148gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G176gat), .B(G204gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n575_), .B(new_n576_), .Z(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n572_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n568_), .A2(new_n571_), .A3(new_n577_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT13), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n579_), .A2(KEYINPUT13), .A3(new_n580_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT71), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n585_), .A2(KEYINPUT71), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n494_), .B(KEYINPUT81), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(new_n544_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(G229gat), .A3(G233gat), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n497_), .A2(new_n544_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n592_), .B(new_n593_), .C1(new_n544_), .C2(new_n589_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G169gat), .B(G197gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G141gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT82), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(G113gat), .Z(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n595_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n591_), .A2(new_n594_), .A3(new_n599_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n587_), .A2(new_n588_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n560_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT103), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT103), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n560_), .A2(new_n608_), .A3(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n258_), .B(KEYINPUT104), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(new_n536_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT38), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n520_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n419_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n605_), .A3(new_n558_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n617_), .B2(new_n418_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n612_), .A2(new_n613_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n614_), .A2(new_n618_), .A3(new_n619_), .ZN(G1324gat));
  AOI22_X1  g419(.A1(new_n302_), .A2(new_n365_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n621_));
  OAI22_X1  g420(.A1(new_n621_), .A2(new_n414_), .B1(new_n258_), .B2(new_n416_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n520_), .A3(new_n558_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n588_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n586_), .ZN(new_n625_));
  NOR4_X1   g424(.A1(new_n623_), .A2(new_n604_), .A3(new_n625_), .A4(new_n365_), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT106), .B1(new_n626_), .B2(new_n537_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT106), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n628_), .B(G8gat), .C1(new_n617_), .C2(new_n365_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n629_), .A3(KEYINPUT39), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n631_));
  OAI211_X1 g430(.A(KEYINPUT106), .B(new_n631_), .C1(new_n626_), .C2(new_n537_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(G8gat), .B1(new_n607_), .B2(new_n609_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT105), .ZN(new_n635_));
  INV_X1    g434(.A(new_n365_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n635_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n633_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n633_), .B(KEYINPUT40), .C1(new_n637_), .C2(new_n638_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1325gat));
  OAI21_X1  g442(.A(G15gat), .B1(new_n617_), .B2(new_n415_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT41), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n606_), .A2(G15gat), .A3(new_n415_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1326gat));
  OAI21_X1  g446(.A(G22gat), .B1(new_n617_), .B2(new_n390_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT42), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n390_), .A2(G22gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n606_), .B2(new_n650_), .ZN(G1327gat));
  NAND4_X1  g450(.A1(new_n605_), .A2(new_n615_), .A3(new_n622_), .A4(new_n559_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n258_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n522_), .A2(new_n524_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n419_), .B2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n525_), .A2(new_n622_), .A3(KEYINPUT43), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n657_), .A2(new_n605_), .A3(new_n559_), .A4(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n661_), .A2(G29gat), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n659_), .A2(new_n660_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n611_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n654_), .B1(new_n662_), .B2(new_n665_), .ZN(G1328gat));
  INV_X1    g465(.A(KEYINPUT46), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n661_), .A2(new_n636_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G36gat), .B1(new_n669_), .B2(new_n663_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT45), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n652_), .A2(G36gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n636_), .ZN(new_n673_));
  NOR4_X1   g472(.A1(new_n652_), .A2(KEYINPUT45), .A3(G36gat), .A4(new_n365_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n668_), .B1(new_n670_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(G36gat), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n659_), .A2(new_n660_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n365_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n681_), .A2(KEYINPUT107), .A3(new_n675_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n667_), .B1(new_n677_), .B2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n670_), .A2(new_n676_), .A3(new_n668_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT107), .B1(new_n681_), .B2(new_n675_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(KEYINPUT46), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(G1329gat));
  OAI21_X1  g486(.A(new_n403_), .B1(new_n652_), .B2(new_n415_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT108), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n679_), .A2(new_n414_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n661_), .A2(G43gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n689_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g492(.A1(new_n297_), .A2(new_n301_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n661_), .A2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G50gat), .B1(new_n695_), .B2(new_n663_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT109), .Z(new_n697_));
  NAND3_X1  g496(.A1(new_n653_), .A2(new_n478_), .A3(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1331gat));
  NOR2_X1   g498(.A1(new_n559_), .A2(new_n603_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n616_), .A2(new_n625_), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(G57gat), .A3(new_n258_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT111), .Z(new_n704_));
  INV_X1    g503(.A(new_n625_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n603_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n560_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G57gat), .B1(new_n708_), .B2(new_n611_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT110), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n704_), .A2(new_n710_), .ZN(G1332gat));
  INV_X1    g510(.A(G64gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n702_), .B2(new_n636_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT112), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n713_), .A2(new_n714_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT48), .ZN(new_n717_));
  OR3_X1    g516(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n708_), .A2(new_n712_), .A3(new_n636_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n718_), .A2(new_n719_), .A3(new_n720_), .ZN(G1333gat));
  OAI21_X1  g520(.A(G71gat), .B1(new_n701_), .B2(new_n415_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT49), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n415_), .A2(G71gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n707_), .B2(new_n724_), .ZN(G1334gat));
  OAI21_X1  g524(.A(G78gat), .B1(new_n701_), .B2(new_n390_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT50), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n390_), .A2(G78gat), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT113), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n707_), .B2(new_n729_), .ZN(G1335gat));
  INV_X1    g529(.A(new_n559_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n419_), .A2(new_n520_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n706_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n439_), .B1(new_n733_), .B2(new_n664_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT114), .Z(new_n735_));
  NAND4_X1  g534(.A1(new_n706_), .A2(new_n657_), .A3(new_n559_), .A4(new_n658_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n258_), .A2(G85gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(G1336gat));
  INV_X1    g538(.A(new_n733_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G92gat), .B1(new_n740_), .B2(new_n636_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n736_), .A2(new_n343_), .A3(new_n365_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n736_), .B2(new_n415_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n740_), .A2(new_n463_), .A3(new_n414_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT51), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n746_), .A2(new_n750_), .A3(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1338gat));
  OAI21_X1  g551(.A(G106gat), .B1(new_n736_), .B2(new_n390_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT52), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n740_), .A2(new_n449_), .A3(new_n694_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT53), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n754_), .A2(new_n758_), .A3(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1339gat));
  AOI21_X1  g559(.A(new_n565_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n568_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n566_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n462_), .A2(new_n551_), .A3(new_n474_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n766_), .B1(new_n570_), .B2(KEYINPUT12), .ZN(new_n767_));
  NOR4_X1   g566(.A1(new_n765_), .A2(new_n767_), .A3(new_n762_), .A4(new_n569_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n577_), .B1(new_n763_), .B2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n770_), .A2(KEYINPUT56), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  AOI211_X1 g571(.A(new_n772_), .B(new_n577_), .C1(new_n763_), .C2(new_n769_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n603_), .B(new_n580_), .C1(new_n771_), .C2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT116), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n765_), .A2(new_n767_), .A3(new_n569_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n569_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(KEYINPUT55), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n578_), .B1(new_n778_), .B2(new_n768_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n772_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n770_), .A2(KEYINPUT56), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n603_), .A4(new_n580_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n599_), .B1(new_n590_), .B2(new_n593_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n592_), .B1(new_n544_), .B2(new_n589_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n593_), .B2(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(new_n602_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n581_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n775_), .A2(new_n784_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n520_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(KEYINPUT57), .A3(new_n520_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n779_), .A2(KEYINPUT117), .A3(new_n772_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n770_), .B2(KEYINPUT56), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n797_), .A3(new_n781_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n788_), .A2(new_n580_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(KEYINPUT58), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT118), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(new_n799_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n798_), .A2(new_n799_), .A3(new_n805_), .A4(KEYINPUT58), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n525_), .A2(new_n801_), .A3(new_n804_), .A4(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n793_), .A2(new_n794_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n558_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n656_), .A2(new_n585_), .A3(new_n700_), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n811_), .A2(KEYINPUT54), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(KEYINPUT54), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n810_), .A2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n416_), .A2(new_n664_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818_), .B2(new_n603_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n808_), .A2(new_n809_), .B1(new_n813_), .B2(new_n812_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n816_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT59), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n814_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824_));
  AND4_X1   g623(.A1(new_n525_), .A2(new_n801_), .A3(new_n804_), .A4(new_n806_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT57), .B1(new_n790_), .B2(new_n520_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n793_), .A2(KEYINPUT119), .A3(new_n807_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n794_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n823_), .B1(new_n829_), .B2(new_n559_), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n821_), .A2(KEYINPUT59), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n603_), .B(new_n822_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n819_), .B1(new_n833_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g633(.A(new_n822_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n835_));
  OAI21_X1  g634(.A(G120gat), .B1(new_n835_), .B2(new_n705_), .ZN(new_n836_));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n705_), .B2(KEYINPUT60), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n818_), .B(new_n838_), .C1(KEYINPUT60), .C2(new_n837_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(G1341gat));
  INV_X1    g639(.A(G127gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n817_), .B2(new_n559_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n842_), .A2(KEYINPUT120), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(KEYINPUT120), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT121), .B(G127gat), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n809_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n822_), .B(new_n846_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n843_), .A2(new_n844_), .A3(new_n848_), .ZN(G1342gat));
  AOI21_X1  g648(.A(G134gat), .B1(new_n818_), .B2(new_n615_), .ZN(new_n850_));
  OAI211_X1 g649(.A(G134gat), .B(new_n822_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n852_), .B2(new_n525_), .ZN(G1343gat));
  NOR2_X1   g652(.A1(new_n390_), .A2(new_n414_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(new_n365_), .A3(new_n611_), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n855_), .B(KEYINPUT122), .Z(new_n856_));
  NAND2_X1  g655(.A1(new_n815_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n604_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT123), .B(G141gat), .Z(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1344gat));
  NOR2_X1   g659(.A1(new_n857_), .A2(new_n705_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(new_n219_), .ZN(G1345gat));
  NOR2_X1   g661(.A1(new_n857_), .A2(new_n559_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT61), .B(G155gat), .Z(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1346gat));
  NOR3_X1   g664(.A1(new_n857_), .A2(new_n422_), .A3(new_n656_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n422_), .B1(new_n857_), .B2(new_n520_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n867_), .A2(KEYINPUT124), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(KEYINPUT124), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n866_), .B1(new_n868_), .B2(new_n869_), .ZN(G1347gat));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n664_), .A2(new_n636_), .A3(new_n414_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT125), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n694_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n830_), .A2(new_n604_), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(G169gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n871_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n829_), .A2(new_n559_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n603_), .B(new_n874_), .C1(new_n879_), .C2(new_n823_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n876_), .A2(new_n323_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n878_), .A2(new_n881_), .A3(new_n882_), .ZN(G1348gat));
  NOR2_X1   g682(.A1(new_n830_), .A2(new_n875_), .ZN(new_n884_));
  AOI21_X1  g683(.A(G176gat), .B1(new_n884_), .B2(new_n625_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n820_), .A2(new_n875_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n705_), .A2(new_n324_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1349gat));
  AOI21_X1  g687(.A(G183gat), .B1(new_n886_), .B2(new_n731_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n558_), .A2(new_n336_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n884_), .B2(new_n890_), .ZN(G1350gat));
  NAND3_X1  g690(.A1(new_n884_), .A2(new_n615_), .A3(new_n309_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n830_), .A2(new_n656_), .A3(new_n875_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n319_), .B2(new_n893_), .ZN(G1351gat));
  INV_X1    g693(.A(new_n854_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n365_), .A2(new_n258_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n820_), .A2(new_n895_), .A3(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n603_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n625_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n902_));
  XOR2_X1   g701(.A(new_n901_), .B(new_n902_), .Z(G1353gat));
  NOR2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906_));
  NOR4_X1   g705(.A1(new_n820_), .A2(new_n809_), .A3(new_n895_), .A4(new_n897_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n815_), .A2(new_n558_), .A3(new_n854_), .A4(new_n896_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n908_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n910_), .A2(KEYINPUT127), .A3(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n905_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n907_), .A2(new_n906_), .A3(new_n908_), .ZN(new_n914_));
  OAI21_X1  g713(.A(KEYINPUT127), .B1(new_n910_), .B2(new_n911_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n914_), .A2(new_n915_), .A3(new_n904_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n913_), .A2(new_n916_), .ZN(G1354gat));
  AND3_X1   g716(.A1(new_n898_), .A2(G218gat), .A3(new_n525_), .ZN(new_n918_));
  AOI21_X1  g717(.A(G218gat), .B1(new_n898_), .B2(new_n615_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1355gat));
endmodule


