//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_;
  XOR2_X1   g000(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n202_));
  XNOR2_X1  g001(.A(G120gat), .B(G148gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G176gat), .B(G204gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G230gat), .A2(G233gat), .ZN(new_n208_));
  INV_X1    g007(.A(G71gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT65), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G71gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n212_), .A3(G78gat), .ZN(new_n213_));
  INV_X1    g012(.A(G57gat), .ZN(new_n214_));
  INV_X1    g013(.A(G64gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G57gat), .A2(G64gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n213_), .A2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(G78gat), .B1(new_n210_), .B2(new_n212_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT66), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n210_), .A2(new_n212_), .ZN(new_n223_));
  INV_X1    g022(.A(G78gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n219_), .A4(new_n213_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(new_n227_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n216_), .A2(new_n218_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(new_n217_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n222_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G85gat), .B(G92gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT9), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT10), .B(G99gat), .Z(new_n237_));
  INV_X1    g036(.A(G106gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G85gat), .ZN(new_n240_));
  INV_X1    g039(.A(G92gat), .ZN(new_n241_));
  OR3_X1    g040(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT9), .ZN(new_n242_));
  NAND3_X1  g041(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n236_), .A2(new_n239_), .A3(new_n242_), .A4(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT7), .ZN(new_n248_));
  INV_X1    g047(.A(G99gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(new_n238_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G99gat), .A2(G106gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT6), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n250_), .A2(new_n253_), .A3(new_n243_), .A4(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n235_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT8), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(KEYINPUT64), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(KEYINPUT64), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(new_n255_), .B2(new_n235_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n259_), .B1(new_n262_), .B2(new_n258_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n232_), .A2(new_n233_), .B1(new_n247_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n232_), .A2(new_n233_), .A3(new_n247_), .A4(new_n263_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n208_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n258_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n254_), .ZN(new_n270_));
  NOR3_X1   g069(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n234_), .B1(new_n272_), .B2(new_n246_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n269_), .B1(new_n273_), .B2(new_n261_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT67), .B1(new_n274_), .B2(new_n259_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n258_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n269_), .B1(new_n255_), .B2(new_n235_), .ZN(new_n278_));
  NOR3_X1   g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n247_), .B1(new_n275_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT12), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n222_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n230_), .B1(new_n222_), .B2(new_n227_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n247_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n274_), .B2(new_n259_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n281_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n283_), .B(new_n208_), .C1(new_n264_), .C2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n207_), .B1(new_n268_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n268_), .A2(new_n290_), .A3(new_n207_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(KEYINPUT69), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n295_));
  INV_X1    g094(.A(new_n293_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n295_), .B1(new_n296_), .B2(new_n291_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n294_), .A2(new_n297_), .A3(KEYINPUT13), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT13), .B1(new_n294_), .B2(new_n297_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT70), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT70), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT23), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n308_), .B1(G183gat), .B2(G190gat), .ZN(new_n309_));
  AND2_X1   g108(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n310_));
  OAI21_X1  g109(.A(G169gat), .B1(new_n310_), .B2(G176gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n309_), .B(new_n311_), .C1(new_n313_), .C2(new_n310_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n308_), .B1(KEYINPUT24), .B2(new_n313_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT81), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G169gat), .ZN(new_n318_));
  INV_X1    g117(.A(G176gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321_));
  NOR3_X1   g120(.A1(new_n320_), .A2(new_n321_), .A3(new_n312_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT25), .B(G183gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT26), .B(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n322_), .B1(KEYINPUT80), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(KEYINPUT80), .B2(new_n325_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n314_), .B1(new_n317_), .B2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT30), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT83), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G71gat), .B(G99gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G227gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G15gat), .B(G43gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n331_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n329_), .B(new_n330_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G127gat), .B(G134gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G113gat), .B(G120gat), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n340_), .B(new_n341_), .Z(new_n342_));
  XOR2_X1   g141(.A(new_n342_), .B(KEYINPUT31), .Z(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n339_), .A2(new_n343_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G155gat), .B(G162gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT86), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349_));
  OR4_X1    g148(.A1(new_n349_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n350_));
  INV_X1    g149(.A(G141gat), .ZN(new_n351_));
  INV_X1    g150(.A(G148gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n353_), .B1(new_n349_), .B2(KEYINPUT3), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT2), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n350_), .A2(new_n354_), .A3(new_n357_), .A4(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n348_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G155gat), .ZN(new_n361_));
  INV_X1    g160(.A(G162gat), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT1), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(G155gat), .B2(G162gat), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n361_), .A2(new_n362_), .A3(KEYINPUT1), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n353_), .B(new_n355_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n360_), .A2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G197gat), .B(G204gat), .Z(new_n368_));
  OR2_X1    g167(.A1(new_n368_), .A2(KEYINPUT21), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(KEYINPUT21), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G211gat), .B(G218gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n370_), .A2(new_n371_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n367_), .A2(KEYINPUT29), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G22gat), .B(G50gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT28), .ZN(new_n376_));
  INV_X1    g175(.A(G233gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT87), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n378_), .A2(G228gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(G228gat), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n377_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n376_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n374_), .B(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n367_), .A2(KEYINPUT29), .ZN(new_n384_));
  XOR2_X1   g183(.A(G78gat), .B(G106gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n383_), .B(new_n386_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n345_), .A2(new_n346_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT4), .B1(new_n367_), .B2(new_n342_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT93), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n367_), .A2(new_n392_), .A3(new_n342_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n390_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(new_n367_), .B(new_n342_), .Z(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n389_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(new_n240_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT0), .B(G57gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n404_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n397_), .A2(new_n399_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n315_), .A2(new_n322_), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n324_), .B(KEYINPUT88), .Z(new_n412_));
  INV_X1    g211(.A(new_n323_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n411_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n309_), .B(KEYINPUT90), .ZN(new_n415_));
  INV_X1    g214(.A(new_n320_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n416_), .A2(KEYINPUT89), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(KEYINPUT89), .ZN(new_n418_));
  XOR2_X1   g217(.A(KEYINPUT22), .B(G169gat), .Z(new_n419_));
  OAI211_X1 g218(.A(new_n417_), .B(new_n418_), .C1(G176gat), .C2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n414_), .B1(new_n415_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n372_), .A2(new_n373_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G226gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT19), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n328_), .B2(new_n422_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n423_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT91), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n427_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(new_n422_), .B2(new_n328_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n425_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT91), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n423_), .A2(new_n428_), .A3(new_n434_), .A4(new_n426_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n430_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G64gat), .B(G92gat), .Z(new_n437_));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n430_), .A2(new_n433_), .A3(new_n443_), .A4(new_n435_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n410_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n432_), .A2(new_n425_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n426_), .B1(new_n423_), .B2(new_n428_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n441_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n448_), .A2(new_n444_), .A3(KEYINPUT27), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n388_), .A2(new_n409_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n409_), .A2(new_n387_), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n445_), .A2(new_n452_), .A3(new_n449_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n442_), .A2(new_n444_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n398_), .A2(new_n390_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n404_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n389_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT94), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n457_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n458_), .A2(new_n459_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n407_), .A2(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n407_), .A2(new_n463_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n462_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n455_), .A2(new_n466_), .A3(KEYINPUT95), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n443_), .A2(KEYINPUT32), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT96), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n469_), .A2(new_n430_), .A3(new_n435_), .A4(new_n433_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n468_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n408_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT95), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n462_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n473_), .B1(new_n474_), .B2(new_n454_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n467_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n387_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n453_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n346_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(KEYINPUT84), .A3(new_n344_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n451_), .B1(new_n478_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G29gat), .B(G36gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G43gat), .B(G50gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n288_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G232gat), .A2(G233gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT34), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(KEYINPUT35), .B2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n277_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n259_), .B(KEYINPUT67), .C1(new_n258_), .C2(new_n262_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n287_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n487_), .B(KEYINPUT15), .Z(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n490_), .A2(KEYINPUT35), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n497_), .B(KEYINPUT71), .Z(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  OR3_X1    g298(.A1(new_n491_), .A2(new_n496_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G190gat), .B(G218gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G134gat), .B(G162gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n502_), .B(new_n503_), .Z(new_n504_));
  OAI21_X1  g303(.A(new_n499_), .B1(new_n491_), .B2(new_n496_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n500_), .A2(new_n501_), .A3(new_n504_), .A4(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT72), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT37), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n500_), .A2(new_n505_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n504_), .B(KEYINPUT36), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n509_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n508_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT73), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n500_), .A2(new_n514_), .A3(new_n505_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n514_), .B1(new_n500_), .B2(new_n505_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n511_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT74), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT74), .B(new_n511_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n507_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n513_), .B1(new_n521_), .B2(KEYINPUT37), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G183gat), .B(G211gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(G127gat), .B(G155gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(G1gat), .ZN(new_n531_));
  INV_X1    g330(.A(G8gat), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT14), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT75), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G15gat), .B(G22gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G1gat), .B(G8gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT76), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n536_), .B(new_n538_), .Z(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G231gat), .A2(G233gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n286_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n286_), .A2(new_n541_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n540_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(new_n542_), .A3(new_n539_), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT17), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n530_), .B1(new_n548_), .B2(new_n528_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n547_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(KEYINPUT78), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(KEYINPUT78), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n552_), .B(new_n530_), .C1(new_n528_), .C2(new_n548_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n523_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n539_), .B(new_n487_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n539_), .A2(new_n495_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n539_), .A2(new_n487_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G169gat), .B(G197gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT79), .B1(new_n564_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT79), .ZN(new_n569_));
  INV_X1    g368(.A(new_n567_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n560_), .A2(new_n569_), .A3(new_n563_), .A4(new_n570_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n568_), .A2(new_n571_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n306_), .A2(new_n484_), .A3(new_n556_), .A4(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(KEYINPUT98), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(KEYINPUT98), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n408_), .B(KEYINPUT99), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(G1gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT100), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT100), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n578_), .A2(new_n583_), .A3(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT38), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n472_), .ZN(new_n588_));
  AOI22_X1  g387(.A1(new_n460_), .A2(new_n461_), .B1(new_n463_), .B2(new_n407_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n589_), .A2(new_n444_), .A3(new_n442_), .A4(new_n465_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n588_), .B1(new_n590_), .B2(new_n473_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n387_), .B1(new_n591_), .B2(new_n467_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n482_), .B(new_n480_), .C1(new_n592_), .C2(new_n453_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n521_), .B1(new_n593_), .B2(new_n451_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n300_), .A2(new_n573_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n554_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G1gat), .B1(new_n598_), .B2(new_n409_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n582_), .A2(KEYINPUT38), .A3(new_n584_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n587_), .A2(new_n599_), .A3(new_n600_), .ZN(G1324gat));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n598_), .B2(new_n450_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n450_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n594_), .A2(KEYINPUT101), .A3(new_n604_), .A4(new_n597_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(G8gat), .A3(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(KEYINPUT102), .A3(KEYINPUT39), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(KEYINPUT39), .B2(new_n606_), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT102), .B1(new_n606_), .B2(KEYINPUT39), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n604_), .A2(new_n532_), .ZN(new_n610_));
  OAI22_X1  g409(.A1(new_n608_), .A2(new_n609_), .B1(new_n577_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT40), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI221_X1 g412(.A(KEYINPUT40), .B1(new_n577_), .B2(new_n610_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1325gat));
  INV_X1    g414(.A(G15gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n483_), .A2(new_n616_), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n577_), .A2(KEYINPUT103), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n598_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n616_), .B1(new_n619_), .B2(new_n483_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT41), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT103), .B1(new_n577_), .B2(new_n617_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n618_), .A2(new_n621_), .A3(new_n622_), .ZN(G1326gat));
  OAI21_X1  g422(.A(G22gat), .B1(new_n598_), .B2(new_n477_), .ZN(new_n624_));
  XOR2_X1   g423(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n625_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n477_), .A2(G22gat), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n626_), .B(new_n627_), .C1(new_n577_), .C2(new_n628_), .ZN(G1327gat));
  NAND2_X1  g428(.A1(new_n521_), .A2(new_n596_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT108), .ZN(new_n631_));
  AND4_X1   g430(.A1(new_n484_), .A2(new_n573_), .A3(new_n300_), .A4(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(G29gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n633_), .A3(new_n408_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n595_), .A2(new_n554_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT43), .B1(new_n523_), .B2(KEYINPUT105), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n484_), .A2(new_n636_), .A3(new_n522_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n636_), .B1(new_n484_), .B2(new_n522_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n579_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n484_), .A2(new_n522_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n636_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n637_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(KEYINPUT44), .A3(new_n635_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n642_), .A2(new_n643_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n633_), .B1(new_n649_), .B2(KEYINPUT106), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT44), .B1(new_n647_), .B2(new_n635_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n635_), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n641_), .B(new_n652_), .C1(new_n646_), .C2(new_n637_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n643_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n650_), .A2(KEYINPUT107), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT107), .B1(new_n650_), .B2(new_n656_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n634_), .B1(new_n657_), .B2(new_n658_), .ZN(G1328gat));
  INV_X1    g458(.A(KEYINPUT46), .ZN(new_n660_));
  INV_X1    g459(.A(G36gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n632_), .A2(new_n661_), .A3(new_n604_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT45), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n642_), .A2(new_n604_), .A3(new_n648_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n665_), .B2(G36gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n660_), .B1(new_n666_), .B2(KEYINPUT109), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT109), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n661_), .B1(new_n654_), .B2(new_n604_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n668_), .B(KEYINPUT46), .C1(new_n669_), .C2(new_n664_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n667_), .A2(new_n670_), .ZN(G1329gat));
  INV_X1    g470(.A(G43gat), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n632_), .A2(new_n672_), .A3(new_n483_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n345_), .A2(new_n346_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n654_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n675_), .B2(G43gat), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g476(.A(G50gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n632_), .A2(new_n678_), .A3(new_n387_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n651_), .A2(new_n653_), .A3(new_n477_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n680_), .B2(new_n678_), .ZN(G1331gat));
  NAND2_X1  g480(.A1(new_n484_), .A2(new_n572_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT110), .Z(new_n683_));
  AND3_X1   g482(.A1(new_n683_), .A2(new_n556_), .A3(new_n301_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G57gat), .B1(new_n684_), .B2(new_n643_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n594_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n554_), .A2(new_n572_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n305_), .A2(new_n687_), .ZN(new_n688_));
  OR3_X1    g487(.A1(new_n686_), .A2(new_n688_), .A3(KEYINPUT111), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT111), .B1(new_n686_), .B2(new_n688_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n409_), .A2(new_n214_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n685_), .B1(new_n691_), .B2(new_n692_), .ZN(G1332gat));
  NAND3_X1  g492(.A1(new_n684_), .A2(new_n215_), .A3(new_n604_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT48), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n691_), .A2(new_n604_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(G64gat), .ZN(new_n697_));
  AOI211_X1 g496(.A(KEYINPUT48), .B(new_n215_), .C1(new_n691_), .C2(new_n604_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1333gat));
  NAND3_X1  g498(.A1(new_n684_), .A2(new_n209_), .A3(new_n483_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT49), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n691_), .A2(new_n483_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(G71gat), .ZN(new_n703_));
  AOI211_X1 g502(.A(KEYINPUT49), .B(new_n209_), .C1(new_n691_), .C2(new_n483_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(G1334gat));
  NAND3_X1  g504(.A1(new_n684_), .A2(new_n224_), .A3(new_n387_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n689_), .A2(new_n387_), .A3(new_n690_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT50), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(G78gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n707_), .B2(G78gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n706_), .B(KEYINPUT112), .C1(new_n710_), .C2(new_n709_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1335gat));
  AND3_X1   g514(.A1(new_n683_), .A2(new_n305_), .A3(new_n631_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G85gat), .B1(new_n716_), .B2(new_n643_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n301_), .A2(new_n596_), .A3(new_n572_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n646_), .B2(new_n637_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n409_), .A2(new_n240_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n717_), .B1(new_n719_), .B2(new_n720_), .ZN(G1336gat));
  INV_X1    g520(.A(KEYINPUT113), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n716_), .A2(new_n604_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n241_), .ZN(new_n724_));
  AOI211_X1 g523(.A(KEYINPUT113), .B(G92gat), .C1(new_n716_), .C2(new_n604_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n719_), .A2(G92gat), .A3(new_n604_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(G1337gat));
  NAND3_X1  g526(.A1(new_n716_), .A2(new_n674_), .A3(new_n237_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n719_), .A2(new_n483_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n249_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT51), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n728_), .B(new_n732_), .C1(new_n249_), .C2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1338gat));
  NAND3_X1  g533(.A1(new_n716_), .A2(new_n238_), .A3(new_n387_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n719_), .A2(new_n387_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G106gat), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT52), .B(new_n238_), .C1(new_n719_), .C2(new_n387_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT53), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT53), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n735_), .B(new_n742_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1339gat));
  INV_X1    g543(.A(new_n521_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT117), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n572_), .A2(new_n296_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n283_), .B1(new_n289_), .B2(new_n264_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n208_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n266_), .A2(KEYINPUT12), .ZN(new_n753_));
  AOI22_X1  g552(.A1(new_n753_), .A2(new_n265_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n754_), .B2(new_n208_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n264_), .B1(KEYINPUT12), .B2(new_n266_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT12), .B1(new_n284_), .B2(new_n285_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n494_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n752_), .ZN(new_n759_));
  NOR4_X1   g558(.A1(new_n756_), .A2(new_n758_), .A3(new_n750_), .A4(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n751_), .B1(new_n755_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT116), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n763_), .B(new_n751_), .C1(new_n755_), .C2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n206_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n767_), .B(new_n207_), .C1(new_n762_), .C2(new_n764_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n746_), .B(new_n747_), .C1(new_n766_), .C2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n561_), .A2(new_n559_), .A3(new_n562_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n570_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n568_), .A2(new_n571_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n294_), .A3(new_n297_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n769_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n764_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n290_), .A2(new_n759_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n754_), .A2(new_n208_), .A3(new_n752_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n763_), .B1(new_n778_), .B2(new_n751_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n206_), .B1(new_n775_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n767_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n207_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT56), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n746_), .B1(new_n784_), .B2(new_n747_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n745_), .B1(new_n774_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT57), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n782_), .B2(KEYINPUT56), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n780_), .A2(KEYINPUT118), .A3(new_n767_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n783_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n772_), .A2(new_n293_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n792_), .A2(KEYINPUT58), .A3(new_n793_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n522_), .A3(new_n797_), .ZN(new_n798_));
  OAI211_X1 g597(.A(KEYINPUT57), .B(new_n745_), .C1(new_n774_), .C2(new_n785_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n788_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n596_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n300_), .A2(new_n687_), .A3(KEYINPUT114), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n554_), .B(new_n572_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n802_), .B1(new_n807_), .B2(new_n523_), .ZN(new_n808_));
  AOI211_X1 g607(.A(KEYINPUT54), .B(new_n522_), .C1(new_n803_), .C2(new_n806_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n801_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n388_), .A2(new_n450_), .A3(new_n643_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(new_n813_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n810_), .B1(new_n800_), .B2(new_n596_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT59), .B1(new_n817_), .B2(new_n814_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n816_), .A2(new_n573_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G113gat), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n812_), .A2(new_n815_), .ZN(new_n821_));
  OR3_X1    g620(.A1(new_n821_), .A2(G113gat), .A3(new_n572_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT119), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n820_), .A2(new_n825_), .A3(new_n822_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1340gat));
  NAND3_X1  g626(.A1(new_n816_), .A2(new_n305_), .A3(new_n818_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(G120gat), .B1(new_n828_), .B2(new_n829_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT60), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(G120gat), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n300_), .A2(KEYINPUT60), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(G120gat), .ZN(new_n835_));
  OAI22_X1  g634(.A1(new_n830_), .A2(new_n831_), .B1(new_n821_), .B2(new_n835_), .ZN(G1341gat));
  NAND4_X1  g635(.A1(new_n816_), .A2(new_n818_), .A3(G127gat), .A4(new_n554_), .ZN(new_n837_));
  INV_X1    g636(.A(G127gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n821_), .B2(new_n596_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(G1342gat));
  XNOR2_X1  g641(.A(KEYINPUT122), .B(G134gat), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n816_), .A2(new_n818_), .A3(new_n522_), .A4(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(G134gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n821_), .B2(new_n745_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1343gat));
  NOR4_X1   g646(.A1(new_n483_), .A2(new_n604_), .A3(new_n477_), .A4(new_n579_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n812_), .A2(new_n848_), .ZN(new_n849_));
  OR3_X1    g648(.A1(new_n849_), .A2(KEYINPUT124), .A3(new_n572_), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT124), .B1(new_n849_), .B2(new_n572_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT123), .B(G141gat), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1344gat));
  NOR2_X1   g654(.A1(new_n849_), .A2(new_n306_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(new_n352_), .ZN(G1345gat));
  NOR2_X1   g656(.A1(new_n849_), .A2(new_n596_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT61), .B(G155gat), .Z(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1346gat));
  NOR3_X1   g659(.A1(new_n849_), .A2(new_n362_), .A3(new_n523_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n849_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n521_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n362_), .B2(new_n863_), .ZN(G1347gat));
  NOR2_X1   g663(.A1(new_n817_), .A2(new_n450_), .ZN(new_n865_));
  AOI211_X1 g664(.A(new_n387_), .B(new_n643_), .C1(new_n480_), .C2(new_n482_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n573_), .A3(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n867_), .A2(new_n868_), .A3(G169gat), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n867_), .B2(G169gat), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n865_), .A2(new_n866_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n572_), .A2(new_n419_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT125), .ZN(new_n873_));
  OAI22_X1  g672(.A1(new_n869_), .A2(new_n870_), .B1(new_n871_), .B2(new_n873_), .ZN(G1348gat));
  NOR3_X1   g673(.A1(new_n871_), .A2(new_n319_), .A3(new_n306_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n871_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n301_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n319_), .B2(new_n877_), .ZN(G1349gat));
  NOR2_X1   g677(.A1(new_n871_), .A2(new_n596_), .ZN(new_n879_));
  MUX2_X1   g678(.A(G183gat), .B(new_n323_), .S(new_n879_), .Z(G1350gat));
  OAI21_X1  g679(.A(G190gat), .B1(new_n871_), .B2(new_n523_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n745_), .A2(new_n412_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n871_), .B2(new_n882_), .ZN(G1351gat));
  NOR2_X1   g682(.A1(new_n483_), .A2(new_n452_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n865_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n573_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n305_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g688(.A(new_n596_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n812_), .A2(new_n604_), .A3(new_n884_), .A4(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT126), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n865_), .A2(new_n893_), .A3(new_n884_), .A4(new_n890_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1354gat));
  AOI21_X1  g696(.A(G218gat), .B1(new_n885_), .B2(new_n521_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n522_), .A2(G218gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n885_), .B2(new_n899_), .ZN(G1355gat));
endmodule


