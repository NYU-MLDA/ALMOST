//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT1), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT82), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(new_n213_), .A3(new_n206_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT81), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n209_), .A2(new_n214_), .A3(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G141gat), .B(G148gat), .Z(new_n221_));
  AND3_X1   g020(.A1(new_n220_), .A2(KEYINPUT83), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT83), .B1(new_n220_), .B2(new_n221_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n219_), .B1(new_n208_), .B2(new_n207_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G141gat), .A2(G148gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT2), .ZN(new_n227_));
  OR4_X1    g026(.A1(KEYINPUT84), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n228_));
  OAI22_X1  g027(.A1(KEYINPUT84), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT85), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT85), .A4(new_n229_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n225_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT86), .B1(new_n224_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n220_), .A2(new_n221_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT83), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n220_), .A2(KEYINPUT83), .A3(new_n221_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(new_n233_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n225_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT86), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n205_), .B1(new_n235_), .B2(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n246_), .A2(KEYINPUT4), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n240_), .A2(new_n243_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n205_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT4), .B1(new_n246_), .B2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n202_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n246_), .A2(new_n250_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n202_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT94), .B(KEYINPUT0), .Z(new_n257_));
  XNOR2_X1  g056(.A(G1gat), .B(G29gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G57gat), .B(G85gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n252_), .A2(new_n255_), .A3(new_n261_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G197gat), .B(G204gat), .Z(new_n266_));
  NOR2_X1   g065(.A1(G211gat), .A2(G218gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT21), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G211gat), .A2(G218gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(G211gat), .A2(G218gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT88), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n272_), .A2(new_n267_), .A3(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n266_), .B(new_n271_), .C1(new_n274_), .C2(new_n269_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n268_), .A2(KEYINPUT88), .A3(new_n270_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G197gat), .B(G204gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(KEYINPUT21), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n248_), .B2(KEYINPUT29), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G228gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT87), .ZN(new_n283_));
  OR3_X1    g082(.A1(new_n281_), .A2(KEYINPUT89), .A3(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT89), .B1(new_n281_), .B2(new_n283_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n235_), .A2(new_n245_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT29), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n279_), .B(new_n283_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G78gat), .B(G106gat), .Z(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n235_), .A2(new_n245_), .A3(new_n288_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n293_), .A2(KEYINPUT28), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(KEYINPUT28), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G22gat), .B(G50gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n296_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n290_), .B(new_n292_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n291_), .B1(new_n286_), .B2(new_n289_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT90), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n293_), .B(KEYINPUT28), .ZN(new_n303_));
  INV_X1    g102(.A(new_n296_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n302_), .B1(new_n305_), .B2(new_n297_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n300_), .B1(new_n301_), .B2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n290_), .A2(new_n292_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT80), .ZN(new_n311_));
  AND3_X1   g110(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT78), .B1(G183gat), .B2(G190gat), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n311_), .B(KEYINPUT23), .C1(new_n312_), .C2(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n316_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT80), .B1(new_n317_), .B2(KEYINPUT23), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n314_), .B(new_n315_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT79), .B(G176gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT22), .B(G169gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n330_));
  OR2_X1    g129(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n329_), .A2(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT24), .ZN(new_n334_));
  INV_X1    g133(.A(G169gat), .ZN(new_n335_));
  INV_X1    g134(.A(G176gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n337_), .B1(new_n325_), .B2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n333_), .A2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n316_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n317_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT23), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n323_), .A2(new_n328_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT30), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(new_n205_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G227gat), .A2(G233gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT31), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n347_), .B(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G15gat), .B(G43gat), .Z(new_n351_));
  XOR2_X1   g150(.A(G71gat), .B(G99gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n350_), .B(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n308_), .A2(new_n306_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n310_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT20), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n323_), .A2(new_n328_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n340_), .A2(new_n344_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n357_), .B1(new_n360_), .B2(new_n279_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G226gat), .A2(G233gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT19), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT23), .B1(new_n312_), .B2(new_n313_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n311_), .B1(new_n342_), .B2(new_n316_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n329_), .A2(new_n330_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n331_), .A2(new_n332_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NOR3_X1   g169(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n338_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(new_n324_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n367_), .A2(new_n314_), .A3(new_n370_), .A4(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n341_), .A2(new_n315_), .A3(new_n343_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n328_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n361_), .B(new_n364_), .C1(new_n279_), .C2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n279_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT91), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n357_), .B1(new_n345_), .B2(new_n280_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n377_), .A2(new_n382_), .A3(new_n279_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT92), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n384_), .A2(new_n385_), .A3(new_n363_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n385_), .B1(new_n384_), .B2(new_n363_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n378_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G64gat), .B(G92gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n388_), .B(new_n393_), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n394_), .A2(KEYINPUT27), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n378_), .B(new_n393_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT100), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT20), .B1(new_n360_), .B2(new_n279_), .ZN(new_n398_));
  AOI221_X4 g197(.A(KEYINPUT91), .B1(new_n275_), .B2(new_n278_), .C1(new_n374_), .C2(new_n376_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n382_), .B1(new_n377_), .B2(new_n279_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT92), .B1(new_n401_), .B2(new_n364_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n384_), .A2(new_n385_), .A3(new_n363_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT100), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n404_), .A2(new_n405_), .A3(new_n378_), .A4(new_n393_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n377_), .A2(KEYINPUT98), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n377_), .A2(KEYINPUT98), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n280_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n361_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n363_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n363_), .B2(new_n384_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n393_), .B(KEYINPUT99), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n397_), .A2(new_n406_), .A3(KEYINPUT27), .A4(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n415_), .A2(KEYINPUT101), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(KEYINPUT101), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n395_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT102), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n415_), .B(KEYINPUT101), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT102), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(new_n395_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n356_), .B1(new_n419_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n354_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT90), .B1(new_n298_), .B2(new_n299_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n301_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n308_), .B1(new_n427_), .B2(new_n300_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n355_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n424_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n430_), .A2(new_n418_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n265_), .B1(new_n423_), .B2(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT96), .B(KEYINPUT33), .Z(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT95), .B1(new_n256_), .B2(new_n262_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT95), .ZN(new_n435_));
  NOR4_X1   g234(.A1(new_n252_), .A2(new_n255_), .A3(new_n435_), .A4(new_n261_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n433_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT97), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n254_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n261_), .B1(new_n253_), .B2(new_n202_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n394_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(KEYINPUT33), .B2(new_n264_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT97), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n443_), .B(new_n433_), .C1(new_n434_), .C2(new_n436_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n438_), .A2(new_n442_), .A3(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n393_), .A2(KEYINPUT32), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n412_), .A2(new_n446_), .ZN(new_n447_));
  OAI221_X1 g246(.A(new_n447_), .B1(new_n388_), .B2(new_n446_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n428_), .A2(new_n429_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n424_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n432_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT76), .B(G15gat), .ZN(new_n453_));
  INV_X1    g252(.A(G22gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G1gat), .ZN(new_n456_));
  INV_X1    g255(.A(G8gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT14), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G8gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G231gat), .A2(G233gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n461_), .B(new_n462_), .Z(new_n463_));
  XNOR2_X1  g262(.A(G57gat), .B(G64gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT71), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n465_), .A2(KEYINPUT11), .ZN(new_n466_));
  XOR2_X1   g265(.A(G71gat), .B(G78gat), .Z(new_n467_));
  OR2_X1    g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n465_), .A2(KEYINPUT11), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n467_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n463_), .B(new_n471_), .Z(new_n472_));
  XOR2_X1   g271(.A(G183gat), .B(G211gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(G127gat), .B(G155gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n477_), .A2(KEYINPUT17), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n477_), .A2(KEYINPUT17), .ZN(new_n479_));
  OR3_X1    g278(.A1(new_n472_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n471_), .A2(KEYINPUT72), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n471_), .A2(KEYINPUT72), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(new_n463_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n479_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n480_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(G99gat), .ZN(new_n488_));
  INV_X1    g287(.A(G106gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(KEYINPUT69), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n490_), .A2(KEYINPUT7), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G99gat), .A2(G106gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT6), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(KEYINPUT7), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G85gat), .B(G92gat), .Z(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT70), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(KEYINPUT70), .A3(new_n496_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(KEYINPUT8), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT8), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G92gat), .ZN(new_n504_));
  OR3_X1    g303(.A1(new_n504_), .A2(KEYINPUT67), .A3(KEYINPUT9), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(KEYINPUT67), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n507_), .A2(G85gat), .B1(KEYINPUT9), .B2(new_n496_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT68), .ZN(new_n509_));
  XOR2_X1   g308(.A(KEYINPUT10), .B(G99gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT65), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT66), .B(G106gat), .Z(new_n512_));
  OAI21_X1  g311(.A(new_n493_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n501_), .B(new_n503_), .C1(new_n509_), .C2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G29gat), .B(G36gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G43gat), .B(G50gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT15), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G232gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT34), .ZN(new_n521_));
  INV_X1    g320(.A(new_n517_), .ZN(new_n522_));
  OAI221_X1 g321(.A(new_n519_), .B1(KEYINPUT35), .B2(new_n521_), .C1(new_n522_), .C2(new_n514_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n521_), .A2(KEYINPUT35), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  XNOR2_X1  g324(.A(G190gat), .B(G218gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G134gat), .B(G162gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n526_), .B(new_n527_), .Z(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT36), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n531_), .A2(KEYINPUT74), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n529_), .A2(KEYINPUT36), .ZN(new_n533_));
  OR3_X1    g332(.A1(new_n525_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(KEYINPUT74), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n532_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT37), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n531_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(KEYINPUT75), .B(KEYINPUT37), .Z(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n537_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n452_), .A2(new_n487_), .A3(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n481_), .A2(KEYINPUT12), .A3(new_n514_), .A4(new_n482_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n514_), .A2(new_n471_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n514_), .A2(new_n471_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT12), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(new_n545_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n550_), .B(KEYINPUT64), .Z(new_n551_));
  NOR2_X1   g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n545_), .A2(new_n546_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n551_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G176gat), .B(G204gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n556_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n553_), .A2(new_n555_), .A3(new_n561_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT13), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT13), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n563_), .A2(new_n567_), .A3(new_n564_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n461_), .A2(new_n522_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n461_), .B2(new_n518_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G229gat), .A2(G233gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n461_), .B(new_n522_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(G229gat), .A3(G233gat), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G113gat), .B(G141gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G169gat), .B(G197gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(new_n579_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n569_), .A2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n543_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n265_), .B(KEYINPUT103), .Z(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n456_), .A3(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT38), .ZN(new_n589_));
  AOI211_X1 g388(.A(new_n539_), .B(new_n486_), .C1(new_n432_), .C2(new_n451_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n584_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G1gat), .B1(new_n592_), .B2(new_n265_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n593_), .ZN(G1324gat));
  NOR2_X1   g393(.A1(new_n418_), .A2(KEYINPUT102), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n421_), .B1(new_n420_), .B2(new_n395_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n585_), .A2(new_n457_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n599_));
  INV_X1    g398(.A(new_n592_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n597_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n601_), .B2(G8gat), .ZN(new_n602_));
  AOI211_X1 g401(.A(KEYINPUT39), .B(new_n457_), .C1(new_n600_), .C2(new_n597_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n598_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g404(.A(G15gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n585_), .A2(new_n606_), .A3(new_n354_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n600_), .B2(new_n354_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n607_), .B1(new_n610_), .B2(new_n611_), .ZN(G1326gat));
  XNOR2_X1  g411(.A(new_n450_), .B(KEYINPUT105), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n585_), .A2(new_n454_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT42), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n600_), .A2(new_n614_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n616_), .B1(new_n617_), .B2(G22gat), .ZN(new_n618_));
  AOI211_X1 g417(.A(KEYINPUT42), .B(new_n454_), .C1(new_n600_), .C2(new_n614_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n615_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT106), .Z(G1327gat));
  NAND3_X1  g420(.A1(new_n569_), .A2(new_n583_), .A3(new_n486_), .ZN(new_n622_));
  AOI211_X1 g421(.A(new_n538_), .B(new_n622_), .C1(new_n432_), .C2(new_n451_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  OR3_X1    g423(.A1(new_n624_), .A2(G29gat), .A3(new_n265_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n622_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n542_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT107), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT43), .B1(new_n542_), .B2(new_n628_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n452_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n452_), .B2(new_n627_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n626_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT44), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n452_), .A2(new_n627_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n629_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n452_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(KEYINPUT44), .A3(new_n626_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n634_), .A2(new_n640_), .A3(new_n587_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT108), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n641_), .A2(new_n642_), .A3(G29gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n641_), .B2(G29gat), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n625_), .B1(new_n643_), .B2(new_n644_), .ZN(G1328gat));
  INV_X1    g444(.A(KEYINPUT112), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n538_), .B1(new_n432_), .B2(new_n451_), .ZN(new_n647_));
  INV_X1    g446(.A(G36gat), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n647_), .A2(new_n648_), .A3(new_n597_), .A4(new_n626_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT110), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n623_), .A2(KEYINPUT110), .A3(new_n648_), .A4(new_n597_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n651_), .A2(new_n652_), .A3(new_n654_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n634_), .A2(new_n640_), .A3(new_n597_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(G36gat), .B2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(KEYINPUT111), .B(KEYINPUT46), .Z(new_n661_));
  OAI21_X1  g460(.A(new_n646_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(KEYINPUT46), .ZN(new_n663_));
  INV_X1    g462(.A(new_n661_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n659_), .A2(G36gat), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT112), .B(new_n664_), .C1(new_n665_), .C2(new_n658_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n662_), .A2(new_n663_), .A3(new_n666_), .ZN(G1329gat));
  NAND4_X1  g466(.A1(new_n634_), .A2(new_n640_), .A3(G43gat), .A4(new_n354_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G43gat), .B1(new_n623_), .B2(new_n354_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT113), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g471(.A(new_n450_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n634_), .A2(new_n640_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT114), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n675_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(G50gat), .A3(new_n677_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n613_), .A2(G50gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n624_), .B2(new_n679_), .ZN(G1331gat));
  NOR2_X1   g479(.A1(new_n569_), .A2(new_n583_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n543_), .A2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G57gat), .B1(new_n683_), .B2(new_n587_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n590_), .A2(new_n681_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(new_n265_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n686_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g486(.A(G64gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n683_), .A2(new_n688_), .A3(new_n597_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n597_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G64gat), .B1(new_n685_), .B2(new_n690_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n691_), .A2(KEYINPUT116), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(KEYINPUT116), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n689_), .B1(new_n695_), .B2(new_n696_), .ZN(G1333gat));
  OAI21_X1  g496(.A(G71gat), .B1(new_n685_), .B2(new_n424_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT49), .ZN(new_n699_));
  INV_X1    g498(.A(new_n683_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n424_), .A2(G71gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT117), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n699_), .B1(new_n700_), .B2(new_n702_), .ZN(G1334gat));
  OR3_X1    g502(.A1(new_n700_), .A2(G78gat), .A3(new_n613_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G78gat), .B1(new_n685_), .B2(new_n613_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(KEYINPUT50), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(KEYINPUT50), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT118), .ZN(G1335gat));
  INV_X1    g508(.A(KEYINPUT119), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n639_), .A2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n682_), .A2(new_n487_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n637_), .A2(KEYINPUT119), .A3(new_n638_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n711_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G85gat), .B1(new_n714_), .B2(new_n265_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n647_), .A2(new_n712_), .ZN(new_n716_));
  OR3_X1    g515(.A1(new_n716_), .A2(G85gat), .A3(new_n586_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT120), .ZN(G1336gat));
  INV_X1    g518(.A(KEYINPUT67), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G92gat), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n690_), .B(new_n714_), .C1(new_n506_), .C2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n716_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G92gat), .B1(new_n723_), .B2(new_n597_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1337gat));
  OAI21_X1  g524(.A(G99gat), .B1(new_n714_), .B2(new_n424_), .ZN(new_n726_));
  OR3_X1    g525(.A1(new_n716_), .A2(new_n511_), .A3(new_n424_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g528(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT52), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n639_), .A2(new_n673_), .A3(new_n712_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(G106gat), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(new_n731_), .A3(G106gat), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OR3_X1    g535(.A1(new_n716_), .A2(new_n512_), .A3(new_n450_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n730_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n735_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n737_), .B(new_n730_), .C1(new_n739_), .C2(new_n733_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n738_), .A2(new_n741_), .ZN(G1339gat));
  INV_X1    g541(.A(KEYINPUT57), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n745_), .A2(new_n552_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n552_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n561_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n748_), .A2(KEYINPUT56), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT56), .ZN(new_n750_));
  AOI211_X1 g549(.A(new_n750_), .B(new_n561_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n583_), .B(new_n564_), .C1(new_n749_), .C2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n574_), .A2(new_n572_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n571_), .B(KEYINPUT122), .Z(new_n754_));
  OAI211_X1 g553(.A(new_n579_), .B(new_n753_), .C1(new_n754_), .C2(new_n572_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(new_n580_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n565_), .A2(new_n756_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n752_), .A2(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(KEYINPUT123), .B(new_n743_), .C1(new_n758_), .C2(new_n539_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n539_), .B1(new_n752_), .B2(new_n757_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT123), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT57), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT124), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n746_), .A2(new_n747_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n562_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n766_), .B2(new_n750_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n751_), .A2(KEYINPUT124), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT125), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(new_n769_), .A3(new_n750_), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT125), .B1(new_n748_), .B2(KEYINPUT56), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n767_), .A2(new_n768_), .A3(new_n770_), .A4(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n756_), .A2(new_n564_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n772_), .A2(KEYINPUT58), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT58), .B1(new_n772_), .B2(new_n773_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n542_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n486_), .B1(new_n763_), .B2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n542_), .A2(new_n582_), .A3(new_n569_), .A4(new_n487_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT54), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n597_), .A2(new_n356_), .A3(new_n586_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(G113gat), .B1(new_n783_), .B2(new_n583_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(KEYINPUT126), .A3(KEYINPUT59), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT59), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT126), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n782_), .B2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n582_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n784_), .B1(new_n789_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g589(.A(G120gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n569_), .B2(KEYINPUT60), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n783_), .B(new_n792_), .C1(KEYINPUT60), .C2(new_n791_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n569_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(new_n791_), .ZN(G1341gat));
  AOI21_X1  g594(.A(G127gat), .B1(new_n783_), .B2(new_n487_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n486_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g597(.A(G134gat), .B1(new_n783_), .B2(new_n539_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n542_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(G134gat), .ZN(G1343gat));
  AOI21_X1  g600(.A(new_n430_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n597_), .A2(new_n586_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n583_), .ZN(new_n805_));
  XOR2_X1   g604(.A(KEYINPUT127), .B(G141gat), .Z(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1344gat));
  INV_X1    g606(.A(new_n569_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n804_), .A2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g609(.A1(new_n804_), .A2(new_n487_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(KEYINPUT61), .B(G155gat), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n811_), .B(new_n812_), .ZN(G1346gat));
  AOI21_X1  g612(.A(G162gat), .B1(new_n804_), .B2(new_n539_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n627_), .A2(G162gat), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n804_), .B2(new_n815_), .ZN(G1347gat));
  AOI21_X1  g615(.A(new_n690_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n817_), .A2(new_n354_), .A3(new_n586_), .A4(new_n613_), .ZN(new_n818_));
  OAI21_X1  g617(.A(G169gat), .B1(new_n818_), .B2(new_n582_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT62), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n818_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n583_), .A3(new_n327_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT62), .B(G169gat), .C1(new_n818_), .C2(new_n582_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(new_n823_), .A3(new_n824_), .ZN(G1348gat));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n808_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n356_), .ZN(new_n827_));
  AND4_X1   g626(.A1(G176gat), .A2(new_n817_), .A3(new_n827_), .A4(new_n586_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n826_), .A2(new_n326_), .B1(new_n828_), .B2(new_n808_), .ZN(G1349gat));
  NOR3_X1   g628(.A1(new_n818_), .A2(new_n368_), .A3(new_n486_), .ZN(new_n830_));
  INV_X1    g629(.A(G183gat), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n817_), .A2(new_n827_), .A3(new_n487_), .A4(new_n586_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n830_), .B1(new_n831_), .B2(new_n832_), .ZN(G1350gat));
  OAI21_X1  g632(.A(G190gat), .B1(new_n818_), .B2(new_n542_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n539_), .A2(new_n369_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n818_), .B2(new_n835_), .ZN(G1351gat));
  AND2_X1   g635(.A1(new_n802_), .A2(new_n265_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n583_), .A3(new_n597_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n808_), .A3(new_n597_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g640(.A(KEYINPUT63), .B(G211gat), .Z(new_n842_));
  AND4_X1   g641(.A1(new_n597_), .A2(new_n837_), .A3(new_n487_), .A4(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n837_), .A2(new_n597_), .A3(new_n487_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(G1354gat));
  AND3_X1   g645(.A1(new_n837_), .A2(G218gat), .A3(new_n597_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n837_), .A2(new_n539_), .A3(new_n597_), .ZN(new_n848_));
  INV_X1    g647(.A(G218gat), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n847_), .A2(new_n627_), .B1(new_n848_), .B2(new_n849_), .ZN(G1355gat));
endmodule


