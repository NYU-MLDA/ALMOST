//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G15gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT77), .B(G43gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G99gat), .Z(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT23), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n209_), .B1(G183gat), .B2(G190gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(G169gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n208_), .B(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(KEYINPUT24), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n215_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT26), .B(G190gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n221_), .A2(new_n222_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT76), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n220_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n221_), .A2(new_n222_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n224_), .A2(new_n225_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(KEYINPUT76), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n213_), .B1(new_n228_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT30), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n207_), .B1(new_n235_), .B2(KEYINPUT78), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(KEYINPUT78), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n236_), .B(new_n237_), .Z(new_n238_));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G113gat), .B(G120gat), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n240_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT80), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(KEYINPUT80), .A3(new_n242_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n247_), .A2(KEYINPUT31), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(KEYINPUT31), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n248_), .A2(KEYINPUT79), .A3(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n238_), .B(new_n250_), .Z(new_n251_));
  NOR2_X1   g050(.A1(G155gat), .A2(G162gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G155gat), .A2(G162gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n252_), .B1(KEYINPUT1), .B2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(KEYINPUT1), .B2(new_n253_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G141gat), .A2(G148gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT82), .ZN(new_n260_));
  XOR2_X1   g059(.A(G155gat), .B(G162gat), .Z(new_n261_));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n256_), .A2(KEYINPUT81), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT2), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n264_), .B1(G141gat), .B2(G148gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n258_), .A2(KEYINPUT2), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n263_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n268_));
  NOR3_X1   g067(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n268_), .B1(new_n269_), .B2(KEYINPUT81), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n260_), .B(new_n261_), .C1(new_n267_), .C2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G141gat), .ZN(new_n273_));
  INV_X1    g072(.A(G148gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n262_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT81), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n258_), .A2(KEYINPUT2), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n264_), .A2(G141gat), .A3(G148gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n277_), .A2(new_n280_), .A3(new_n268_), .A4(new_n263_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n260_), .B1(new_n281_), .B2(new_n261_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n259_), .B(new_n243_), .C1(new_n272_), .C2(new_n282_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n255_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n261_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT82), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n284_), .B1(new_n286_), .B2(new_n271_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n245_), .A2(new_n246_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n283_), .B(KEYINPUT4), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G225gat), .A2(G233gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n259_), .B1(new_n272_), .B2(new_n282_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n247_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n289_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G1gat), .B(G29gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G57gat), .B(G85gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n283_), .B(new_n290_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n295_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n301_), .B1(new_n295_), .B2(new_n302_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT98), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  AOI211_X1 g105(.A(KEYINPUT98), .B(new_n301_), .C1(new_n295_), .C2(new_n302_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n251_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT19), .ZN(new_n311_));
  INV_X1    g110(.A(G211gat), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n312_), .A2(G218gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(G218gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G197gat), .A2(G204gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(KEYINPUT86), .B(G197gat), .Z(new_n319_));
  INV_X1    g118(.A(G204gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT21), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n316_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(KEYINPUT86), .A2(G197gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(KEYINPUT86), .A2(G197gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n320_), .A3(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n322_), .B1(G197gat), .B2(G204gat), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n326_), .A2(KEYINPUT87), .A3(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT87), .B1(new_n326_), .B2(new_n327_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT21), .B1(new_n313_), .B2(new_n314_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n324_), .A2(new_n325_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n317_), .B1(new_n332_), .B2(G204gat), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n333_), .B2(KEYINPUT88), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT88), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n320_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n335_), .B1(new_n336_), .B2(new_n317_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n323_), .A2(new_n330_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT90), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT25), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n340_), .A2(G183gat), .ZN(new_n341_));
  INV_X1    g140(.A(G183gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n342_), .A2(KEYINPUT25), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n339_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(KEYINPUT25), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(G183gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(KEYINPUT90), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n344_), .A2(new_n347_), .A3(new_n222_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n348_), .A2(KEYINPUT91), .A3(new_n230_), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT91), .B1(new_n348_), .B2(new_n230_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n220_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT92), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n210_), .A2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n209_), .B(KEYINPUT92), .C1(G183gat), .C2(G190gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(new_n212_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n338_), .B1(new_n351_), .B2(new_n355_), .ZN(new_n356_));
  OAI211_X1 g155(.A(KEYINPUT88), .B(new_n318_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n331_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(new_n337_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n326_), .A2(new_n327_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT87), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n326_), .A2(KEYINPUT87), .A3(new_n327_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n315_), .B1(new_n333_), .B2(KEYINPUT21), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n359_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT20), .B1(new_n233_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n311_), .B1(new_n356_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n351_), .A2(new_n338_), .A3(new_n355_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT20), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n233_), .B2(new_n366_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n311_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n369_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT18), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n377_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n380_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n368_), .A2(new_n373_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT27), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n367_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n351_), .A2(new_n355_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n387_), .B(new_n372_), .C1(new_n388_), .C2(new_n338_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n369_), .A2(new_n371_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n311_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n380_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(KEYINPUT27), .A3(new_n383_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n386_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n287_), .A2(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n398_), .A2(KEYINPUT28), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(KEYINPUT28), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G22gat), .B(G50gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n401_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT83), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n399_), .A2(new_n400_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n401_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT83), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n402_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n405_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT89), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n338_), .A2(KEYINPUT85), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n397_), .B2(new_n287_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(KEYINPUT84), .A2(G233gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(KEYINPUT84), .A2(G233gat), .ZN(new_n419_));
  OAI21_X1  g218(.A(G228gat), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n415_), .B(new_n420_), .C1(new_n397_), .C2(new_n287_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n414_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n424_), .A3(new_n413_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n427_), .A2(new_n408_), .A3(new_n402_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n412_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n411_), .A2(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n396_), .A2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n309_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n283_), .B(new_n291_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n434_), .A2(new_n300_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n289_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n295_), .A2(KEYINPUT33), .A3(new_n301_), .A4(new_n302_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n302_), .A2(new_n301_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n294_), .A2(new_n291_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n439_), .B1(new_n289_), .B2(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n437_), .B(new_n438_), .C1(new_n441_), .C2(KEYINPUT33), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT94), .B1(new_n442_), .B2(new_n384_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n368_), .A2(new_n373_), .A3(new_n382_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n382_), .B1(new_n368_), .B2(new_n373_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT94), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT33), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n303_), .A2(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n302_), .A2(KEYINPUT33), .A3(new_n301_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n450_), .A2(new_n295_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n446_), .A2(new_n447_), .A3(new_n449_), .A4(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n378_), .A2(KEYINPUT32), .A3(new_n379_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT95), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n368_), .A2(new_n373_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT96), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n368_), .A2(KEYINPUT96), .A3(new_n455_), .A4(new_n373_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n453_), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT97), .B1(new_n392_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT97), .ZN(new_n463_));
  AOI211_X1 g262(.A(new_n463_), .B(new_n453_), .C1(new_n389_), .C2(new_n391_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n460_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n443_), .B(new_n452_), .C1(new_n465_), .C2(new_n308_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n431_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT99), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT99), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n466_), .A2(new_n469_), .A3(new_n431_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n308_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n431_), .A2(new_n471_), .A3(new_n395_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n468_), .A2(new_n470_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n251_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n433_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT14), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT70), .B(G1gat), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n477_), .B1(new_n478_), .B2(G8gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT71), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT71), .ZN(new_n481_));
  INV_X1    g280(.A(G8gat), .ZN(new_n482_));
  OR2_X1    g281(.A1(KEYINPUT70), .A2(G1gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(KEYINPUT70), .A2(G1gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n482_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n481_), .B1(new_n485_), .B2(new_n477_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n480_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n487_), .A2(KEYINPUT72), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT72), .B1(new_n487_), .B2(new_n488_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G8gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n489_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n486_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n485_), .A2(new_n481_), .A3(new_n477_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n488_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT72), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n487_), .A2(KEYINPUT72), .A3(new_n488_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n491_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n493_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G29gat), .B(G36gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT68), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G43gat), .B(G50gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT15), .ZN(new_n506_));
  INV_X1    g305(.A(new_n504_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n503_), .B(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT15), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n501_), .A2(new_n506_), .A3(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n492_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n498_), .A2(new_n499_), .A3(new_n491_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n508_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n511_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n516_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n512_), .A2(new_n513_), .A3(new_n505_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n505_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n518_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G113gat), .B(G141gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT74), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G169gat), .B(G197gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n525_), .B(new_n526_), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n517_), .A2(new_n522_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT75), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n531_), .A2(new_n532_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n476_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G230gat), .A2(G233gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G57gat), .B(G64gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n542_));
  XOR2_X1   g341(.A(G71gat), .B(G78gat), .Z(new_n543_));
  OR2_X1    g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n543_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(KEYINPUT10), .B(G99gat), .Z(new_n548_));
  INV_X1    g347(.A(G106gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G85gat), .B(G92gat), .Z(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT9), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT9), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(G85gat), .A3(G92gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G99gat), .A2(G106gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT6), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n550_), .A2(new_n552_), .A3(new_n554_), .A4(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT7), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT6), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n555_), .B(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n551_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n563_), .A2(KEYINPUT8), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G85gat), .B(G92gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n558_), .B(KEYINPUT7), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n565_), .B1(new_n566_), .B2(new_n556_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT8), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n547_), .B(new_n557_), .C1(new_n564_), .C2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT64), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n557_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n563_), .A2(KEYINPUT8), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n567_), .A2(new_n568_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(new_n547_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n540_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n576_), .A2(KEYINPUT12), .A3(new_n547_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT12), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n557_), .B1(new_n564_), .B2(new_n569_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n547_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n580_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n539_), .B(new_n570_), .C1(new_n579_), .C2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n578_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G120gat), .B(G148gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G176gat), .B(G204gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT65), .B(KEYINPUT5), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n585_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT13), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n592_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT66), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n506_), .A2(new_n510_), .A3(new_n581_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n576_), .A2(new_n508_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT35), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n597_), .A2(new_n598_), .A3(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n601_), .A2(new_n602_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(KEYINPUT36), .ZN(new_n610_));
  INV_X1    g409(.A(new_n605_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n597_), .A2(new_n598_), .A3(new_n611_), .A4(new_n603_), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n606_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n609_), .B(KEYINPUT36), .Z(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n606_), .B2(new_n612_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT37), .B1(new_n617_), .B2(KEYINPUT69), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT69), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT37), .ZN(new_n620_));
  NOR4_X1   g419(.A1(new_n613_), .A2(new_n616_), .A3(new_n619_), .A4(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(G231gat), .ZN(new_n623_));
  INV_X1    g422(.A(G233gat), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n514_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n514_), .A2(new_n625_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n547_), .B(KEYINPUT73), .Z(new_n628_));
  OR3_X1    g427(.A1(new_n626_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(G127gat), .B(G155gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT16), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G183gat), .B(G211gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT17), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n628_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n629_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n633_), .A2(new_n634_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n629_), .B2(new_n636_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n622_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n596_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n538_), .A2(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n644_), .A2(new_n308_), .A3(new_n478_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n645_), .A2(KEYINPUT38), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(KEYINPUT38), .ZN(new_n647_));
  INV_X1    g446(.A(new_n617_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n593_), .A2(new_n594_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(new_n531_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(new_n640_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n472_), .B1(new_n467_), .B2(KEYINPUT99), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n251_), .B1(new_n652_), .B2(new_n470_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n648_), .B(new_n651_), .C1(new_n653_), .C2(new_n433_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G1gat), .B1(new_n654_), .B2(new_n308_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n646_), .A2(new_n647_), .A3(new_n655_), .ZN(G1324gat));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n476_), .A2(new_n617_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n395_), .A3(new_n651_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n657_), .B1(new_n659_), .B2(G8gat), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n657_), .B(G8gat), .C1(new_n654_), .C2(new_n396_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n395_), .A2(new_n482_), .ZN(new_n663_));
  OAI22_X1  g462(.A1(new_n660_), .A2(new_n662_), .B1(new_n644_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT101), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n666_));
  OAI221_X1 g465(.A(new_n666_), .B1(new_n644_), .B2(new_n663_), .C1(new_n660_), .C2(new_n662_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n665_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1325gat));
  INV_X1    g470(.A(G15gat), .ZN(new_n672_));
  INV_X1    g471(.A(new_n654_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n673_), .B2(new_n251_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT102), .B(KEYINPUT41), .Z(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n538_), .A2(new_n672_), .A3(new_n251_), .A4(new_n643_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n674_), .A2(new_n675_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT103), .Z(G1326gat));
  OAI21_X1  g480(.A(G22gat), .B1(new_n654_), .B2(new_n431_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT42), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n431_), .A2(G22gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n644_), .B2(new_n684_), .ZN(G1327gat));
  NAND2_X1  g484(.A1(new_n640_), .A2(new_n617_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n595_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n538_), .A2(new_n687_), .ZN(new_n688_));
  OR3_X1    g487(.A1(new_n688_), .A2(G29gat), .A3(new_n308_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n622_), .B(KEYINPUT104), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT43), .B1(new_n476_), .B2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n622_), .A2(KEYINPUT43), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT105), .B1(new_n476_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n695_), .B(new_n692_), .C1(new_n653_), .C2(new_n433_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n691_), .A2(new_n694_), .A3(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n650_), .A2(new_n641_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n697_), .A2(new_n702_), .A3(new_n698_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(KEYINPUT107), .A3(new_n471_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G29gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT107), .B1(new_n704_), .B2(new_n471_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n689_), .B1(new_n706_), .B2(new_n707_), .ZN(G1328gat));
  INV_X1    g507(.A(new_n688_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n396_), .A2(G36gat), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT45), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n396_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n713_));
  INV_X1    g512(.A(G36gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n712_), .B(KEYINPUT46), .C1(new_n713_), .C2(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1329gat));
  INV_X1    g518(.A(G43gat), .ZN(new_n720_));
  AOI211_X1 g519(.A(new_n720_), .B(new_n475_), .C1(new_n701_), .C2(new_n703_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT108), .B(G43gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n709_), .B2(new_n251_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT47), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n475_), .A2(new_n720_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n723_), .B1(new_n704_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n724_), .A2(new_n728_), .ZN(G1330gat));
  INV_X1    g528(.A(new_n431_), .ZN(new_n730_));
  AOI21_X1  g529(.A(G50gat), .B1(new_n709_), .B2(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n730_), .A2(G50gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n704_), .B2(new_n732_), .ZN(G1331gat));
  XNOR2_X1  g532(.A(new_n649_), .B(KEYINPUT66), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n641_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n658_), .A2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n308_), .ZN(new_n738_));
  NOR4_X1   g537(.A1(new_n476_), .A2(new_n531_), .A3(new_n649_), .A4(new_n642_), .ZN(new_n739_));
  INV_X1    g538(.A(G57gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n471_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n741_), .ZN(G1332gat));
  OAI21_X1  g541(.A(G64gat), .B1(new_n737_), .B2(new_n396_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT48), .ZN(new_n744_));
  INV_X1    g543(.A(G64gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n739_), .A2(new_n745_), .A3(new_n395_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n737_), .B2(new_n475_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT49), .ZN(new_n749_));
  INV_X1    g548(.A(G71gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n739_), .A2(new_n750_), .A3(new_n251_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1334gat));
  INV_X1    g551(.A(G78gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n739_), .A2(new_n753_), .A3(new_n730_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n658_), .A2(new_n736_), .A3(new_n730_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(G78gat), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n755_), .B2(G78gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n754_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT109), .Z(G1335gat));
  INV_X1    g560(.A(G85gat), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n476_), .A2(new_n531_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n734_), .A2(new_n686_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n762_), .B1(new_n765_), .B2(new_n308_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT110), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n649_), .A2(new_n531_), .A3(new_n641_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n697_), .A2(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n308_), .A2(new_n762_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n767_), .B1(new_n769_), .B2(new_n770_), .ZN(G1336gat));
  NOR3_X1   g570(.A1(new_n765_), .A2(G92gat), .A3(new_n396_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n697_), .A2(new_n395_), .A3(new_n768_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(G92gat), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n774_), .B(KEYINPUT111), .Z(G1337gat));
  AND4_X1   g574(.A1(new_n251_), .A2(new_n763_), .A3(new_n548_), .A4(new_n764_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT112), .Z(new_n777_));
  NAND2_X1  g576(.A1(new_n769_), .A2(new_n251_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G99gat), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(KEYINPUT113), .A3(KEYINPUT51), .ZN(new_n781_));
  NAND2_X1  g580(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n777_), .A2(new_n779_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1338gat));
  XNOR2_X1  g583(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n697_), .A2(new_n730_), .A3(new_n768_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(G106gat), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT52), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n789_), .A3(G106gat), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n763_), .A2(new_n764_), .A3(new_n549_), .A4(new_n730_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n785_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n786_), .A2(new_n789_), .A3(G106gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n789_), .B1(new_n786_), .B2(G106gat), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n792_), .B(new_n785_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n793_), .A2(new_n797_), .ZN(G1339gat));
  INV_X1    g597(.A(KEYINPUT58), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n584_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n579_), .A2(new_n583_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n540_), .B1(new_n803_), .B2(new_n572_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n570_), .A2(new_n539_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT12), .B1(new_n576_), .B2(new_n547_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n581_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n805_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT115), .B1(new_n808_), .B2(KEYINPUT55), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(KEYINPUT55), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n802_), .A2(new_n804_), .A3(new_n809_), .A4(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n590_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT56), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n585_), .A2(new_n590_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n811_), .A2(new_n815_), .A3(new_n590_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n813_), .A2(new_n814_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n518_), .B1(new_n515_), .B2(new_n519_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT116), .B1(new_n818_), .B2(new_n529_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n516_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n527_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n511_), .A2(new_n515_), .A3(new_n518_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n819_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n530_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n799_), .B1(new_n817_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n816_), .A2(new_n814_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n815_), .B1(new_n811_), .B2(new_n590_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n825_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(KEYINPUT58), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n622_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n826_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n813_), .A2(new_n531_), .A3(new_n814_), .A4(new_n816_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n591_), .A2(new_n530_), .A3(new_n824_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n617_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT57), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n833_), .A2(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n640_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n535_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n640_), .B1(new_n842_), .B2(new_n533_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n843_), .A2(new_n649_), .A3(new_n844_), .A4(new_n622_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n622_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT54), .B1(new_n735_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n841_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n475_), .A2(new_n308_), .A3(new_n432_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n836_), .A2(new_n839_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n853_), .A2(KEYINPUT118), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(KEYINPUT118), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n838_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n848_), .B1(new_n856_), .B2(new_n641_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n857_), .A2(new_n851_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n852_), .B1(new_n858_), .B2(new_n850_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G113gat), .B1(new_n859_), .B2(new_n537_), .ZN(new_n860_));
  INV_X1    g659(.A(G113gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n858_), .A2(new_n861_), .A3(new_n531_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1340gat));
  OAI21_X1  g662(.A(G120gat), .B1(new_n859_), .B2(new_n734_), .ZN(new_n864_));
  INV_X1    g663(.A(G120gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n649_), .B2(KEYINPUT60), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n858_), .B(new_n866_), .C1(KEYINPUT60), .C2(new_n865_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(G1341gat));
  OAI21_X1  g667(.A(G127gat), .B1(new_n859_), .B2(new_n640_), .ZN(new_n869_));
  INV_X1    g668(.A(G127gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n858_), .A2(new_n870_), .A3(new_n641_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1342gat));
  OAI21_X1  g671(.A(G134gat), .B1(new_n859_), .B2(new_n622_), .ZN(new_n873_));
  INV_X1    g672(.A(G134gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n858_), .A2(new_n874_), .A3(new_n617_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1343gat));
  NOR4_X1   g675(.A1(new_n251_), .A2(new_n431_), .A3(new_n308_), .A4(new_n395_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n857_), .A2(KEYINPUT119), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT119), .B1(new_n857_), .B2(new_n877_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n531_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g680(.A(new_n596_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g682(.A(new_n641_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT61), .B(G155gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1346gat));
  OR2_X1    g685(.A1(new_n878_), .A2(new_n879_), .ZN(new_n887_));
  INV_X1    g686(.A(G162gat), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n690_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n617_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n887_), .A2(new_n889_), .B1(new_n890_), .B2(new_n888_), .ZN(G1347gat));
  OR3_X1    g690(.A1(new_n309_), .A2(KEYINPUT120), .A3(new_n396_), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT120), .B1(new_n309_), .B2(new_n396_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n730_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n827_), .A2(new_n825_), .A3(new_n828_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n622_), .B1(new_n895_), .B2(KEYINPUT58), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n896_), .A2(new_n826_), .B1(KEYINPUT57), .B2(new_n836_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n641_), .B1(new_n897_), .B2(new_n853_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n845_), .A2(new_n847_), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n531_), .B(new_n894_), .C1(new_n898_), .C2(new_n899_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT22), .B(G169gat), .Z(new_n901_));
  OR2_X1    g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n900_), .A2(KEYINPUT121), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n849_), .A2(new_n905_), .A3(new_n531_), .A4(new_n894_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n216_), .B1(KEYINPUT122), .B2(KEYINPUT62), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n903_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n903_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n908_), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n910_), .B(new_n911_), .C1(new_n904_), .C2(new_n906_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n902_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT123), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n915_), .B(new_n902_), .C1(new_n909_), .C2(new_n912_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1348gat));
  NAND2_X1  g716(.A1(new_n849_), .A2(new_n894_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G176gat), .B1(new_n919_), .B2(new_n595_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n857_), .A2(new_n431_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n892_), .A2(new_n893_), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n922_), .A2(G176gat), .A3(new_n596_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n920_), .B1(new_n921_), .B2(new_n923_), .ZN(G1349gat));
  AOI211_X1 g723(.A(new_n640_), .B(new_n918_), .C1(new_n344_), .C2(new_n347_), .ZN(new_n925_));
  AND4_X1   g724(.A1(new_n431_), .A2(new_n857_), .A3(new_n641_), .A4(new_n922_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n926_), .A2(KEYINPUT124), .ZN(new_n927_));
  AOI21_X1  g726(.A(G183gat), .B1(new_n926_), .B2(KEYINPUT124), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n925_), .B1(new_n927_), .B2(new_n928_), .ZN(G1350gat));
  OAI21_X1  g728(.A(G190gat), .B1(new_n918_), .B2(new_n622_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n617_), .A2(new_n222_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n918_), .B2(new_n931_), .ZN(G1351gat));
  NOR4_X1   g731(.A1(new_n251_), .A2(new_n431_), .A3(new_n471_), .A4(new_n396_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n857_), .A2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n531_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g736(.A1(new_n934_), .A2(new_n734_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n320_), .ZN(G1353gat));
  AOI21_X1  g738(.A(new_n640_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(KEYINPUT125), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n935_), .A2(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  XOR2_X1   g742(.A(new_n942_), .B(new_n943_), .Z(G1354gat));
  NOR3_X1   g743(.A1(new_n934_), .A2(KEYINPUT126), .A3(new_n648_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(G218gat), .ZN(new_n946_));
  OAI21_X1  g745(.A(KEYINPUT126), .B1(new_n934_), .B2(new_n648_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n832_), .A2(G218gat), .ZN(new_n948_));
  XOR2_X1   g747(.A(new_n948_), .B(KEYINPUT127), .Z(new_n949_));
  AOI22_X1  g748(.A1(new_n946_), .A2(new_n947_), .B1(new_n935_), .B2(new_n949_), .ZN(G1355gat));
endmodule


