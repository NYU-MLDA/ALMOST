//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G1gat), .B(G8gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT71), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G15gat), .ZN(new_n209_));
  INV_X1    g008(.A(G22gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G15gat), .A2(G22gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G1gat), .A2(G8gat), .ZN(new_n213_));
  AOI22_X1  g012(.A1(new_n211_), .A2(new_n212_), .B1(KEYINPUT14), .B2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n208_), .B(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G43gat), .B(G50gat), .Z(new_n217_));
  INV_X1    g016(.A(G36gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G29gat), .ZN(new_n219_));
  INV_X1    g018(.A(G29gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G36gat), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT68), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT68), .B1(new_n219_), .B2(new_n221_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n217_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n220_), .A2(G36gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n218_), .A2(G29gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT68), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G43gat), .B(G50gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n224_), .A2(KEYINPUT15), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT15), .B1(new_n224_), .B2(new_n231_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n216_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n224_), .A2(new_n231_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT73), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n236_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n215_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n234_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n239_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n216_), .B1(new_n237_), .B2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n241_), .B1(new_n244_), .B2(new_n240_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n205_), .B1(new_n242_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n241_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n240_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n215_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n234_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(new_n204_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(new_n252_), .A3(KEYINPUT74), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT74), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n254_), .B(new_n205_), .C1(new_n242_), .C2(new_n245_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(KEYINPUT67), .B(KEYINPUT34), .Z(new_n258_));
  NAND2_X1  g057(.A1(G232gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT35), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n264_));
  INV_X1    g063(.A(G106gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(G85gat), .A2(G92gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G85gat), .A2(G92gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(KEYINPUT9), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G99gat), .A2(G106gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT6), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(G99gat), .A3(G106gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n269_), .A2(KEYINPUT9), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n267_), .A2(new_n270_), .A3(new_n275_), .A4(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n268_), .A2(new_n269_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT65), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n281_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT7), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G99gat), .A2(G106gat), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n272_), .A2(new_n274_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n278_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n277_), .B1(new_n287_), .B2(KEYINPUT8), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n284_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n275_), .A2(new_n289_), .A3(new_n280_), .A4(new_n282_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n278_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT8), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  OAI22_X1  g093(.A1(new_n288_), .A2(new_n294_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n263_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  AND4_X1   g096(.A1(new_n275_), .A2(new_n267_), .A3(new_n270_), .A4(new_n276_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n298_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n287_), .A2(KEYINPUT8), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n299_), .A2(new_n231_), .A3(new_n224_), .A4(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n295_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n260_), .A2(new_n261_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n295_), .A2(new_n301_), .A3(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n297_), .A2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT70), .B1(new_n304_), .B2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G190gat), .B(G218gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G134gat), .B(G162gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(KEYINPUT36), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n304_), .A2(new_n307_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(KEYINPUT36), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n308_), .B(new_n313_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n295_), .A2(new_n301_), .A3(new_n305_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT15), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n222_), .A2(new_n223_), .A3(new_n217_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n230_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n319_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n224_), .A2(new_n231_), .A3(KEYINPUT15), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n299_), .A2(new_n300_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n262_), .B1(new_n324_), .B2(KEYINPUT69), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n318_), .A2(new_n325_), .ZN(new_n326_));
  AOI221_X4 g125(.A(new_n317_), .B1(new_n313_), .B2(new_n315_), .C1(new_n326_), .C2(new_n303_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n316_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(G183gat), .A3(G190gat), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n331_), .A2(KEYINPUT76), .ZN(new_n332_));
  INV_X1    g131(.A(G183gat), .ZN(new_n333_));
  INV_X1    g132(.A(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT23), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(new_n331_), .A3(KEYINPUT76), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n332_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(G169gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT25), .B(G183gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT26), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G190gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n334_), .A2(KEYINPUT26), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n344_), .A2(KEYINPUT75), .A3(G190gat), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n343_), .A2(new_n347_), .A3(new_n348_), .A4(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n337_), .A2(new_n331_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G169gat), .A2(G176gat), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n352_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n350_), .A2(new_n351_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n342_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT30), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G15gat), .B(G43gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT77), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(G99gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G227gat), .A2(G233gat), .ZN(new_n364_));
  INV_X1    g163(.A(G71gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n363_), .B(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n360_), .B1(new_n367_), .B2(KEYINPUT78), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n358_), .A2(new_n359_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n368_), .B(new_n369_), .C1(KEYINPUT78), .C2(new_n367_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n367_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n372_));
  INV_X1    g171(.A(new_n369_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n371_), .B(new_n372_), .C1(new_n373_), .C2(new_n360_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n370_), .A2(KEYINPUT80), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n376_));
  INV_X1    g175(.A(G134gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G127gat), .ZN(new_n378_));
  INV_X1    g177(.A(G127gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G134gat), .ZN(new_n380_));
  INV_X1    g179(.A(G120gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G113gat), .ZN(new_n382_));
  INV_X1    g181(.A(G113gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G120gat), .ZN(new_n384_));
  AND4_X1   g183(.A1(new_n378_), .A2(new_n380_), .A3(new_n382_), .A4(new_n384_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n378_), .A2(new_n380_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n376_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n378_), .A2(new_n380_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n382_), .A2(new_n384_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n378_), .A2(new_n380_), .A3(new_n382_), .A4(new_n384_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(KEYINPUT79), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n387_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT31), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n375_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397_));
  INV_X1    g196(.A(G141gat), .ZN(new_n398_));
  INV_X1    g197(.A(G148gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G141gat), .A2(G148gat), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT2), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n400_), .A2(new_n403_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G155gat), .B(G162gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(G141gat), .A2(G148gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(G141gat), .A2(G148gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n412_), .B(new_n413_), .C1(new_n407_), .C2(KEYINPUT1), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT82), .B1(new_n415_), .B2(KEYINPUT29), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G211gat), .B(G218gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT21), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(G204gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G197gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT83), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n420_), .A3(G197gat), .ZN(new_n424_));
  INV_X1    g223(.A(G197gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(G204gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n419_), .A2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n422_), .A2(new_n424_), .A3(new_n418_), .A4(new_n426_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n421_), .A2(new_n426_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT21), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n417_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n428_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n416_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G228gat), .ZN(new_n436_));
  INV_X1    g235(.A(G233gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n435_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n416_), .A2(new_n440_), .A3(new_n434_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G78gat), .B(G106gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT85), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G22gat), .B(G50gat), .Z(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(KEYINPUT81), .B(KEYINPUT28), .Z(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n415_), .B2(KEYINPUT29), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n415_), .A2(KEYINPUT29), .A3(new_n449_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n448_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n415_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT29), .ZN(new_n455_));
  INV_X1    g254(.A(new_n449_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n453_), .A2(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n439_), .A2(new_n441_), .A3(KEYINPUT85), .A4(new_n443_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n446_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n453_), .A2(new_n462_), .A3(new_n458_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n441_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n440_), .B1(new_n416_), .B2(new_n434_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n442_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n463_), .A2(new_n466_), .A3(new_n444_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n443_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n459_), .B2(KEYINPUT84), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n461_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT86), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n461_), .A2(new_n467_), .A3(new_n472_), .A4(new_n469_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G226gat), .A2(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n356_), .A2(new_n332_), .A3(new_n338_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n333_), .A2(KEYINPUT25), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n333_), .A2(KEYINPUT25), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n343_), .A2(KEYINPUT88), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n348_), .A2(new_n345_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT89), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n351_), .A2(new_n488_), .A3(new_n335_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n488_), .B1(new_n351_), .B2(new_n335_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n341_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n478_), .B1(new_n493_), .B2(new_n434_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G211gat), .B(G218gat), .Z(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(KEYINPUT21), .B2(new_n431_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n496_), .A2(new_n429_), .B1(new_n427_), .B2(new_n419_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(new_n342_), .A3(new_n357_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n477_), .B1(new_n494_), .B2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n487_), .A2(new_n497_), .A3(new_n492_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n358_), .A2(new_n434_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT20), .A4(new_n477_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G8gat), .B(G36gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G64gat), .B(G92gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n499_), .A2(new_n503_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n508_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n491_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n489_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n512_), .A2(new_n341_), .B1(new_n479_), .B2(new_n486_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n498_), .B(KEYINPUT20), .C1(new_n513_), .C2(new_n497_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n477_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n510_), .B1(new_n516_), .B2(new_n502_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n509_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT95), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(KEYINPUT33), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n415_), .A2(new_n387_), .A3(new_n392_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n409_), .B(new_n414_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(KEYINPUT91), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT91), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n415_), .A2(new_n387_), .A3(new_n524_), .A4(new_n392_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G225gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT92), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT94), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT94), .ZN(new_n531_));
  AOI211_X1 g330(.A(new_n531_), .B(new_n528_), .C1(new_n523_), .C2(new_n525_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G1gat), .B(G29gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(G85gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT0), .B(G57gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  INV_X1    g336(.A(KEYINPUT4), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n415_), .A2(new_n387_), .A3(new_n538_), .A4(new_n392_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT93), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n539_), .A2(new_n540_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n528_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n538_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n537_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n520_), .B1(new_n533_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n537_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n526_), .A2(KEYINPUT4), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n393_), .A2(KEYINPUT93), .A3(new_n538_), .A4(new_n415_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n539_), .A2(new_n540_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n529_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n547_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n520_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n552_), .B(new_n553_), .C1(new_n530_), .C2(new_n532_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n537_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n529_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n555_), .B1(new_n544_), .B2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n518_), .A2(new_n546_), .A3(new_n554_), .A4(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n543_), .A2(new_n544_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n547_), .B1(new_n533_), .B2(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n530_), .A2(new_n532_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n552_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n494_), .A2(new_n477_), .A3(new_n498_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n500_), .A2(new_n501_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n515_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n516_), .A2(new_n502_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n510_), .A2(KEYINPUT32), .ZN(new_n570_));
  MUX2_X1   g369(.A(new_n568_), .B(new_n569_), .S(new_n570_), .Z(new_n571_));
  AOI22_X1  g370(.A1(new_n558_), .A2(KEYINPUT96), .B1(new_n563_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n508_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n516_), .A2(new_n510_), .A3(new_n502_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n573_), .A2(new_n574_), .A3(new_n557_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT96), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n575_), .A2(new_n576_), .A3(new_n546_), .A4(new_n554_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n474_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT98), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n560_), .A2(new_n562_), .A3(new_n579_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT27), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n509_), .B2(new_n517_), .ZN(new_n584_));
  OAI211_X1 g383(.A(KEYINPUT27), .B(new_n574_), .C1(new_n568_), .C2(new_n510_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AND4_X1   g386(.A1(new_n581_), .A2(new_n474_), .A3(new_n582_), .A4(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n396_), .B1(new_n578_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n582_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(new_n580_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n474_), .A2(new_n586_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n395_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n329_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G57gat), .B(G64gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G71gat), .B(G78gat), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n596_), .A3(KEYINPUT11), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(KEYINPUT11), .ZN(new_n598_));
  INV_X1    g397(.A(new_n596_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n595_), .A2(KEYINPUT11), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n597_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n215_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT16), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT17), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n602_), .B(new_n603_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n216_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n605_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT72), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n605_), .A2(new_n613_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n609_), .B(KEYINPUT17), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n602_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n288_), .B2(new_n294_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n299_), .A2(new_n300_), .A3(new_n602_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(KEYINPUT12), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT12), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n625_), .B(new_n621_), .C1(new_n288_), .C2(new_n294_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT64), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT5), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n633_), .B(new_n634_), .Z(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n622_), .A2(new_n623_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n631_), .B(new_n636_), .C1(new_n630_), .C2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n630_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n629_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n635_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT13), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(KEYINPUT66), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n638_), .A2(new_n641_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n642_), .A2(KEYINPUT66), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n638_), .A2(new_n641_), .B1(new_n646_), .B2(new_n644_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AND4_X1   g448(.A1(new_n257_), .A2(new_n594_), .A3(new_n620_), .A4(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n581_), .A2(new_n582_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(G1gat), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT38), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n256_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n620_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n316_), .A2(KEYINPUT37), .A3(new_n328_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT37), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n315_), .B1(new_n326_), .B2(new_n303_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n317_), .B1(new_n326_), .B2(new_n303_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n312_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n662_), .B2(new_n327_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n657_), .B1(new_n658_), .B2(new_n663_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n656_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n653_), .A3(new_n651_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n654_), .B1(new_n655_), .B2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n667_), .B1(new_n655_), .B2(new_n666_), .ZN(G1324gat));
  INV_X1    g467(.A(G8gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n665_), .A2(new_n669_), .A3(new_n586_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n650_), .A2(new_n586_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT39), .ZN(new_n673_));
  AND4_X1   g472(.A1(new_n671_), .A2(new_n672_), .A3(new_n673_), .A4(G8gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n669_), .B1(KEYINPUT99), .B2(KEYINPUT39), .ZN(new_n675_));
  AOI22_X1  g474(.A1(new_n672_), .A2(new_n675_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n670_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(G1325gat));
  NAND2_X1  g478(.A1(new_n650_), .A2(new_n395_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G15gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT100), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n681_), .B(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT41), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n665_), .A2(new_n209_), .A3(new_n395_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n684_), .A2(new_n687_), .A3(new_n688_), .ZN(G1326gat));
  AOI21_X1  g488(.A(new_n210_), .B1(new_n650_), .B2(new_n474_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n665_), .A2(new_n210_), .A3(new_n474_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1327gat));
  INV_X1    g493(.A(new_n329_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n695_), .A2(new_n648_), .A3(new_n620_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n656_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n651_), .A2(new_n220_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT106), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n648_), .A2(new_n256_), .A3(new_n620_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT102), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n663_), .A2(new_n658_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(KEYINPUT103), .ZN(new_n706_));
  AOI211_X1 g505(.A(new_n704_), .B(new_n706_), .C1(new_n589_), .C2(new_n593_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n546_), .A2(new_n554_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n573_), .A2(new_n574_), .A3(new_n557_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT96), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n563_), .A2(new_n571_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n577_), .A3(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n474_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n586_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n715_));
  AOI22_X1  g514(.A1(new_n713_), .A2(new_n714_), .B1(new_n591_), .B2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n593_), .B1(new_n716_), .B2(new_n395_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n704_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n708_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n703_), .B1(new_n707_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723_));
  OAI211_X1 g522(.A(KEYINPUT44), .B(new_n703_), .C1(new_n707_), .C2(new_n719_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n722_), .A2(new_n723_), .A3(new_n651_), .A4(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(G29gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n722_), .A2(new_n651_), .A3(new_n724_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT104), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n701_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  AND4_X1   g528(.A1(new_n701_), .A2(new_n728_), .A3(G29gat), .A4(new_n725_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n700_), .B1(new_n729_), .B2(new_n730_), .ZN(G1328gat));
  NAND3_X1  g530(.A1(new_n697_), .A2(new_n218_), .A3(new_n586_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT45), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n717_), .B(new_n718_), .C1(KEYINPUT103), .C2(new_n705_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n704_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(new_n708_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT44), .B1(new_n736_), .B2(new_n703_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n724_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n587_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n733_), .B1(new_n739_), .B2(new_n218_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(G1329gat));
  NOR2_X1   g541(.A1(new_n737_), .A2(new_n738_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(G43gat), .A3(new_n395_), .ZN(new_n744_));
  INV_X1    g543(.A(G43gat), .ZN(new_n745_));
  INV_X1    g544(.A(new_n697_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(new_n396_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n744_), .A2(KEYINPUT47), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT47), .B1(new_n744_), .B2(new_n747_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1330gat));
  AOI21_X1  g549(.A(G50gat), .B1(new_n697_), .B2(new_n474_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n474_), .A2(G50gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n743_), .B2(new_n752_), .ZN(G1331gat));
  AOI21_X1  g552(.A(new_n257_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n754_));
  AND4_X1   g553(.A1(new_n704_), .A2(new_n754_), .A3(new_n620_), .A4(new_n648_), .ZN(new_n755_));
  INV_X1    g554(.A(G57gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n651_), .ZN(new_n757_));
  AND4_X1   g556(.A1(new_n256_), .A2(new_n594_), .A3(new_n620_), .A4(new_n648_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(new_n651_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n757_), .B1(new_n759_), .B2(new_n756_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT107), .ZN(G1332gat));
  INV_X1    g560(.A(G64gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n758_), .B2(new_n586_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT48), .Z(new_n764_));
  NAND3_X1  g563(.A1(new_n755_), .A2(new_n762_), .A3(new_n586_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1333gat));
  AOI21_X1  g565(.A(new_n365_), .B1(new_n758_), .B2(new_n395_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT49), .Z(new_n768_));
  NAND3_X1  g567(.A1(new_n755_), .A2(new_n365_), .A3(new_n395_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1334gat));
  INV_X1    g569(.A(G78gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n758_), .B2(new_n474_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n474_), .A2(new_n771_), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT109), .Z(new_n776_));
  NAND2_X1  g575(.A1(new_n755_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n774_), .A2(new_n777_), .ZN(G1335gat));
  NAND2_X1  g577(.A1(new_n616_), .A2(new_n619_), .ZN(new_n779_));
  AND4_X1   g578(.A1(new_n329_), .A2(new_n754_), .A3(new_n779_), .A4(new_n648_), .ZN(new_n780_));
  INV_X1    g579(.A(G85gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n651_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n649_), .A2(new_n257_), .A3(new_n620_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT110), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n736_), .A2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(new_n651_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n782_), .B1(new_n787_), .B2(new_n781_), .ZN(G1336gat));
  AOI21_X1  g587(.A(G92gat), .B1(new_n780_), .B2(new_n586_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n586_), .A2(G92gat), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT111), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(new_n786_), .B2(new_n791_), .ZN(G1337gat));
  NAND4_X1  g591(.A1(new_n780_), .A2(new_n395_), .A3(new_n264_), .A4(new_n266_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n736_), .A2(new_n395_), .A3(new_n785_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n794_), .A2(KEYINPUT112), .A3(G99gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT112), .B1(new_n794_), .B2(G99gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n793_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g597(.A1(new_n780_), .A2(new_n265_), .A3(new_n474_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n736_), .A2(new_n474_), .A3(new_n785_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n800_), .A2(new_n801_), .A3(G106gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n800_), .B2(G106gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n799_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g604(.A1(new_n395_), .A2(new_n651_), .A3(new_n592_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n806_), .A2(KEYINPUT119), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(KEYINPUT119), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810_));
  INV_X1    g609(.A(new_n638_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n256_), .A2(new_n811_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n629_), .A2(KEYINPUT116), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n627_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n624_), .A2(new_n626_), .B1(new_n815_), .B2(new_n630_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n814_), .B1(new_n816_), .B2(new_n813_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n631_), .A2(KEYINPUT115), .A3(new_n815_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n640_), .B2(KEYINPUT55), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n635_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n635_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n812_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n241_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n234_), .A2(new_n240_), .A3(new_n247_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n205_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n252_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n641_), .B2(new_n638_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n329_), .B1(new_n824_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n810_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n821_), .A2(new_n635_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n635_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n829_), .B1(new_n838_), .B2(new_n812_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT117), .B(KEYINPUT57), .C1(new_n839_), .C2(new_n329_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n833_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n811_), .A2(new_n828_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n704_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT58), .B(new_n843_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n846_), .A2(KEYINPUT118), .A3(new_n847_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n779_), .B1(new_n842_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n638_), .A2(new_n641_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n644_), .A2(new_n646_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n638_), .A2(new_n641_), .A3(new_n644_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n779_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n704_), .A2(new_n256_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT114), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT54), .B1(new_n859_), .B2(new_n860_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n664_), .A2(KEYINPUT113), .A3(new_n863_), .A4(new_n256_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n861_), .A2(new_n862_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n862_), .B1(new_n864_), .B2(new_n861_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n809_), .B1(new_n853_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G113gat), .B1(new_n868_), .B2(new_n257_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n809_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n844_), .A2(new_n845_), .ZN(new_n871_));
  AND4_X1   g670(.A1(KEYINPUT118), .A2(new_n871_), .A3(new_n718_), .A4(new_n847_), .ZN(new_n872_));
  AOI21_X1  g671(.A(KEYINPUT118), .B1(new_n846_), .B2(new_n847_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n620_), .B1(new_n874_), .B2(new_n841_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n865_), .A2(new_n866_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n870_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n833_), .A2(new_n840_), .B1(new_n847_), .B2(new_n846_), .ZN(new_n878_));
  OAI22_X1  g677(.A1(new_n878_), .A2(new_n620_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n809_), .B2(KEYINPUT120), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(KEYINPUT120), .B2(new_n809_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n877_), .A2(KEYINPUT59), .B1(new_n879_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n257_), .A2(G113gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(KEYINPUT121), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n869_), .B1(new_n883_), .B2(new_n885_), .ZN(G1340gat));
  AOI21_X1  g685(.A(new_n381_), .B1(new_n883_), .B2(new_n648_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n381_), .B1(new_n649_), .B2(KEYINPUT60), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(KEYINPUT60), .B2(new_n381_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n877_), .A2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(KEYINPUT122), .B1(new_n887_), .B2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n882_), .A2(new_n879_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n648_), .B(new_n892_), .C1(new_n868_), .C2(new_n880_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G120gat), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895_));
  INV_X1    g694(.A(new_n890_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n894_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n891_), .A2(new_n897_), .ZN(G1341gat));
  AOI21_X1  g697(.A(G127gat), .B1(new_n868_), .B2(new_n620_), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n899_), .A2(KEYINPUT123), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(KEYINPUT123), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT124), .B(G127gat), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n779_), .A2(new_n902_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n900_), .A2(new_n901_), .B1(new_n883_), .B2(new_n903_), .ZN(G1342gat));
  NAND3_X1  g703(.A1(new_n868_), .A2(new_n377_), .A3(new_n329_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n883_), .A2(new_n718_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n377_), .ZN(G1343gat));
  NAND2_X1  g706(.A1(new_n853_), .A2(new_n867_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n908_), .A2(new_n651_), .A3(new_n715_), .A4(new_n396_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n256_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(new_n398_), .ZN(G1344gat));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n649_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n399_), .ZN(G1345gat));
  NOR2_X1   g712(.A1(new_n909_), .A2(new_n779_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT61), .B(G155gat), .Z(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1346gat));
  OAI21_X1  g715(.A(G162gat), .B1(new_n909_), .B2(new_n704_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n695_), .A2(G162gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n909_), .B2(new_n918_), .ZN(G1347gat));
  INV_X1    g718(.A(new_n879_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n395_), .A2(new_n591_), .A3(new_n586_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(KEYINPUT125), .Z(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n714_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n920_), .A2(new_n923_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT22), .B(G169gat), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n257_), .A2(new_n925_), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT126), .Z(new_n927_));
  NAND2_X1  g726(.A1(new_n924_), .A2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n924_), .A2(new_n257_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n929_), .A2(new_n930_), .A3(G169gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n929_), .B2(G169gat), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n928_), .B1(new_n931_), .B2(new_n932_), .ZN(G1348gat));
  AOI21_X1  g732(.A(G176gat), .B1(new_n924_), .B2(new_n648_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n474_), .B1(new_n853_), .B2(new_n867_), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n922_), .A2(G176gat), .A3(new_n648_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n934_), .B1(new_n935_), .B2(new_n936_), .ZN(G1349gat));
  NAND3_X1  g736(.A1(new_n935_), .A2(new_n620_), .A3(new_n922_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n779_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n939_));
  AOI22_X1  g738(.A1(new_n938_), .A2(new_n333_), .B1(new_n924_), .B2(new_n939_), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n924_), .A2(new_n485_), .A3(new_n329_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n920_), .A2(new_n704_), .A3(new_n923_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n334_), .B2(new_n942_), .ZN(G1351gat));
  NOR4_X1   g742(.A1(new_n395_), .A2(new_n651_), .A3(new_n714_), .A4(new_n587_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n908_), .A2(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n256_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(new_n425_), .ZN(G1352gat));
  NOR2_X1   g746(.A1(new_n945_), .A2(new_n649_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(new_n420_), .ZN(G1353gat));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n950_));
  INV_X1    g749(.A(G211gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n620_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(KEYINPUT127), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n908_), .A2(new_n944_), .A3(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n950_), .A2(new_n951_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n954_), .B(new_n955_), .ZN(G1354gat));
  OAI21_X1  g755(.A(G218gat), .B1(new_n945_), .B2(new_n704_), .ZN(new_n957_));
  OR2_X1    g756(.A1(new_n695_), .A2(G218gat), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n945_), .B2(new_n958_), .ZN(G1355gat));
endmodule


