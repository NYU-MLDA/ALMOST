//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT26), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT26), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n204_), .B(new_n206_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  OR2_X1    g010(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n212_));
  NAND2_X1  g011(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n211_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n211_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n210_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  INV_X1    g018(.A(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT24), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n222_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n212_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n215_), .A2(new_n216_), .ZN(new_n228_));
  INV_X1    g027(.A(G183gat), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n227_), .A2(new_n228_), .B1(new_n229_), .B2(new_n203_), .ZN(new_n230_));
  AND2_X1   g029(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n221_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(new_n223_), .ZN(new_n234_));
  OAI22_X1  g033(.A1(new_n218_), .A2(new_n226_), .B1(new_n230_), .B2(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(G211gat), .A2(G218gat), .ZN(new_n236_));
  INV_X1    g035(.A(G204gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G197gat), .ZN(new_n238_));
  INV_X1    g037(.A(G197gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G204gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G211gat), .A2(G218gat), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n236_), .A2(new_n238_), .A3(new_n240_), .A4(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n240_), .A3(KEYINPUT85), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n236_), .A2(new_n241_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n242_), .A2(KEYINPUT21), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n243_), .A2(KEYINPUT21), .A3(new_n244_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n235_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n243_), .A2(KEYINPUT21), .A3(new_n244_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  INV_X1    g049(.A(new_n241_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(G211gat), .A2(G218gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G197gat), .B(G204gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n250_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n254_), .A2(KEYINPUT85), .B1(new_n236_), .B2(new_n241_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n249_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n229_), .A2(new_n203_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n233_), .A2(new_n223_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT25), .B(G183gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT79), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n206_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n205_), .A2(KEYINPUT79), .A3(G190gat), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n262_), .A2(new_n264_), .A3(new_n204_), .A4(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n226_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n227_), .A2(new_n228_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n257_), .A2(new_n261_), .A3(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n248_), .A2(KEYINPUT20), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G226gat), .A2(G233gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n272_), .B(KEYINPUT19), .Z(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n209_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n276_), .A2(new_n207_), .B1(new_n206_), .B2(new_n263_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n265_), .A2(new_n204_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n226_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n279_), .A2(new_n268_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT90), .B1(new_n280_), .B2(new_n257_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n261_), .A2(new_n269_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT90), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(new_n247_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n286_));
  OAI211_X1 g085(.A(KEYINPUT98), .B(new_n286_), .C1(new_n235_), .C2(new_n247_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n286_), .B1(new_n235_), .B2(new_n247_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT98), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n285_), .A2(new_n287_), .A3(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n275_), .B1(new_n291_), .B2(new_n274_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G8gat), .B(G36gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT100), .B1(new_n292_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n273_), .A2(KEYINPUT20), .ZN(new_n299_));
  INV_X1    g098(.A(new_n218_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n268_), .A2(new_n258_), .ZN(new_n301_));
  AOI22_X1  g100(.A1(new_n300_), .A2(new_n267_), .B1(new_n301_), .B2(new_n260_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n299_), .B1(new_n302_), .B2(new_n257_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n280_), .A2(KEYINPUT90), .A3(new_n257_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n283_), .B1(new_n282_), .B2(new_n247_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT91), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n303_), .B(KEYINPUT91), .C1(new_n304_), .C2(new_n305_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n271_), .A2(new_n274_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT89), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n271_), .A2(KEYINPUT89), .A3(new_n274_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n315_), .A3(new_n297_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT100), .ZN(new_n317_));
  INV_X1    g116(.A(new_n297_), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n281_), .A2(new_n284_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n273_), .B1(new_n319_), .B2(new_n287_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n317_), .B(new_n318_), .C1(new_n320_), .C2(new_n275_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n298_), .A2(new_n316_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT27), .ZN(new_n323_));
  INV_X1    g122(.A(new_n309_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT91), .B1(new_n285_), .B2(new_n303_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n314_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT89), .B1(new_n271_), .B2(new_n274_), .ZN(new_n327_));
  OAI22_X1  g126(.A1(new_n324_), .A2(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n318_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT27), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n330_), .A3(new_n316_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n323_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G113gat), .A2(G120gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G113gat), .A2(G120gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G127gat), .A2(G134gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G127gat), .A2(G134gat), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n335_), .B(new_n336_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G127gat), .ZN(new_n341_));
  INV_X1    g140(.A(G134gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n336_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n343_), .B(new_n337_), .C1(new_n344_), .C2(new_n334_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n333_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348_));
  INV_X1    g147(.A(G141gat), .ZN(new_n349_));
  INV_X1    g148(.A(G148gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT2), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n351_), .A2(new_n354_), .A3(new_n355_), .A4(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(KEYINPUT1), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT1), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(G155gat), .A3(G162gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n363_), .A3(new_n358_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G141gat), .B(G148gat), .Z(new_n365_));
  AOI22_X1  g164(.A1(new_n357_), .A2(new_n360_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n340_), .A2(new_n333_), .A3(new_n345_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n347_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n357_), .A2(new_n360_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n365_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n340_), .A2(new_n333_), .A3(new_n345_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(new_n346_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n368_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n371_), .B(new_n376_), .C1(new_n372_), .C2(new_n346_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT94), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n368_), .A2(new_n373_), .A3(KEYINPUT4), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n374_), .B(KEYINPUT93), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n375_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G57gat), .B(G85gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT99), .ZN(new_n389_));
  INV_X1    g188(.A(new_n387_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n375_), .B(new_n390_), .C1(new_n378_), .C2(new_n381_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n382_), .A2(KEYINPUT99), .A3(new_n387_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n372_), .A2(new_n346_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(KEYINPUT30), .B(G15gat), .Z(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n396_), .A2(new_n398_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT31), .B(G43gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n402_), .B(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n282_), .B(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G71gat), .B(G99gat), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n407_), .B(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n405_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n405_), .A2(new_n410_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n395_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(G50gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n371_), .A2(KEYINPUT29), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT28), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n416_), .A2(new_n417_), .ZN(new_n420_));
  OAI21_X1  g219(.A(G22gat), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n420_), .ZN(new_n422_));
  INV_X1    g221(.A(G22gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n418_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n415_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n421_), .A2(new_n424_), .A3(new_n415_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n371_), .A2(KEYINPUT29), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT84), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G233gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n430_), .A2(G233gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(G228gat), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n429_), .A2(new_n247_), .A3(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G78gat), .B(G106gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT87), .ZN(new_n437_));
  INV_X1    g236(.A(new_n434_), .ZN(new_n438_));
  XOR2_X1   g237(.A(KEYINPUT86), .B(KEYINPUT29), .Z(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n437_), .B(new_n438_), .C1(new_n440_), .C2(new_n257_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n242_), .A2(KEYINPUT21), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n243_), .A2(new_n244_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n445_), .B(new_n249_), .C1(new_n366_), .C2(new_n439_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n437_), .B1(new_n446_), .B2(new_n438_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n435_), .B(new_n436_), .C1(new_n442_), .C2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT83), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n438_), .B1(new_n440_), .B2(new_n257_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT87), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n441_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n436_), .B1(new_n453_), .B2(new_n435_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n450_), .A2(new_n454_), .A3(KEYINPUT88), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT88), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n429_), .A2(new_n247_), .A3(new_n434_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n452_), .B2(new_n441_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT83), .B1(new_n458_), .B2(new_n436_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n435_), .B1(new_n442_), .B2(new_n447_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n436_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n456_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n428_), .B1(new_n455_), .B2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT88), .B1(new_n450_), .B2(new_n454_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n459_), .A2(new_n456_), .A3(new_n462_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n426_), .A4(new_n427_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n332_), .A2(new_n414_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n464_), .A2(new_n394_), .A3(new_n467_), .ZN(new_n471_));
  OAI211_X1 g270(.A(KEYINPUT32), .B(new_n297_), .C1(new_n320_), .C2(new_n275_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n297_), .A2(KEYINPUT32), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n310_), .A2(new_n315_), .A3(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n392_), .A2(new_n472_), .A3(new_n474_), .A4(new_n393_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n391_), .A2(KEYINPUT96), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT33), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n391_), .A2(KEYINPUT96), .A3(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n368_), .A2(new_n373_), .A3(new_n380_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n379_), .A2(new_n374_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n387_), .B(new_n480_), .C1(new_n378_), .C2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n477_), .A2(new_n479_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n329_), .A2(new_n316_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n475_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n332_), .A2(new_n471_), .B1(new_n485_), .B2(new_n468_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n413_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT101), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT101), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n464_), .A2(new_n394_), .A3(new_n467_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n331_), .B2(new_n323_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n479_), .A2(new_n482_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n492_), .A2(new_n316_), .A3(new_n329_), .A4(new_n477_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n493_), .A2(new_n475_), .B1(new_n467_), .B2(new_n464_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n489_), .B(new_n413_), .C1(new_n491_), .C2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n470_), .B1(new_n488_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G71gat), .B(G78gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(KEYINPUT11), .B2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n499_), .B1(KEYINPUT11), .B2(new_n498_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n497_), .A3(KEYINPUT11), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G231gat), .A2(G233gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n502_), .B(new_n503_), .Z(new_n504_));
  XNOR2_X1  g303(.A(G1gat), .B(G8gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT73), .ZN(new_n506_));
  INV_X1    g305(.A(G15gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n423_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G15gat), .A2(G22gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G1gat), .A2(G8gat), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n508_), .A2(new_n509_), .B1(KEYINPUT14), .B2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n506_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n504_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G127gat), .B(G155gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(G211gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT16), .B(G183gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n517_), .A2(KEYINPUT17), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n513_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n517_), .B(KEYINPUT17), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n513_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G232gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT34), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n525_), .A2(KEYINPUT35), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G43gat), .B(G50gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT69), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G29gat), .B(G36gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT15), .ZN(new_n531_));
  XOR2_X1   g330(.A(G85gat), .B(G92gat), .Z(new_n532_));
  NAND2_X1  g331(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n533_));
  INV_X1    g332(.A(G99gat), .ZN(new_n534_));
  INV_X1    g333(.A(G106gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  OAI211_X1 g335(.A(KEYINPUT64), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n536_), .B(new_n537_), .C1(KEYINPUT64), .C2(KEYINPUT7), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT6), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n532_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  AOI21_X1  g343(.A(new_n541_), .B1(KEYINPUT9), .B2(new_n532_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G85gat), .A2(G92gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT10), .B(G99gat), .ZN(new_n547_));
  OAI221_X1 g346(.A(new_n545_), .B1(KEYINPUT9), .B2(new_n546_), .C1(G106gat), .C2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  AOI211_X1 g348(.A(KEYINPUT72), .B(new_n526_), .C1(new_n531_), .C2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n530_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n552_), .A2(KEYINPUT70), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(KEYINPUT70), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n550_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n525_), .A2(KEYINPUT35), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT71), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n550_), .B(new_n556_), .C1(new_n554_), .C2(new_n553_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n561_), .A2(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n558_), .A2(new_n559_), .A3(new_n566_), .A4(new_n560_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n558_), .A2(new_n560_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n564_), .A2(new_n565_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n568_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n496_), .A2(new_n523_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT12), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT66), .ZN(new_n576_));
  INV_X1    g375(.A(new_n502_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n549_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n549_), .A2(new_n577_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n544_), .A2(new_n502_), .A3(new_n548_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n579_), .B(new_n580_), .C1(KEYINPUT66), .C2(new_n575_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n578_), .B1(new_n581_), .B2(new_n576_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G230gat), .A2(G233gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n579_), .A2(new_n580_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(G230gat), .A3(G233gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n588_));
  XNOR2_X1  g387(.A(G120gat), .B(G148gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G176gat), .B(G204gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n587_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n592_), .B(KEYINPUT68), .Z(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n587_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT13), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT13), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n593_), .A2(new_n599_), .A3(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT77), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n512_), .A2(new_n530_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n512_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n531_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n551_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n605_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n609_), .B1(new_n611_), .B2(new_n608_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G169gat), .B(G197gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT75), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G113gat), .B(G141gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT76), .Z(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n612_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n605_), .A2(new_n610_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(G229gat), .A3(G233gat), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n609_), .A3(new_n616_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n602_), .B1(new_n619_), .B2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n617_), .B1(new_n621_), .B2(new_n609_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(KEYINPUT77), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT78), .B1(new_n623_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n622_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT77), .B1(new_n627_), .B2(new_n624_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT78), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n619_), .A2(new_n602_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n626_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n601_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n601_), .A2(KEYINPUT102), .A3(new_n632_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n574_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n202_), .B1(new_n637_), .B2(new_n395_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT37), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n573_), .A2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n568_), .A2(new_n572_), .A3(KEYINPUT37), .A4(new_n569_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n523_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n643_), .A2(new_n496_), .A3(new_n633_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(new_n202_), .A3(new_n395_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n638_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n648_), .B1(new_n646_), .B2(new_n645_), .ZN(G1324gat));
  INV_X1    g448(.A(G8gat), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n323_), .A2(new_n331_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n637_), .B2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT39), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n644_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n655_), .B(new_n656_), .Z(G1325gat));
  AOI21_X1  g456(.A(new_n507_), .B1(new_n637_), .B2(new_n487_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n659_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n644_), .A2(new_n507_), .A3(new_n487_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(G1326gat));
  INV_X1    g462(.A(new_n468_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n423_), .B1(new_n637_), .B2(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT42), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n644_), .A2(new_n423_), .A3(new_n664_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1327gat));
  INV_X1    g467(.A(new_n573_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(new_n522_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n496_), .A2(new_n633_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G29gat), .B1(new_n672_), .B2(new_n395_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n485_), .A2(new_n468_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n674_), .B1(new_n651_), .B2(new_n490_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n489_), .B1(new_n675_), .B2(new_n413_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n486_), .A2(KEYINPUT101), .A3(new_n487_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n469_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n640_), .A2(new_n641_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n678_), .A2(new_n679_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n496_), .B2(new_n680_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT105), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n687_), .B(KEYINPUT43), .C1(new_n496_), .C2(new_n680_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n678_), .A2(KEYINPUT106), .A3(new_n679_), .A4(new_n681_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n684_), .A2(new_n686_), .A3(new_n688_), .A4(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n635_), .A2(new_n523_), .A3(new_n636_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT104), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n635_), .A2(new_n693_), .A3(new_n523_), .A4(new_n636_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n690_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT44), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  AOI211_X1 g499(.A(KEYINPUT107), .B(new_n700_), .C1(new_n690_), .C2(new_n695_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n699_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n395_), .A2(G29gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n673_), .B1(new_n703_), .B2(new_n704_), .ZN(G1328gat));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT108), .ZN(new_n707_));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n672_), .A2(new_n708_), .A3(new_n651_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT45), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT45), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n651_), .B1(new_n698_), .B2(new_n701_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(G36gat), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n706_), .A2(KEYINPUT108), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(G1329gat));
  OAI21_X1  g515(.A(new_n487_), .B1(new_n698_), .B2(new_n701_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n413_), .A2(G43gat), .ZN(new_n718_));
  AOI22_X1  g517(.A1(new_n717_), .A2(G43gat), .B1(new_n672_), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g519(.A1(new_n468_), .A2(G50gat), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT109), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n672_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n468_), .B1(new_n699_), .B2(new_n702_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(new_n415_), .ZN(G1331gat));
  INV_X1    g524(.A(new_n601_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n626_), .A2(new_n631_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n574_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(G57gat), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n728_), .A2(new_n729_), .A3(new_n394_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n678_), .A2(new_n727_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT110), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n726_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n643_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n395_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n730_), .B1(new_n735_), .B2(new_n729_), .ZN(G1332gat));
  INV_X1    g535(.A(G64gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n734_), .A2(new_n737_), .A3(new_n651_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G64gat), .B1(new_n728_), .B2(new_n332_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT48), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1333gat));
  INV_X1    g540(.A(G71gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n734_), .A2(new_n742_), .A3(new_n487_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G71gat), .B1(new_n728_), .B2(new_n413_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT49), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1334gat));
  INV_X1    g545(.A(G78gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n734_), .A2(new_n747_), .A3(new_n664_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G78gat), .B1(new_n728_), .B2(new_n468_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT50), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1335gat));
  NOR2_X1   g550(.A1(new_n733_), .A2(new_n671_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n395_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n601_), .A2(new_n522_), .A3(new_n632_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n690_), .B2(KEYINPUT111), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n496_), .A2(new_n680_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT106), .B1(new_n757_), .B2(new_n679_), .ZN(new_n758_));
  NOR4_X1   g557(.A1(new_n496_), .A2(new_n680_), .A3(new_n683_), .A4(KEYINPUT43), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n688_), .A4(new_n686_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n756_), .A2(KEYINPUT112), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT112), .B1(new_n756_), .B2(new_n762_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n395_), .A2(G85gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n753_), .B1(new_n765_), .B2(new_n766_), .ZN(G1336gat));
  AOI21_X1  g566(.A(G92gat), .B1(new_n752_), .B2(new_n651_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n651_), .A2(G92gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n765_), .B2(new_n769_), .ZN(G1337gat));
  NOR2_X1   g569(.A1(new_n413_), .A2(new_n547_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT113), .B1(new_n752_), .B2(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n763_), .A2(new_n764_), .A3(new_n413_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(new_n534_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n772_), .B(new_n775_), .C1(new_n773_), .C2(new_n534_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1338gat));
  NOR2_X1   g578(.A1(new_n755_), .A2(new_n468_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n535_), .B1(new_n690_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782_));
  XOR2_X1   g581(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n783_));
  OR3_X1    g582(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n783_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n781_), .A2(KEYINPUT116), .A3(new_n783_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n782_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n784_), .A2(new_n787_), .A3(new_n788_), .A4(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n752_), .A2(new_n535_), .A3(new_n664_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n790_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(new_n794_), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT57), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n605_), .A2(new_n607_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n608_), .B1(new_n797_), .B2(KEYINPUT119), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(KEYINPUT119), .B2(new_n797_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n616_), .B1(new_n620_), .B2(new_n608_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n627_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n597_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT55), .B1(new_n582_), .B2(new_n583_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n584_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n582_), .A2(KEYINPUT55), .A3(new_n583_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n594_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT56), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n593_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n802_), .B1(new_n811_), .B2(new_n632_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n796_), .B1(new_n812_), .B2(new_n573_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n727_), .A2(new_n810_), .A3(new_n809_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT57), .B(new_n669_), .C1(new_n814_), .C2(new_n802_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n811_), .A2(KEYINPUT58), .A3(new_n801_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n806_), .A2(new_n807_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n817_), .A2(new_n593_), .A3(new_n808_), .A4(new_n801_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(new_n820_), .A3(new_n681_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n813_), .A2(new_n815_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n523_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n632_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n642_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n824_), .B2(new_n642_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n664_), .B1(new_n823_), .B2(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n651_), .A2(new_n394_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n487_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT120), .B1(new_n830_), .B2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n828_), .B1(new_n822_), .B2(new_n523_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n836_));
  NOR4_X1   g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n664_), .A4(new_n832_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n632_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(G113gat), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n841_));
  NOR4_X1   g640(.A1(new_n835_), .A2(KEYINPUT59), .A3(new_n664_), .A4(new_n832_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n727_), .A2(new_n839_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n838_), .A2(new_n839_), .B1(new_n843_), .B2(new_n844_), .ZN(G1340gat));
  INV_X1    g644(.A(KEYINPUT60), .ZN(new_n846_));
  AOI21_X1  g645(.A(G120gat), .B1(new_n726_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848_));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI22_X1  g648(.A1(new_n847_), .A2(new_n848_), .B1(KEYINPUT60), .B2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n848_), .B2(new_n847_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n841_), .A2(new_n842_), .A3(new_n601_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n849_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(KEYINPUT122), .B(new_n852_), .C1(new_n853_), .C2(new_n849_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1341gat));
  OAI21_X1  g657(.A(new_n522_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n522_), .A2(G127gat), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT123), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n859_), .A2(new_n341_), .B1(new_n843_), .B2(new_n861_), .ZN(G1342gat));
  OAI21_X1  g661(.A(new_n573_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n680_), .A2(new_n342_), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n863_), .A2(new_n342_), .B1(new_n843_), .B2(new_n864_), .ZN(G1343gat));
  NAND3_X1  g664(.A1(new_n831_), .A2(new_n413_), .A3(new_n664_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n835_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n632_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n726_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT124), .B(G148gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1345gat));
  NAND2_X1  g671(.A1(new_n867_), .A2(new_n522_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  AOI21_X1  g674(.A(G162gat), .B1(new_n867_), .B2(new_n573_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n681_), .A2(G162gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT125), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n867_), .B2(new_n878_), .ZN(G1347gat));
  NAND2_X1  g678(.A1(new_n651_), .A2(new_n414_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n835_), .A2(new_n664_), .A3(new_n880_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n881_), .B(new_n632_), .C1(new_n232_), .C2(new_n231_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  INV_X1    g682(.A(new_n880_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n632_), .A2(new_n884_), .ZN(new_n885_));
  XOR2_X1   g684(.A(new_n885_), .B(KEYINPUT126), .Z(new_n886_));
  NAND2_X1  g685(.A1(new_n830_), .A2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n883_), .B1(new_n887_), .B2(G169gat), .ZN(new_n888_));
  AOI211_X1 g687(.A(KEYINPUT62), .B(new_n220_), .C1(new_n830_), .C2(new_n886_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n882_), .B1(new_n888_), .B2(new_n889_), .ZN(G1348gat));
  NAND2_X1  g689(.A1(new_n881_), .A2(new_n726_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g691(.A1(new_n881_), .A2(new_n522_), .ZN(new_n893_));
  MUX2_X1   g692(.A(new_n262_), .B(G183gat), .S(new_n893_), .Z(G1350gat));
  NAND4_X1  g693(.A1(new_n881_), .A2(new_n573_), .A3(new_n204_), .A4(new_n206_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n881_), .A2(new_n681_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n203_), .ZN(G1351gat));
  NOR3_X1   g696(.A1(new_n332_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n835_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n632_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n726_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g703(.A1(new_n835_), .A2(new_n523_), .A3(new_n899_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n905_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n906_));
  XOR2_X1   g705(.A(KEYINPUT63), .B(G211gat), .Z(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n905_), .B2(new_n907_), .ZN(G1354gat));
  AOI21_X1  g707(.A(G218gat), .B1(new_n900_), .B2(new_n573_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n681_), .A2(G218gat), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT127), .Z(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n900_), .B2(new_n911_), .ZN(G1355gat));
endmodule


