//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G99gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT30), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205_));
  INV_X1    g004(.A(G71gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n204_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT81), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT22), .B(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT81), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n211_), .A2(new_n212_), .A3(new_n221_), .A4(new_n213_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n215_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n211_), .B(new_n213_), .C1(new_n225_), .C2(KEYINPUT24), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n216_), .A2(KEYINPUT24), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(new_n224_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT25), .B(G183gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT26), .B(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT80), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT80), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n229_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n208_), .A2(new_n223_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n207_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n204_), .B(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n223_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT82), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n243_), .A2(KEYINPUT31), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(KEYINPUT31), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G113gat), .B(G120gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n244_), .A2(new_n249_), .A3(new_n245_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT95), .ZN(new_n254_));
  OR2_X1    g053(.A1(G155gat), .A2(G162gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G155gat), .A2(G162gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT84), .ZN(new_n258_));
  NOR2_X1   g057(.A1(G141gat), .A2(G148gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT3), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G141gat), .A2(G148gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT2), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n261_), .A2(new_n264_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT84), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n255_), .A2(new_n268_), .A3(new_n256_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n258_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n256_), .A2(KEYINPUT1), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(G155gat), .A3(G162gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n273_), .A3(new_n255_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n262_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n275_), .A2(new_n259_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n274_), .A2(KEYINPUT83), .A3(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT83), .B1(new_n274_), .B2(new_n276_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n270_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n250_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n249_), .B(new_n270_), .C1(new_n278_), .C2(new_n277_), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n280_), .A2(KEYINPUT4), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(new_n283_), .A3(new_n250_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G225gat), .A2(G233gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n254_), .B1(new_n282_), .B2(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n280_), .A2(new_n281_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n285_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n280_), .A2(KEYINPUT4), .A3(new_n281_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n291_), .A2(KEYINPUT95), .A3(new_n286_), .A4(new_n284_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G1gat), .B(G29gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT97), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G57gat), .B(G85gat), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n295_), .A2(new_n296_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  OR3_X1    g099(.A1(new_n297_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n300_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n293_), .A2(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n301_), .A2(new_n302_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n288_), .A2(new_n305_), .A3(new_n290_), .A4(new_n292_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(KEYINPUT99), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT99), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n293_), .A2(new_n308_), .A3(new_n303_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n253_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G8gat), .B(G36gat), .ZN(new_n312_));
  INV_X1    g111(.A(G92gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT18), .B(G64gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT21), .ZN(new_n318_));
  INV_X1    g117(.A(G204gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n319_), .A2(G197gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT86), .B(G204gat), .ZN(new_n322_));
  INV_X1    g121(.A(G197gat), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n318_), .B(new_n321_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G197gat), .A2(G204gat), .ZN(new_n325_));
  OAI211_X1 g124(.A(KEYINPUT21), .B(new_n325_), .C1(new_n322_), .C2(G197gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(G211gat), .B(G218gat), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n319_), .A2(KEYINPUT86), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G204gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n320_), .B1(new_n333_), .B2(G197gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT21), .B1(new_n334_), .B2(KEYINPUT87), .ZN(new_n335_));
  OAI211_X1 g134(.A(KEYINPUT87), .B(new_n321_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n327_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n329_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n220_), .A2(new_n214_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n227_), .A2(KEYINPUT92), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n225_), .B1(new_n227_), .B2(KEYINPUT92), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n232_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n339_), .B1(new_n342_), .B2(new_n226_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n338_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT87), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n323_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n345_), .B1(new_n346_), .B2(new_n320_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n347_), .A2(KEYINPUT21), .A3(new_n327_), .A4(new_n336_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n236_), .A2(new_n348_), .A3(new_n223_), .A4(new_n329_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(KEYINPUT20), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n351_), .B(KEYINPUT19), .Z(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT91), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n350_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT93), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT20), .B1(new_n338_), .B2(new_n343_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n240_), .A2(new_n338_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT94), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT94), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n240_), .A2(new_n338_), .A3(new_n361_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n358_), .A2(new_n360_), .A3(new_n352_), .A4(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT93), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n350_), .A2(new_n364_), .A3(new_n354_), .ZN(new_n365_));
  AND4_X1   g164(.A1(new_n317_), .A2(new_n356_), .A3(new_n363_), .A4(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT101), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT20), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n338_), .B2(new_n343_), .ZN(new_n369_));
  AOI211_X1 g168(.A(KEYINPUT93), .B(new_n353_), .C1(new_n369_), .C2(new_n349_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n364_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(new_n317_), .A3(new_n363_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT101), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT27), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n358_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n377_));
  OAI22_X1  g176(.A1(new_n377_), .A2(new_n352_), .B1(new_n354_), .B2(new_n350_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n376_), .B1(new_n378_), .B2(new_n316_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n367_), .A2(new_n375_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n317_), .B1(new_n372_), .B2(new_n363_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n376_), .B1(new_n381_), .B2(new_n366_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G78gat), .B(G106gat), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n279_), .A2(KEYINPUT29), .ZN(new_n386_));
  INV_X1    g185(.A(G228gat), .ZN(new_n387_));
  INV_X1    g186(.A(G233gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n386_), .A2(new_n390_), .A3(new_n338_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n390_), .B1(new_n386_), .B2(new_n338_), .ZN(new_n393_));
  OAI211_X1 g192(.A(KEYINPUT89), .B(new_n385_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G22gat), .B(G50gat), .Z(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n279_), .B2(KEYINPUT29), .ZN(new_n396_));
  INV_X1    g195(.A(new_n278_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n274_), .A2(KEYINPUT83), .A3(new_n276_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400_));
  INV_X1    g199(.A(new_n395_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n270_), .A4(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n396_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n396_), .B2(new_n402_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n393_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n385_), .A2(KEYINPUT89), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n391_), .A3(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n394_), .A2(new_n406_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT90), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n394_), .A2(new_n406_), .A3(new_n409_), .A4(KEYINPUT90), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n385_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n407_), .A2(new_n391_), .A3(new_n384_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT88), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n406_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n418_), .B(new_n419_), .C1(new_n417_), .C2(new_n416_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n414_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n383_), .A2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n311_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n378_), .A2(KEYINPUT32), .A3(new_n317_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n317_), .A2(KEYINPUT32), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n372_), .A2(new_n363_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n356_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n316_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n289_), .A2(new_n286_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n303_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT98), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT98), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n303_), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n291_), .A2(new_n285_), .A3(new_n284_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n430_), .A2(new_n373_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n292_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n284_), .A2(new_n286_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT95), .B1(new_n440_), .B2(new_n291_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n442_), .A2(KEYINPUT33), .A3(new_n305_), .A4(new_n290_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT33), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n306_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  OAI22_X1  g245(.A1(new_n310_), .A2(new_n428_), .B1(new_n438_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n422_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT100), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n310_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n422_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n383_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n447_), .A2(KEYINPUT100), .A3(new_n422_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n450_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n253_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n424_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G113gat), .B(G141gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G169gat), .B(G197gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G29gat), .B(G36gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(G43gat), .B(G50gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G43gat), .B(G50gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(G29gat), .B(G36gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT75), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G1gat), .B(G8gat), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G1gat), .ZN(new_n472_));
  INV_X1    g271(.A(G8gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT14), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G15gat), .ZN(new_n475_));
  INV_X1    g274(.A(G22gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(G15gat), .A2(G22gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n474_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT74), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n479_), .A2(KEYINPUT74), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n471_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n482_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(new_n470_), .A3(new_n480_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n469_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT76), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT76), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n469_), .A2(new_n489_), .A3(new_n486_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT15), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n467_), .B(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT78), .B1(new_n494_), .B2(new_n486_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n467_), .B(KEYINPUT15), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT78), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n485_), .A4(new_n483_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n491_), .A2(new_n492_), .A3(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n469_), .A2(new_n486_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n491_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n492_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n500_), .A2(KEYINPUT77), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n469_), .A2(new_n486_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT77), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n492_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n460_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n506_), .A2(new_n492_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT77), .ZN(new_n511_));
  INV_X1    g310(.A(new_n460_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n488_), .A2(new_n490_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n507_), .B1(new_n513_), .B2(new_n492_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n511_), .B(new_n512_), .C1(new_n510_), .C2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT79), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n509_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT79), .B(new_n460_), .C1(new_n504_), .C2(new_n508_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT102), .B1(new_n457_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT102), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n517_), .A2(new_n518_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n381_), .A2(new_n366_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n306_), .B(KEYINPUT33), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n437_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n307_), .A2(new_n425_), .A3(new_n309_), .A4(new_n427_), .ZN(new_n526_));
  AOI211_X1 g325(.A(new_n449_), .B(new_n421_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT100), .B1(new_n447_), .B2(new_n422_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n253_), .B1(new_n529_), .B2(new_n453_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n521_), .B(new_n522_), .C1(new_n530_), .C2(new_n424_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT67), .B(G71gat), .ZN(new_n532_));
  INV_X1    g331(.A(G78gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G57gat), .B(G64gat), .Z(new_n535_));
  INV_X1    g334(.A(KEYINPUT11), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n536_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n534_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n532_), .B(G78gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n537_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(new_n486_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G127gat), .B(G155gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(G211gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(KEYINPUT16), .B(G183gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT17), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n550_), .A2(KEYINPUT17), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n546_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n553_), .B1(new_n551_), .B2(new_n546_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT34), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT10), .B(G99gat), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT65), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(G106gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT6), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(G85gat), .A3(G92gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G85gat), .B(G92gat), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n564_), .B(new_n566_), .C1(new_n565_), .C2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n562_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT68), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n568_), .B1(new_n561_), .B2(new_n560_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT68), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n576_));
  OR3_X1    g375(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n564_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n567_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT8), .B1(new_n579_), .B2(KEYINPUT66), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n578_), .B(new_n579_), .C1(KEYINPUT66), .C2(KEYINPUT8), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n494_), .B1(new_n575_), .B2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n467_), .A3(new_n570_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n556_), .B(new_n557_), .C1(new_n586_), .C2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n573_), .B(new_n571_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n496_), .B1(new_n590_), .B2(new_n584_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n556_), .A2(new_n557_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n556_), .A2(new_n557_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n591_), .A2(new_n587_), .A3(new_n592_), .A4(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(G190gat), .B(G218gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT72), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n589_), .A2(new_n594_), .A3(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n601_), .A2(KEYINPUT73), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(KEYINPUT73), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n589_), .A2(new_n594_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n597_), .B(KEYINPUT36), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT37), .ZN(new_n609_));
  INV_X1    g408(.A(new_n607_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT37), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n554_), .B1(new_n609_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT70), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n543_), .A2(KEYINPUT12), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n590_), .B2(new_n584_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT64), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n570_), .A2(new_n583_), .A3(new_n582_), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT12), .B1(new_n621_), .B2(new_n543_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(new_n543_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n617_), .A2(new_n620_), .A3(new_n623_), .A4(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n621_), .A2(new_n543_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n619_), .ZN(new_n629_));
  XOR2_X1   g428(.A(G176gat), .B(G204gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n626_), .A2(new_n629_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n626_), .B2(new_n629_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n615_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n626_), .A2(new_n629_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n634_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n626_), .A2(new_n629_), .A3(new_n635_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(KEYINPUT70), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n638_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT13), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n520_), .A2(new_n531_), .A3(new_n614_), .A4(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n645_), .A2(G1gat), .A3(new_n310_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(KEYINPUT38), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n647_), .A2(KEYINPUT103), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n457_), .A2(new_n611_), .A3(new_n554_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n638_), .A2(new_n642_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT13), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n519_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n649_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n472_), .B1(new_n653_), .B2(new_n451_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n646_), .B2(KEYINPUT38), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n647_), .A2(KEYINPUT103), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n648_), .A2(new_n655_), .A3(new_n656_), .ZN(G1324gat));
  INV_X1    g456(.A(new_n383_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n473_), .B1(new_n653_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n645_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n473_), .A3(new_n658_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(KEYINPUT40), .A3(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1325gat));
  AOI21_X1  g467(.A(new_n475_), .B1(new_n653_), .B2(new_n253_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT41), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n253_), .A2(new_n475_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n645_), .B2(new_n671_), .ZN(G1326gat));
  AOI21_X1  g471(.A(new_n476_), .B1(new_n653_), .B2(new_n421_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT42), .Z(new_n674_));
  NAND2_X1  g473(.A1(new_n421_), .A2(new_n476_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n645_), .B2(new_n675_), .ZN(G1327gat));
  NOR2_X1   g475(.A1(new_n611_), .A2(new_n612_), .ZN(new_n677_));
  AOI211_X1 g476(.A(KEYINPUT37), .B(new_n610_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT43), .B1(new_n457_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n682_), .B(new_n679_), .C1(new_n530_), .C2(new_n424_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n652_), .A2(new_n554_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n685_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT44), .ZN(new_n691_));
  AND4_X1   g490(.A1(G29gat), .A2(new_n689_), .A3(new_n451_), .A4(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n520_), .A2(new_n531_), .A3(new_n611_), .A4(new_n644_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n554_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n451_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n692_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT104), .ZN(G1328gat));
  XNOR2_X1  g497(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n383_), .A2(G36gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n695_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n701_), .ZN(new_n703_));
  NOR4_X1   g502(.A1(new_n693_), .A2(new_n694_), .A3(new_n699_), .A4(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n689_), .A2(new_n658_), .A3(new_n691_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(G36gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n658_), .B1(new_n690_), .B2(KEYINPUT44), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n688_), .B(new_n685_), .C1(new_n681_), .C2(new_n683_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n706_), .B(G36gat), .C1(new_n709_), .C2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n705_), .B1(new_n708_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(KEYINPUT46), .B(new_n705_), .C1(new_n708_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  NAND4_X1  g516(.A1(new_n689_), .A2(G43gat), .A3(new_n253_), .A4(new_n691_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n695_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n719_), .A2(new_n456_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n718_), .B1(new_n720_), .B2(G43gat), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g521(.A(G50gat), .B1(new_n695_), .B2(new_n421_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n689_), .A2(G50gat), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n710_), .A2(new_n422_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n723_), .B1(new_n724_), .B2(new_n725_), .ZN(G1331gat));
  NAND2_X1  g525(.A1(new_n651_), .A2(new_n519_), .ZN(new_n727_));
  NOR4_X1   g526(.A1(new_n457_), .A2(new_n727_), .A3(new_n679_), .A4(new_n554_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G57gat), .B1(new_n728_), .B2(new_n451_), .ZN(new_n729_));
  NOR4_X1   g528(.A1(new_n457_), .A2(new_n727_), .A3(new_n611_), .A4(new_n554_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n730_), .A2(KEYINPUT107), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(KEYINPUT107), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n451_), .A2(G57gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n729_), .B1(new_n733_), .B2(new_n734_), .ZN(G1332gat));
  NAND3_X1  g534(.A1(new_n731_), .A2(new_n658_), .A3(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G64gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT108), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(new_n739_), .A3(G64gat), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n738_), .A2(KEYINPUT48), .A3(new_n740_), .ZN(new_n744_));
  INV_X1    g543(.A(G64gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n728_), .A2(new_n745_), .A3(new_n658_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n743_), .A2(new_n744_), .A3(new_n746_), .ZN(G1333gat));
  NAND3_X1  g546(.A1(new_n728_), .A2(new_n206_), .A3(new_n253_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n733_), .A2(new_n253_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G71gat), .ZN(new_n751_));
  AOI211_X1 g550(.A(KEYINPUT49), .B(new_n206_), .C1(new_n733_), .C2(new_n253_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1334gat));
  NAND3_X1  g552(.A1(new_n728_), .A2(new_n533_), .A3(new_n421_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n733_), .A2(new_n421_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G78gat), .ZN(new_n757_));
  AOI211_X1 g556(.A(KEYINPUT50), .B(new_n533_), .C1(new_n733_), .C2(new_n421_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n727_), .A2(new_n694_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n611_), .C1(new_n530_), .C2(new_n424_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT109), .ZN(new_n762_));
  AOI21_X1  g561(.A(G85gat), .B1(new_n762_), .B2(new_n451_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT110), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n684_), .A2(new_n760_), .ZN(new_n765_));
  INV_X1    g564(.A(G85gat), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n310_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n764_), .A2(new_n767_), .ZN(G1336gat));
  NOR3_X1   g567(.A1(new_n765_), .A2(new_n313_), .A3(new_n383_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n762_), .A2(new_n658_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(new_n313_), .ZN(G1337gat));
  NAND3_X1  g570(.A1(new_n762_), .A2(new_n560_), .A3(new_n253_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n684_), .A2(new_n253_), .A3(new_n760_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(G99gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(G99gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n778_), .A2(KEYINPUT112), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n777_), .B(new_n779_), .ZN(G1338gat));
  NAND3_X1  g579(.A1(new_n762_), .A2(new_n561_), .A3(new_n421_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n684_), .A2(new_n421_), .A3(new_n760_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n782_), .A2(new_n783_), .A3(G106gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n782_), .B2(G106gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g586(.A(G113gat), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n543_), .A2(KEYINPUT12), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n575_), .B2(new_n585_), .ZN(new_n791_));
  NOR4_X1   g590(.A1(new_n791_), .A2(new_n622_), .A3(new_n619_), .A4(new_n624_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT55), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n792_), .B2(KEYINPUT115), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n617_), .A2(new_n625_), .A3(new_n623_), .ZN(new_n796_));
  AOI22_X1  g595(.A1(new_n794_), .A2(new_n795_), .B1(new_n619_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT116), .B1(new_n626_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT55), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n635_), .B1(new_n797_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n789_), .B1(new_n801_), .B2(KEYINPUT56), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n796_), .A2(new_n619_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n626_), .B2(KEYINPUT116), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n800_), .B(new_n803_), .C1(new_n805_), .C2(new_n799_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(KEYINPUT56), .A3(new_n634_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n805_), .B2(new_n799_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n799_), .A2(KEYINPUT55), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n634_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(KEYINPUT119), .A3(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n802_), .A2(new_n807_), .A3(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n460_), .B1(new_n506_), .B2(new_n503_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n513_), .A2(new_n503_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT117), .B(new_n460_), .C1(new_n506_), .C2(new_n503_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n816_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n515_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT118), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n515_), .A2(new_n819_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n636_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n813_), .A2(KEYINPUT58), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT58), .B1(new_n813_), .B2(new_n824_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n680_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n650_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n810_), .A2(new_n811_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n636_), .B1(new_n830_), .B2(new_n807_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n831_), .B2(new_n522_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n828_), .B1(new_n832_), .B2(new_n611_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n810_), .A2(new_n811_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT56), .B1(new_n806_), .B2(new_n634_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n522_), .B(new_n641_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n829_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(KEYINPUT57), .A3(new_n608_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n833_), .A2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n554_), .B1(new_n827_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n694_), .B(new_n519_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n651_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n614_), .A2(KEYINPUT54), .A3(new_n644_), .A4(new_n519_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT113), .B(KEYINPUT114), .Z(new_n846_));
  AND3_X1   g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n421_), .B1(new_n841_), .B2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n658_), .A2(new_n310_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n253_), .A3(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n788_), .B1(new_n852_), .B2(new_n519_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(KEYINPUT120), .B(new_n788_), .C1(new_n852_), .C2(new_n519_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n838_), .B2(new_n608_), .ZN(new_n857_));
  AOI211_X1 g656(.A(new_n828_), .B(new_n611_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n826_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n813_), .A2(KEYINPUT58), .A3(new_n824_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n679_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n694_), .B1(new_n859_), .B2(new_n862_), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n847_), .A2(new_n848_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n422_), .B(new_n851_), .C1(new_n863_), .C2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT59), .B1(new_n865_), .B2(new_n456_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n850_), .A2(new_n867_), .A3(new_n253_), .A4(new_n851_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n522_), .A2(G113gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT121), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n855_), .A2(new_n856_), .B1(new_n869_), .B2(new_n871_), .ZN(G1340gat));
  NAND3_X1  g671(.A1(new_n866_), .A2(new_n651_), .A3(new_n868_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G120gat), .ZN(new_n874_));
  INV_X1    g673(.A(G120gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n644_), .B2(KEYINPUT60), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n850_), .A2(new_n253_), .A3(new_n851_), .A4(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n875_), .A2(KEYINPUT60), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(KEYINPUT122), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n877_), .A2(new_n881_), .A3(new_n878_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n874_), .B1(new_n880_), .B2(new_n882_), .ZN(G1341gat));
  INV_X1    g682(.A(G127gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n554_), .A2(new_n884_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n852_), .A2(new_n554_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n869_), .A2(new_n885_), .B1(new_n886_), .B2(new_n884_), .ZN(G1342gat));
  NAND4_X1  g686(.A1(new_n866_), .A2(G134gat), .A3(new_n679_), .A4(new_n868_), .ZN(new_n888_));
  INV_X1    g687(.A(G134gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n852_), .B2(new_n608_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1343gat));
  AOI21_X1  g690(.A(new_n253_), .B1(new_n841_), .B2(new_n849_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n892_), .A2(new_n421_), .A3(new_n851_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n522_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n651_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g696(.A1(new_n892_), .A2(new_n694_), .A3(new_n421_), .A4(new_n851_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT123), .ZN(new_n899_));
  AOI211_X1 g698(.A(new_n253_), .B(new_n422_), .C1(new_n841_), .C2(new_n849_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n900_), .A2(new_n901_), .A3(new_n694_), .A4(new_n851_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT61), .B(G155gat), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n899_), .A2(new_n902_), .A3(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n899_), .B2(new_n902_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1346gat));
  AOI21_X1  g705(.A(G162gat), .B1(new_n893_), .B2(new_n611_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n893_), .A2(G162gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n679_), .B2(new_n908_), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n311_), .A2(new_n383_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n850_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n912_), .A2(new_n522_), .A3(new_n218_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n522_), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(KEYINPUT124), .Z(new_n915_));
  NAND2_X1  g714(.A1(new_n850_), .A2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G169gat), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n917_), .A2(KEYINPUT62), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(KEYINPUT62), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n913_), .B1(new_n918_), .B2(new_n919_), .ZN(G1348gat));
  NOR2_X1   g719(.A1(new_n911_), .A2(new_n644_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT125), .B(G176gat), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1349gat));
  NOR2_X1   g722(.A1(new_n911_), .A2(new_n554_), .ZN(new_n924_));
  MUX2_X1   g723(.A(G183gat), .B(new_n230_), .S(new_n924_), .Z(G1350gat));
  NAND3_X1  g724(.A1(new_n912_), .A2(new_n611_), .A3(new_n231_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n850_), .A2(new_n679_), .A3(new_n910_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n927_), .A2(new_n928_), .A3(G190gat), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n928_), .B1(new_n927_), .B2(G190gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n926_), .B1(new_n930_), .B2(new_n931_), .ZN(G1351gat));
  NAND3_X1  g731(.A1(new_n892_), .A2(new_n452_), .A3(new_n658_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n519_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(new_n323_), .ZN(G1352gat));
  INV_X1    g734(.A(new_n933_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n651_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(G204gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n938_), .B1(new_n322_), .B2(new_n937_), .ZN(G1353gat));
  XOR2_X1   g738(.A(KEYINPUT63), .B(G211gat), .Z(new_n940_));
  NAND3_X1  g739(.A1(new_n936_), .A2(new_n694_), .A3(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n942_), .B1(new_n933_), .B2(new_n554_), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1354gat));
  NAND4_X1  g743(.A1(new_n892_), .A2(new_n611_), .A3(new_n452_), .A4(new_n658_), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n452_), .ZN(new_n948_));
  AOI211_X1 g747(.A(new_n253_), .B(new_n948_), .C1(new_n841_), .C2(new_n849_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n949_), .A2(KEYINPUT127), .A3(new_n611_), .A4(new_n658_), .ZN(new_n950_));
  INV_X1    g749(.A(G218gat), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n947_), .A2(new_n950_), .A3(new_n951_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n936_), .A2(G218gat), .A3(new_n679_), .ZN(new_n953_));
  AND2_X1   g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1355gat));
endmodule


