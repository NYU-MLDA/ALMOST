//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n891_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT6), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT67), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n202_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(KEYINPUT68), .A2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(G99gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT7), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(new_n212_), .A3(new_n209_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n202_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n205_), .A2(KEYINPUT67), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n203_), .A2(KEYINPUT6), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n207_), .A2(new_n211_), .A3(new_n213_), .A4(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT69), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT8), .ZN(new_n221_));
  XOR2_X1   g020(.A(G85gat), .B(G92gat), .Z(new_n222_));
  NOR4_X1   g021(.A1(KEYINPUT68), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n212_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n225_), .A2(KEYINPUT69), .A3(new_n217_), .A4(new_n207_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .A4(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(KEYINPUT70), .A2(KEYINPUT6), .ZN(new_n228_));
  NAND2_X1  g027(.A1(KEYINPUT70), .A2(KEYINPUT6), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n202_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n214_), .A3(new_n229_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n225_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(new_n222_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT8), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n227_), .A2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT10), .B(G99gat), .Z(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT66), .B(G106gat), .Z(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT9), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(G85gat), .A3(G92gat), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n239_), .A2(new_n217_), .A3(new_n207_), .A4(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n222_), .A2(KEYINPUT9), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n236_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G57gat), .B(G64gat), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n248_), .A2(KEYINPUT11), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(KEYINPUT11), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G71gat), .B(G78gat), .ZN(new_n251_));
  OR3_X1    g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n248_), .A2(new_n251_), .A3(KEYINPUT11), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n247_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT12), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n245_), .B1(new_n227_), .B2(new_n235_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(new_n254_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G230gat), .A2(G233gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n261_), .B(KEYINPUT64), .Z(new_n262_));
  XOR2_X1   g061(.A(new_n262_), .B(KEYINPUT65), .Z(new_n263_));
  AND3_X1   g062(.A1(new_n239_), .A2(new_n217_), .A3(new_n207_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n264_), .A2(KEYINPUT71), .A3(new_n243_), .A4(new_n241_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n236_), .A2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n254_), .A2(new_n257_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n258_), .A2(new_n260_), .A3(new_n263_), .A4(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n256_), .A2(new_n260_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n263_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G120gat), .B(G148gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G176gat), .B(G204gat), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n278_), .B(new_n279_), .Z(new_n280_));
  NAND3_X1  g079(.A1(new_n272_), .A2(new_n275_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n272_), .A2(KEYINPUT73), .A3(new_n275_), .A4(new_n280_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n280_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT74), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n285_), .A2(new_n290_), .A3(new_n287_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(KEYINPUT13), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT13), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n290_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n294_));
  AOI211_X1 g093(.A(KEYINPUT74), .B(new_n286_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(KEYINPUT78), .B(G1gat), .Z(new_n298_));
  INV_X1    g097(.A(G8gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT14), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT79), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G15gat), .B(G22gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n301_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n305_));
  OAI21_X1  g104(.A(G1gat), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n305_), .ZN(new_n307_));
  INV_X1    g106(.A(G1gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(new_n308_), .A3(new_n303_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n309_), .A3(G8gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(G8gat), .B1(new_n306_), .B2(new_n309_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(G29gat), .A2(G36gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G29gat), .A2(G36gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(G43gat), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G29gat), .ZN(new_n317_));
  INV_X1    g116(.A(G36gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G43gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G29gat), .A2(G36gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n316_), .A2(new_n322_), .A3(G50gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(G50gat), .B1(new_n316_), .B2(new_n322_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT75), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n316_), .A2(new_n322_), .ZN(new_n326_));
  INV_X1    g125(.A(G50gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n316_), .A2(new_n322_), .A3(G50gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n325_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT15), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n325_), .A2(new_n331_), .A3(KEYINPUT15), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT83), .B1(new_n313_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G229gat), .A2(G233gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n312_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n323_), .A2(new_n324_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n310_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT83), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n325_), .A2(new_n331_), .A3(KEYINPUT15), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT15), .B1(new_n325_), .B2(new_n331_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n342_), .B(new_n345_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n337_), .A2(new_n338_), .A3(new_n341_), .A4(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n338_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n340_), .B1(new_n339_), .B2(new_n310_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n340_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n311_), .A2(new_n312_), .A3(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n348_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G113gat), .B(G141gat), .ZN(new_n354_));
  INV_X1    g153(.A(G169gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G197gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n353_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n358_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n347_), .A2(new_n352_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n297_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT18), .B(G64gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(G92gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G8gat), .B(G36gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT32), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(KEYINPUT93), .A2(G204gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(KEYINPUT93), .A2(G204gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(G197gat), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G204gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(G197gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT21), .ZN(new_n379_));
  OR2_X1    g178(.A1(G211gat), .A2(G218gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G211gat), .A2(G218gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT97), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT97), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n380_), .A2(new_n384_), .A3(new_n381_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n379_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT93), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n375_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(KEYINPUT93), .A2(G204gat), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n357_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT94), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n375_), .A2(G197gat), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT94), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n389_), .A2(new_n394_), .A3(new_n357_), .A4(new_n390_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n392_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n396_), .A2(KEYINPUT21), .B1(new_n383_), .B2(new_n385_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n374_), .A2(new_n377_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT96), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n374_), .A2(KEYINPUT96), .A3(new_n377_), .A4(new_n398_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n387_), .B1(new_n397_), .B2(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT99), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(KEYINPUT99), .A3(new_n406_), .ZN(new_n410_));
  AOI21_X1  g209(.A(G176gat), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G169gat), .A2(G176gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G183gat), .A2(G190gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT23), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(G183gat), .A2(G190gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n412_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n411_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT24), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT86), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT85), .B1(G169gat), .B2(G176gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(KEYINPUT85), .A2(G169gat), .A3(G176gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n420_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT85), .ZN(new_n425_));
  INV_X1    g224(.A(G176gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n355_), .A3(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(KEYINPUT86), .A3(new_n421_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n419_), .B1(new_n424_), .B2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n415_), .B1(new_n429_), .B2(new_n412_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT24), .B1(new_n427_), .B2(new_n421_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT25), .B(G183gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT26), .B(G190gat), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n418_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT20), .B1(new_n404_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n396_), .A2(KEYINPUT21), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n437_), .A2(new_n386_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n387_), .ZN(new_n439_));
  AOI21_X1  g238(.A(G176gat), .B1(new_n405_), .B2(new_n406_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n417_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT84), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n432_), .A2(new_n433_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n427_), .A2(KEYINPUT86), .A3(new_n421_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT86), .B1(new_n427_), .B2(new_n421_), .ZN(new_n447_));
  OAI211_X1 g246(.A(KEYINPUT24), .B(new_n412_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n415_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n424_), .A2(new_n419_), .A3(new_n428_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n445_), .A2(new_n448_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  AND4_X1   g250(.A1(new_n438_), .A2(new_n439_), .A3(new_n441_), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G226gat), .A2(G233gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT19), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n436_), .A2(new_n452_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n454_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n404_), .B2(new_n435_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n438_), .A2(new_n439_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n451_), .A2(new_n441_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n456_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n371_), .B1(new_n455_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT102), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT3), .ZN(new_n465_));
  INV_X1    g264(.A(G141gat), .ZN(new_n466_));
  INV_X1    g265(.A(G148gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G141gat), .A2(G148gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT2), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n468_), .A2(new_n471_), .A3(new_n472_), .A4(new_n473_), .ZN(new_n474_));
  OR2_X1    g273(.A1(G155gat), .A2(G162gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G155gat), .A2(G162gat), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT90), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(G155gat), .A2(G162gat), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n481_), .A2(KEYINPUT1), .B1(new_n466_), .B2(new_n467_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT1), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n483_), .A3(new_n476_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n484_), .A3(new_n469_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n474_), .A2(KEYINPUT90), .A3(new_n477_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n480_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G127gat), .B(G134gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G113gat), .B(G120gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT87), .ZN(new_n491_));
  INV_X1    g290(.A(new_n488_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G113gat), .B(G120gat), .Z(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(KEYINPUT88), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n488_), .A2(new_n489_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n498_));
  AND4_X1   g297(.A1(new_n491_), .A2(new_n494_), .A3(new_n496_), .A4(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n487_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n492_), .A2(new_n493_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n490_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n480_), .A2(new_n502_), .A3(new_n485_), .A4(new_n486_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G225gat), .A2(G233gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n504_), .B(KEYINPUT100), .Z(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n500_), .A2(new_n503_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT4), .B1(new_n487_), .B2(new_n499_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n474_), .A2(KEYINPUT90), .A3(new_n477_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT90), .B1(new_n474_), .B2(new_n477_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n482_), .A2(new_n484_), .A3(new_n469_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n491_), .A2(new_n494_), .A3(new_n496_), .A4(new_n498_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n503_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n508_), .B1(new_n514_), .B2(KEYINPUT4), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n505_), .B(KEYINPUT101), .Z(new_n516_));
  OAI21_X1  g315(.A(new_n507_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT0), .B(G57gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(G85gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(G1gat), .B(G29gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n507_), .B(new_n521_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n454_), .B1(new_n436_), .B2(new_n452_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n458_), .A2(new_n456_), .A3(new_n461_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n370_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT102), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n529_), .B(new_n371_), .C1(new_n455_), .C2(new_n462_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n464_), .A2(new_n525_), .A3(new_n528_), .A4(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n515_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n521_), .B1(new_n532_), .B2(new_n506_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n516_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT33), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n533_), .A2(new_n535_), .B1(new_n524_), .B2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n526_), .A2(new_n369_), .A3(new_n527_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n369_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n524_), .A2(new_n536_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n537_), .A2(new_n538_), .A3(new_n540_), .A4(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n531_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G78gat), .B(G106gat), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT92), .B1(new_n438_), .B2(new_n439_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G228gat), .A2(G233gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n544_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n404_), .B1(KEYINPUT29), .B2(new_n487_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n544_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n550_), .B(new_n546_), .C1(new_n404_), .C2(KEYINPUT92), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n548_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n549_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT98), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n548_), .A2(new_n551_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n549_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT98), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n548_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n487_), .A2(KEYINPUT29), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G22gat), .B(G50gat), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n563_), .B(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n554_), .A2(new_n560_), .A3(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n563_), .B(new_n564_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n568_), .A2(new_n558_), .A3(new_n559_), .A4(new_n557_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n543_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT103), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT27), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n526_), .A2(new_n369_), .A3(new_n527_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(new_n539_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n369_), .B(KEYINPUT105), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n455_), .B2(new_n462_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(new_n538_), .A3(KEYINPUT27), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n570_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT104), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n525_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n523_), .A2(KEYINPUT104), .A3(new_n524_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT103), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n543_), .A2(new_n587_), .A3(new_n570_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n572_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G15gat), .B(G43gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT31), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT30), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n460_), .B(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n499_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n460_), .B(KEYINPUT30), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n513_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n592_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G71gat), .B(G99gat), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G227gat), .A2(G233gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n595_), .A2(new_n597_), .A3(new_n592_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n599_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n602_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n603_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n605_), .B1(new_n606_), .B2(new_n598_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT89), .ZN(new_n609_));
  INV_X1    g408(.A(new_n579_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n608_), .A2(new_n570_), .A3(new_n610_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n589_), .A2(new_n609_), .B1(new_n585_), .B2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n365_), .A2(new_n612_), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n269_), .A2(new_n345_), .B1(new_n340_), .B2(new_n259_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT34), .Z(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n614_), .B2(KEYINPUT76), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n236_), .A2(new_n246_), .A3(new_n340_), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n235_), .A2(new_n227_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n622_), .B(KEYINPUT76), .C1(new_n623_), .C2(new_n336_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n619_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n617_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n614_), .A2(KEYINPUT76), .A3(new_n620_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n619_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(KEYINPUT35), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n626_), .A2(KEYINPUT77), .A3(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G190gat), .B(G218gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(G134gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(G162gat), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(KEYINPUT36), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n630_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n629_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n616_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n637_));
  OAI211_X1 g436(.A(KEYINPUT36), .B(new_n633_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n634_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n626_), .A2(KEYINPUT77), .A3(new_n639_), .A4(new_n629_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n635_), .A2(new_n638_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT37), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT37), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n635_), .A2(new_n638_), .A3(new_n643_), .A4(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n254_), .B(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n313_), .B(new_n647_), .Z(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G127gat), .B(G155gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(G183gat), .B(G211gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT17), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n649_), .A2(KEYINPUT81), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT81), .B1(new_n649_), .B2(new_n656_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n654_), .B(KEYINPUT17), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT82), .Z(new_n660_));
  NOR2_X1   g459(.A1(new_n649_), .A2(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n657_), .A2(new_n658_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n645_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n613_), .A2(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n665_), .A2(KEYINPUT106), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(KEYINPUT106), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n584_), .B(KEYINPUT107), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n298_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT38), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n663_), .A2(new_n641_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n613_), .A2(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G1gat), .B1(new_n675_), .B2(new_n585_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n669_), .A2(KEYINPUT38), .A3(new_n298_), .A4(new_n670_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n673_), .A2(new_n676_), .A3(new_n677_), .ZN(G1324gat));
  INV_X1    g477(.A(KEYINPUT39), .ZN(new_n679_));
  INV_X1    g478(.A(new_n675_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n579_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n681_), .B2(G8gat), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT39), .B(new_n299_), .C1(new_n680_), .C2(new_n579_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n579_), .A2(new_n299_), .ZN(new_n684_));
  OAI22_X1  g483(.A1(new_n682_), .A2(new_n683_), .B1(new_n668_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(G1325gat));
  OAI21_X1  g486(.A(G15gat), .B1(new_n675_), .B2(new_n609_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT41), .Z(new_n689_));
  NOR3_X1   g488(.A1(new_n665_), .A2(G15gat), .A3(new_n609_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT108), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1326gat));
  OR3_X1    g491(.A1(new_n665_), .A2(G22gat), .A3(new_n570_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G22gat), .B1(new_n675_), .B2(new_n570_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(KEYINPUT42), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(KEYINPUT42), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n693_), .B1(new_n695_), .B2(new_n696_), .ZN(G1327gat));
  INV_X1    g496(.A(new_n641_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n612_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n364_), .A2(new_n663_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G29gat), .B1(new_n702_), .B2(new_n584_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n642_), .A2(new_n644_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n612_), .A2(KEYINPUT43), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n645_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n642_), .A2(KEYINPUT109), .A3(new_n644_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n710_), .B2(new_n612_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT110), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n642_), .A2(KEYINPUT109), .A3(new_n644_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT109), .B1(new_n642_), .B2(new_n644_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n611_), .A2(new_n585_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n543_), .A2(new_n587_), .A3(new_n570_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n587_), .B1(new_n543_), .B2(new_n570_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n570_), .A2(new_n584_), .A3(new_n579_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n717_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT89), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n608_), .B(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n716_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n715_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(KEYINPUT43), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n706_), .B1(new_n712_), .B2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n704_), .B1(new_n727_), .B2(new_n701_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(new_n317_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n706_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n725_), .B1(new_n724_), .B2(KEYINPUT43), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n733_));
  AOI211_X1 g532(.A(KEYINPUT110), .B(new_n733_), .C1(new_n715_), .C2(new_n723_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n731_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n701_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(KEYINPUT44), .A3(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n737_), .A2(new_n670_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n703_), .B1(new_n730_), .B2(new_n738_), .ZN(G1328gat));
  XNOR2_X1  g538(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n728_), .A2(new_n737_), .A3(new_n579_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G36gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n702_), .A2(new_n318_), .A3(new_n579_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n702_), .A2(KEYINPUT45), .A3(new_n318_), .A4(new_n579_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n740_), .B1(new_n742_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n740_), .ZN(new_n750_));
  AOI211_X1 g549(.A(new_n750_), .B(new_n747_), .C1(new_n741_), .C2(G36gat), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1329gat));
  NAND4_X1  g551(.A1(new_n728_), .A2(new_n737_), .A3(G43gat), .A4(new_n608_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n702_), .A2(new_n722_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n320_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g556(.A(new_n570_), .ZN(new_n758_));
  AOI21_X1  g557(.A(G50gat), .B1(new_n702_), .B2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n729_), .A2(new_n327_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n737_), .A2(new_n758_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n759_), .B1(new_n760_), .B2(new_n761_), .ZN(G1331gat));
  INV_X1    g561(.A(new_n297_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n612_), .A2(new_n763_), .A3(new_n362_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n674_), .ZN(new_n765_));
  INV_X1    g564(.A(G57gat), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n585_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n664_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT112), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n670_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n767_), .B1(new_n770_), .B2(new_n766_), .ZN(G1332gat));
  OAI21_X1  g570(.A(G64gat), .B1(new_n765_), .B2(new_n610_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT48), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n610_), .A2(G64gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n768_), .B2(new_n774_), .ZN(G1333gat));
  OAI21_X1  g574(.A(G71gat), .B1(new_n765_), .B2(new_n609_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT49), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n609_), .A2(G71gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n768_), .B2(new_n778_), .ZN(G1334gat));
  OAI21_X1  g578(.A(G78gat), .B1(new_n765_), .B2(new_n570_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT50), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n570_), .A2(G78gat), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT113), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n781_), .B1(new_n768_), .B2(new_n783_), .ZN(G1335gat));
  NAND3_X1  g583(.A1(new_n297_), .A2(new_n663_), .A3(new_n363_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n700_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G85gat), .B1(new_n786_), .B2(new_n670_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n785_), .B(KEYINPUT114), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n735_), .A2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(new_n585_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n787_), .B1(new_n790_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g590(.A(G92gat), .B1(new_n786_), .B2(new_n579_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n789_), .A2(new_n610_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g593(.A(G99gat), .B1(new_n789_), .B2(new_n609_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n786_), .A2(new_n237_), .A3(new_n608_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n797_), .B(new_n798_), .ZN(G1338gat));
  NAND3_X1  g598(.A1(new_n786_), .A2(new_n238_), .A3(new_n758_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n735_), .A2(new_n758_), .A3(new_n788_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n801_), .A2(new_n802_), .A3(G106gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n801_), .B2(G106gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT53), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n800_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1339gat));
  NAND2_X1  g608(.A1(new_n611_), .A2(new_n670_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n338_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT117), .A3(new_n358_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n350_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n348_), .B1(new_n341_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n813_), .B1(new_n815_), .B2(new_n360_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n337_), .A2(new_n348_), .A3(new_n341_), .A4(new_n346_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n812_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n361_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n271_), .A2(new_n260_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT12), .B1(new_n247_), .B2(new_n255_), .ZN(new_n823_));
  OR4_X1    g622(.A1(KEYINPUT55), .A2(new_n822_), .A3(new_n274_), .A4(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n280_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n274_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(new_n272_), .A3(KEYINPUT55), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n824_), .A2(new_n825_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n824_), .A2(KEYINPUT56), .A3(new_n827_), .A4(new_n825_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n362_), .A3(new_n285_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n821_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n698_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(KEYINPUT57), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n831_), .A2(KEYINPUT119), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n819_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n830_), .A2(KEYINPUT119), .A3(new_n831_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n285_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n840_), .A2(KEYINPUT58), .A3(new_n285_), .A4(new_n841_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n645_), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n837_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n834_), .A2(new_n698_), .A3(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n838_), .A2(new_n846_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n663_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n705_), .A2(new_n662_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n292_), .A2(new_n296_), .A3(new_n363_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n852_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n664_), .A2(new_n763_), .A3(new_n363_), .A4(new_n851_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n810_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858_), .B2(new_n362_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n850_), .A2(new_n857_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n810_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n863_));
  NOR2_X1   g662(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n860_), .A2(new_n861_), .A3(new_n863_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n363_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n859_), .B1(new_n868_), .B2(G113gat), .ZN(G1340gat));
  AOI211_X1 g668(.A(KEYINPUT121), .B(new_n763_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871_));
  INV_X1    g670(.A(new_n865_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n867_), .B1(new_n858_), .B2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n871_), .B1(new_n873_), .B2(new_n297_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G120gat), .B1(new_n870_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n763_), .B2(G120gat), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n858_), .B(new_n877_), .C1(new_n876_), .C2(G120gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n878_), .ZN(G1341gat));
  AOI21_X1  g678(.A(G127gat), .B1(new_n858_), .B2(new_n662_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT122), .ZN(new_n881_));
  XOR2_X1   g680(.A(KEYINPUT123), .B(G127gat), .Z(new_n882_));
  NAND3_X1  g681(.A1(new_n873_), .A2(new_n662_), .A3(new_n882_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n881_), .A2(new_n883_), .ZN(G1342gat));
  AOI21_X1  g683(.A(G134gat), .B1(new_n858_), .B2(new_n641_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n705_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(G134gat), .ZN(G1343gat));
  NAND4_X1  g686(.A1(new_n860_), .A2(new_n609_), .A3(new_n580_), .A4(new_n670_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n363_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(new_n466_), .ZN(G1344gat));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n763_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n467_), .ZN(G1345gat));
  NOR2_X1   g691(.A1(new_n888_), .A2(new_n663_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT61), .B(G155gat), .Z(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1346gat));
  INV_X1    g694(.A(G162gat), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n888_), .A2(new_n896_), .A3(new_n710_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n888_), .B2(new_n698_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n899_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n897_), .B1(new_n900_), .B2(new_n901_), .ZN(G1347gat));
  AOI21_X1  g701(.A(new_n363_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n609_), .A2(new_n758_), .A3(new_n670_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n847_), .B1(new_n834_), .B2(new_n698_), .ZN(new_n905_));
  AOI211_X1 g704(.A(new_n641_), .B(new_n837_), .C1(new_n821_), .C2(new_n833_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n662_), .B1(new_n907_), .B2(new_n846_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n855_), .A2(new_n856_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n579_), .B(new_n904_), .C1(new_n908_), .C2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n610_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n913_));
  AOI21_X1  g712(.A(KEYINPUT125), .B1(new_n913_), .B2(new_n904_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n903_), .B1(new_n912_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n916_));
  INV_X1    g715(.A(new_n910_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n362_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n918_), .B2(G169gat), .ZN(new_n919_));
  AOI211_X1 g718(.A(KEYINPUT62), .B(new_n355_), .C1(new_n917_), .C2(new_n362_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n915_), .B1(new_n919_), .B2(new_n920_), .ZN(G1348gat));
  OAI211_X1 g720(.A(new_n426_), .B(new_n297_), .C1(new_n912_), .C2(new_n914_), .ZN(new_n922_));
  OAI21_X1  g721(.A(G176gat), .B1(new_n910_), .B2(new_n763_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1349gat));
  AOI21_X1  g723(.A(G183gat), .B1(new_n917_), .B2(new_n662_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n910_), .A2(new_n911_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n913_), .A2(KEYINPUT125), .A3(new_n904_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n663_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n432_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n925_), .B1(new_n928_), .B2(new_n929_), .ZN(G1350gat));
  OAI211_X1 g729(.A(new_n641_), .B(new_n433_), .C1(new_n912_), .C2(new_n914_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n645_), .B1(new_n912_), .B2(new_n914_), .ZN(new_n932_));
  AOI21_X1  g731(.A(KEYINPUT126), .B1(new_n932_), .B2(G190gat), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n705_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935_));
  INV_X1    g734(.A(G190gat), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n934_), .A2(new_n935_), .A3(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n931_), .B1(new_n933_), .B2(new_n937_), .ZN(G1351gat));
  NOR3_X1   g737(.A1(new_n722_), .A2(new_n584_), .A3(new_n570_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(KEYINPUT127), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n913_), .A2(new_n941_), .ZN(new_n942_));
  OR2_X1    g741(.A1(new_n940_), .A2(KEYINPUT127), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n363_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(new_n357_), .ZN(G1352gat));
  NAND2_X1  g745(.A1(new_n389_), .A2(new_n390_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n942_), .A2(new_n297_), .A3(new_n943_), .ZN(new_n948_));
  MUX2_X1   g747(.A(new_n947_), .B(G204gat), .S(new_n948_), .Z(G1353gat));
  XNOR2_X1  g748(.A(KEYINPUT63), .B(G211gat), .ZN(new_n950_));
  OR2_X1    g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n942_), .A2(new_n662_), .A3(new_n943_), .ZN(new_n952_));
  MUX2_X1   g751(.A(new_n950_), .B(new_n951_), .S(new_n952_), .Z(G1354gat));
  INV_X1    g752(.A(G218gat), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n944_), .A2(new_n954_), .A3(new_n705_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n942_), .A2(new_n641_), .A3(new_n943_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n955_), .B1(new_n954_), .B2(new_n956_), .ZN(G1355gat));
endmodule


