//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n945_, new_n946_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n961_, new_n962_;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202_));
  INV_X1    g001(.A(G155gat), .ZN(new_n203_));
  INV_X1    g002(.A(G162gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OAI22_X1  g006(.A1(new_n207_), .A2(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT89), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n208_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n215_), .A2(KEYINPUT87), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(KEYINPUT87), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n214_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n215_), .B(KEYINPUT3), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n214_), .B(KEYINPUT2), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n207_), .B1(G155gat), .B2(G162gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT29), .B1(new_n219_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(G204gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(G197gat), .ZN(new_n227_));
  INV_X1    g026(.A(G197gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(G204gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT21), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT91), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n229_), .B1(new_n232_), .B2(new_n227_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT91), .B1(new_n226_), .B2(G197gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n230_), .B(new_n231_), .C1(new_n235_), .C2(KEYINPUT21), .ZN(new_n236_));
  INV_X1    g035(.A(new_n231_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(KEYINPUT21), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n225_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G228gat), .ZN(new_n241_));
  INV_X1    g040(.A(G233gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n225_), .B(new_n239_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G78gat), .B(G106gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n244_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT92), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n244_), .A2(new_n245_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n246_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT93), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(KEYINPUT93), .A3(new_n246_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n248_), .A2(new_n249_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n250_), .A2(new_n254_), .A3(new_n255_), .A4(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n219_), .A2(new_n224_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT28), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT28), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n258_), .A2(new_n262_), .A3(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT90), .ZN(new_n265_));
  XOR2_X1   g064(.A(G22gat), .B(G50gat), .Z(new_n266_));
  INV_X1    g065(.A(KEYINPUT90), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n261_), .A2(new_n267_), .A3(new_n263_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n265_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n266_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n261_), .A2(new_n267_), .A3(new_n263_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n267_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n257_), .A2(new_n269_), .A3(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT25), .B(G183gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G190gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n275_), .A2(new_n276_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT23), .ZN(new_n282_));
  INV_X1    g081(.A(G169gat), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n280_), .B(new_n282_), .C1(KEYINPUT24), .C2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n282_), .B1(G183gat), .B2(G190gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(G169gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n239_), .A2(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n292_), .A2(KEYINPUT94), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G226gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT19), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT20), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n236_), .A2(new_n238_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n291_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n292_), .A2(KEYINPUT94), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n293_), .A2(new_n296_), .A3(new_n300_), .A4(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n292_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n295_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G8gat), .B(G36gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G64gat), .B(G92gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n302_), .A2(new_n304_), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT27), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n293_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n295_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n300_), .A2(new_n296_), .A3(new_n292_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n312_), .B1(new_n309_), .B2(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(KEYINPUT83), .B(KEYINPUT84), .Z(new_n318_));
  NAND2_X1  g117(.A1(G227gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G71gat), .B(G99gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT86), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n322_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n291_), .B(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G15gat), .B(G43gat), .Z(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n291_), .B(KEYINPUT30), .ZN(new_n331_));
  INV_X1    g130(.A(new_n329_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G127gat), .B(G134gat), .Z(new_n334_));
  XOR2_X1   g133(.A(G113gat), .B(G120gat), .Z(new_n335_));
  XOR2_X1   g134(.A(new_n334_), .B(new_n335_), .Z(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n330_), .A2(new_n333_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n337_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n326_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n330_), .A2(new_n333_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n336_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(new_n338_), .A3(new_n325_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(KEYINPUT99), .B(KEYINPUT27), .Z(new_n346_));
  NAND2_X1  g145(.A1(new_n302_), .A2(new_n304_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n309_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n346_), .B1(new_n348_), .B2(new_n311_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n317_), .A2(new_n345_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n273_), .A2(new_n269_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n252_), .A3(new_n248_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n274_), .A2(new_n350_), .A3(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n336_), .B1(new_n219_), .B2(new_n224_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n354_), .A2(KEYINPUT4), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT96), .ZN(new_n360_));
  OAI221_X1 g159(.A(new_n337_), .B1(new_n222_), .B2(new_n223_), .C1(new_n213_), .C2(new_n218_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n354_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n360_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n354_), .A2(new_n361_), .A3(KEYINPUT96), .A4(KEYINPUT4), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n359_), .A2(new_n366_), .ZN(new_n367_));
  OAI22_X1  g166(.A1(new_n367_), .A2(KEYINPUT97), .B1(new_n362_), .B2(new_n357_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n358_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT97), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G1gat), .B(G29gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G85gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT0), .B(G57gat), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n373_), .B(new_n374_), .Z(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n368_), .A2(new_n371_), .A3(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n362_), .A2(new_n357_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n367_), .A2(KEYINPUT97), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n375_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n377_), .A2(new_n381_), .A3(KEYINPUT98), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT98), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n376_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n379_), .A2(new_n375_), .A3(new_n380_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n353_), .B1(new_n382_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT100), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT98), .B1(new_n377_), .B2(new_n381_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n384_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(KEYINPUT100), .A3(new_n353_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n317_), .A2(new_n349_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n254_), .A2(new_n255_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n248_), .B(KEYINPUT92), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n351_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n351_), .A2(new_n252_), .A3(new_n248_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n395_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n400_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n274_), .A2(new_n352_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n385_), .A2(new_n403_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n379_), .A2(new_n380_), .A3(KEYINPUT33), .A4(new_n375_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n348_), .A2(new_n311_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n366_), .A2(new_n356_), .A3(new_n355_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n362_), .A2(new_n356_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n408_), .A2(new_n375_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n406_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n404_), .A2(new_n405_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n347_), .B1(KEYINPUT32), .B2(new_n310_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n310_), .A2(KEYINPUT32), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n412_), .B1(new_n413_), .B2(new_n316_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n414_), .B1(new_n377_), .B2(new_n381_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n402_), .B1(new_n411_), .B2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n345_), .B1(new_n401_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n394_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G229gat), .A2(G233gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G15gat), .B(G22gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G1gat), .A2(G8gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT77), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(KEYINPUT14), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n423_), .B2(KEYINPUT14), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT78), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(G1gat), .B(G8gat), .Z(new_n429_));
  INV_X1    g228(.A(new_n427_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT78), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n422_), .A4(new_n425_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n428_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n429_), .B1(new_n428_), .B2(new_n432_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G29gat), .B(G36gat), .Z(new_n435_));
  XOR2_X1   g234(.A(G43gat), .B(G50gat), .Z(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G29gat), .B(G36gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G43gat), .B(G50gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(new_n433_), .A2(new_n434_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n428_), .A2(new_n432_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n429_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n428_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n441_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n421_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n437_), .A2(KEYINPUT15), .A3(new_n440_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT15), .B1(new_n437_), .B2(new_n440_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n453_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n446_), .A2(new_n441_), .A3(new_n447_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n420_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n419_), .B1(new_n450_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G113gat), .B(G141gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G169gat), .B(G197gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n459_), .B(new_n460_), .Z(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n449_), .A2(KEYINPUT81), .A3(new_n456_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n458_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n449_), .A2(new_n456_), .A3(new_n461_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT82), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT82), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n449_), .A2(new_n467_), .A3(new_n456_), .A4(new_n461_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n464_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G176gat), .B(G204gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT68), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G120gat), .B(G148gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT69), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G230gat), .A2(G233gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n480_), .B(KEYINPUT64), .Z(new_n481_));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT6), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(G99gat), .A3(G106gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  OR2_X1    g285(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n487_));
  INV_X1    g286(.A(G106gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(G85gat), .ZN(new_n491_));
  INV_X1    g290(.A(G92gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G85gat), .A2(G92gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(KEYINPUT9), .A3(new_n494_), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n494_), .A2(KEYINPUT9), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n486_), .A2(new_n490_), .A3(new_n495_), .A4(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n494_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n483_), .A2(new_n485_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT7), .ZN(new_n502_));
  INV_X1    g301(.A(G99gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n488_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n500_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT8), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n486_), .A2(new_n505_), .A3(new_n504_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT8), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(new_n510_), .A3(new_n500_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n498_), .B1(new_n508_), .B2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G57gat), .B(G64gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G71gat), .B(G78gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(KEYINPUT11), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(KEYINPUT11), .ZN(new_n516_));
  INV_X1    g315(.A(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n513_), .A2(KEYINPUT11), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n515_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n481_), .B1(new_n512_), .B2(new_n520_), .ZN(new_n521_));
  NOR3_X1   g320(.A1(new_n512_), .A2(KEYINPUT12), .A3(new_n520_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT12), .ZN(new_n523_));
  INV_X1    g322(.A(new_n505_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AOI211_X1 g325(.A(KEYINPUT8), .B(new_n499_), .C1(new_n526_), .C2(new_n486_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n510_), .B1(new_n509_), .B2(new_n500_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n497_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n520_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n523_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n521_), .B1(new_n522_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT66), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT66), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n534_), .B(new_n521_), .C1(new_n522_), .C2(new_n531_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n481_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n529_), .A2(new_n530_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n520_), .B(new_n497_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT65), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n479_), .B1(new_n536_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT70), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n540_), .B(KEYINPUT65), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n545_), .A2(new_n477_), .A3(new_n533_), .A4(new_n535_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n543_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n544_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n549_), .A2(KEYINPUT13), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(KEYINPUT13), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT71), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n550_), .A2(KEYINPUT71), .A3(new_n551_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n471_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n418_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n529_), .A2(new_n453_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT34), .ZN(new_n560_));
  OAI221_X1 g359(.A(new_n558_), .B1(KEYINPUT35), .B2(new_n560_), .C1(new_n442_), .C2(new_n529_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(KEYINPUT35), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT72), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n561_), .B(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G134gat), .B(G162gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(G190gat), .B(G218gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT36), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT74), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n564_), .A2(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT75), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(KEYINPUT37), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(KEYINPUT37), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT76), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n580_), .B1(new_n574_), .B2(new_n577_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n520_), .B(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n433_), .A2(new_n434_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n587_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT79), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G127gat), .B(G155gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT16), .ZN(new_n592_));
  XOR2_X1   g391(.A(G183gat), .B(G211gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n594_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n595_), .B1(KEYINPUT17), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n595_), .A2(KEYINPUT17), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(KEYINPUT80), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT80), .ZN(new_n604_));
  INV_X1    g403(.A(new_n601_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n604_), .B1(new_n599_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n584_), .A2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n557_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(G1gat), .ZN(new_n611_));
  INV_X1    g410(.A(new_n392_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n614_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n574_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n599_), .A2(new_n605_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n557_), .A2(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n620_), .A2(new_n612_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n615_), .B(new_n616_), .C1(new_n611_), .C2(new_n621_), .ZN(G1324gat));
  INV_X1    g421(.A(G8gat), .ZN(new_n623_));
  INV_X1    g422(.A(new_n395_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n610_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT102), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n557_), .A2(new_n626_), .A3(new_n624_), .A4(new_n619_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n627_), .A2(G8gat), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n557_), .A2(new_n624_), .A3(new_n619_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT102), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n628_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n629_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n625_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n625_), .B(new_n635_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1325gat));
  INV_X1    g438(.A(G15gat), .ZN(new_n640_));
  INV_X1    g439(.A(new_n345_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n620_), .B2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT41), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n610_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1326gat));
  INV_X1    g444(.A(G22gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n620_), .B2(new_n402_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT42), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n610_), .A2(new_n646_), .A3(new_n402_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1327gat));
  INV_X1    g449(.A(new_n608_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n574_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n557_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n612_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n582_), .A2(new_n583_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n394_), .B2(new_n417_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n608_), .B1(new_n656_), .B2(KEYINPUT43), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n411_), .A2(new_n415_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n402_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n624_), .B1(new_n274_), .B2(new_n352_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n392_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  AOI22_X1  g462(.A1(new_n663_), .A2(new_n345_), .B1(new_n389_), .B2(new_n393_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(new_n655_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n657_), .A2(new_n666_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n667_), .A2(KEYINPUT104), .A3(KEYINPUT44), .A4(new_n556_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n664_), .B2(new_n655_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n418_), .A2(KEYINPUT43), .A3(new_n584_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n670_), .A2(new_n556_), .A3(new_n671_), .A4(new_n608_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n668_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n673_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n612_), .A2(G29gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n654_), .B1(new_n677_), .B2(new_n678_), .ZN(G1328gat));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(G36gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n395_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n675_), .B2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n395_), .A2(G36gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n557_), .A2(new_n652_), .A3(new_n686_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n687_), .A2(KEYINPUT45), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(KEYINPUT45), .ZN(new_n689_));
  AOI22_X1  g488(.A1(new_n688_), .A2(new_n689_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n682_), .B1(new_n685_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n682_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n676_), .A2(new_n624_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n674_), .B2(new_n668_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n693_), .B(new_n690_), .C1(new_n695_), .C2(new_n683_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n692_), .A2(new_n696_), .ZN(G1329gat));
  NAND4_X1  g496(.A1(new_n675_), .A2(G43gat), .A3(new_n641_), .A4(new_n676_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n653_), .A2(new_n641_), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n699_), .A2(G43gat), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT47), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n698_), .A2(new_n703_), .A3(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1330gat));
  AOI21_X1  g504(.A(G50gat), .B1(new_n653_), .B2(new_n402_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n402_), .A2(G50gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n677_), .B2(new_n707_), .ZN(G1331gat));
  NAND2_X1  g507(.A1(new_n554_), .A2(new_n555_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n709_), .A2(new_n470_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n418_), .A2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n608_), .A2(new_n617_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G57gat), .B1(new_n714_), .B2(new_n392_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n711_), .A2(new_n609_), .ZN(new_n716_));
  INV_X1    g515(.A(G57gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n612_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1332gat));
  INV_X1    g518(.A(G64gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n713_), .B2(new_n624_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT106), .B(KEYINPUT48), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n716_), .A2(new_n720_), .A3(new_n624_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1333gat));
  INV_X1    g524(.A(G71gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n716_), .A2(new_n726_), .A3(new_n641_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT49), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n713_), .A2(new_n641_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G71gat), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT49), .B(new_n726_), .C1(new_n713_), .C2(new_n641_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT107), .ZN(G1334gat));
  INV_X1    g532(.A(G78gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n713_), .B2(new_n402_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT50), .Z(new_n736_));
  NAND3_X1  g535(.A1(new_n716_), .A2(new_n734_), .A3(new_n402_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1335gat));
  NAND2_X1  g537(.A1(new_n667_), .A2(new_n710_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739_), .B2(new_n392_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n711_), .A2(new_n652_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(new_n491_), .A3(new_n612_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1336gat));
  AOI21_X1  g542(.A(G92gat), .B1(new_n741_), .B2(new_n624_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT108), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n739_), .A2(new_n492_), .A3(new_n395_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1337gat));
  OAI21_X1  g546(.A(G99gat), .B1(new_n739_), .B2(new_n345_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n741_), .A2(new_n487_), .A3(new_n489_), .A4(new_n641_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g550(.A1(new_n741_), .A2(new_n488_), .A3(new_n402_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n667_), .A2(new_n402_), .A3(new_n710_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(G106gat), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n754_), .B1(new_n753_), .B2(G106gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n752_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n752_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1339gat));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763_));
  INV_X1    g562(.A(new_n618_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n533_), .A2(new_n767_), .A3(new_n535_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n539_), .B1(new_n522_), .B2(new_n531_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n539_), .A2(new_n537_), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT12), .B1(new_n512_), .B2(new_n520_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n529_), .A2(new_n523_), .A3(new_n530_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n481_), .A2(new_n769_), .B1(new_n773_), .B2(KEYINPUT55), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n768_), .A2(KEYINPUT110), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n479_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT110), .B1(new_n768_), .B2(new_n774_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n766_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n777_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n479_), .A4(new_n775_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n470_), .A2(new_n546_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n454_), .A2(new_n455_), .A3(new_n421_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n420_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(new_n462_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n442_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n421_), .B1(new_n789_), .B2(new_n455_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n790_), .A2(KEYINPUT111), .A3(new_n461_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n784_), .B(new_n785_), .C1(new_n788_), .C2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n469_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n787_), .A2(new_n786_), .A3(new_n462_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT111), .B1(new_n790_), .B2(new_n461_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n784_), .B1(new_n796_), .B2(new_n785_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT113), .B1(new_n793_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n785_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT112), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n469_), .A4(new_n792_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n798_), .A2(new_n802_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n781_), .A2(new_n783_), .B1(new_n549_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n765_), .B1(new_n804_), .B2(new_n617_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n549_), .A2(new_n803_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n782_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n807_));
  OAI211_X1 g606(.A(KEYINPUT57), .B(new_n574_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n805_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n778_), .A2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT114), .B(new_n766_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n780_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n803_), .A2(new_n546_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n813_), .A2(new_n814_), .A3(KEYINPUT58), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n584_), .A3(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n809_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n817_), .A2(KEYINPUT115), .A3(new_n584_), .A4(new_n818_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n764_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n470_), .B1(new_n602_), .B2(new_n606_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n549_), .A2(KEYINPUT13), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n549_), .A2(KEYINPUT13), .ZN(new_n826_));
  OAI211_X1 g625(.A(KEYINPUT109), .B(new_n824_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n827_), .A2(new_n655_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n552_), .A2(new_n824_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT109), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n827_), .A2(new_n655_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT109), .B1(new_n552_), .B2(new_n824_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT54), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n833_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n763_), .B1(new_n823_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n803_), .A2(new_n546_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n776_), .A2(new_n766_), .A3(new_n777_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n810_), .B2(new_n778_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n839_), .B1(new_n841_), .B2(new_n812_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n584_), .B1(new_n842_), .B2(KEYINPUT58), .ZN(new_n843_));
  INV_X1    g642(.A(new_n818_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n820_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n809_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n822_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n618_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n833_), .A2(new_n836_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(KEYINPUT116), .A3(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n612_), .A2(new_n353_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n838_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT117), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n838_), .A2(new_n850_), .A3(new_n854_), .A4(new_n851_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n470_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(G113gat), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n856_), .A2(KEYINPUT118), .A3(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n852_), .A2(KEYINPUT59), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT119), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n852_), .A2(new_n864_), .A3(KEYINPUT59), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n846_), .A2(new_n819_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n608_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n837_), .B1(KEYINPUT120), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(KEYINPUT120), .B2(new_n867_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n851_), .A2(new_n870_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n863_), .A2(new_n865_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n471_), .A2(new_n857_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n860_), .A2(new_n861_), .B1(new_n872_), .B2(new_n873_), .ZN(G1340gat));
  NAND2_X1  g673(.A1(new_n869_), .A2(new_n871_), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n852_), .A2(new_n864_), .A3(KEYINPUT59), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n864_), .B1(new_n852_), .B2(KEYINPUT59), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n875_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(G120gat), .B1(new_n878_), .B2(new_n709_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n709_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT60), .ZN(new_n881_));
  AOI21_X1  g680(.A(G120gat), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n881_), .B2(G120gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n853_), .A2(new_n883_), .A3(new_n855_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n853_), .A2(new_n883_), .A3(KEYINPUT121), .A4(new_n855_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n879_), .A2(new_n888_), .ZN(G1341gat));
  INV_X1    g688(.A(G127gat), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n853_), .A2(new_n890_), .A3(new_n651_), .A4(new_n855_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n764_), .B(new_n875_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n891_), .B1(new_n893_), .B2(new_n890_), .ZN(G1342gat));
  INV_X1    g693(.A(G134gat), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n853_), .A2(new_n895_), .A3(new_n617_), .A4(new_n855_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n584_), .B(new_n875_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n898_), .B2(new_n895_), .ZN(G1343gat));
  AND2_X1   g698(.A1(new_n838_), .A2(new_n850_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n612_), .A2(new_n661_), .A3(new_n345_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT122), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n470_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g705(.A1(new_n903_), .A2(new_n709_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT123), .B(G148gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1345gat));
  NOR2_X1   g708(.A1(new_n903_), .A2(new_n608_), .ZN(new_n910_));
  XOR2_X1   g709(.A(KEYINPUT61), .B(G155gat), .Z(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1346gat));
  OAI21_X1  g711(.A(G162gat), .B1(new_n903_), .B2(new_n655_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n617_), .A2(new_n204_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n903_), .B2(new_n914_), .ZN(G1347gat));
  NOR2_X1   g714(.A1(new_n612_), .A2(new_n395_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n641_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT124), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n402_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n869_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n470_), .ZN(new_n921_));
  OAI211_X1 g720(.A(KEYINPUT62), .B(G169gat), .C1(new_n921_), .C2(KEYINPUT22), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n869_), .A2(new_n919_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n471_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT22), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n923_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n283_), .B1(new_n925_), .B2(new_n923_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n922_), .B1(new_n927_), .B2(new_n928_), .ZN(G1348gat));
  AOI21_X1  g728(.A(G176gat), .B1(new_n920_), .B2(new_n880_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n900_), .A2(new_n659_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n918_), .A2(new_n284_), .A3(new_n709_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n930_), .B1(new_n931_), .B2(new_n932_), .ZN(G1349gat));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n618_), .A2(new_n275_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n920_), .A2(new_n934_), .A3(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n935_), .ZN(new_n937_));
  OAI21_X1  g736(.A(KEYINPUT125), .B1(new_n924_), .B2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(G183gat), .ZN(new_n940_));
  INV_X1    g739(.A(new_n918_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n931_), .A2(new_n651_), .A3(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n939_), .B1(new_n940_), .B2(new_n942_), .ZN(G1350gat));
  OAI21_X1  g742(.A(G190gat), .B1(new_n924_), .B2(new_n655_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n617_), .A2(new_n276_), .ZN(new_n945_));
  XOR2_X1   g744(.A(new_n945_), .B(KEYINPUT126), .Z(new_n946_));
  OAI21_X1  g745(.A(new_n944_), .B1(new_n924_), .B2(new_n946_), .ZN(G1351gat));
  NAND3_X1  g746(.A1(new_n916_), .A2(new_n402_), .A3(new_n345_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n900_), .A2(new_n949_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n950_), .A2(new_n471_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(KEYINPUT127), .B(G197gat), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n951_), .B(new_n952_), .ZN(G1352gat));
  NOR2_X1   g752(.A1(new_n950_), .A2(new_n709_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(new_n226_), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n900_), .A2(new_n764_), .A3(new_n949_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n957_));
  AND2_X1   g756(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n956_), .A2(new_n957_), .A3(new_n958_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n959_), .B1(new_n956_), .B2(new_n957_), .ZN(G1354gat));
  OAI21_X1  g759(.A(G218gat), .B1(new_n950_), .B2(new_n655_), .ZN(new_n961_));
  OR2_X1    g760(.A1(new_n574_), .A2(G218gat), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n961_), .B1(new_n950_), .B2(new_n962_), .ZN(G1355gat));
endmodule


