//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202_));
  INV_X1    g001(.A(G204gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G197gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT90), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G197gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G204gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n204_), .A2(new_n205_), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT21), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n204_), .A2(new_n208_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n211_), .B(new_n212_), .C1(KEYINPUT21), .C2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n212_), .B(KEYINPUT91), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(KEYINPUT21), .A3(new_n213_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT92), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  OR2_X1    g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT2), .ZN(new_n223_));
  INV_X1    g022(.A(G141gat), .ZN(new_n224_));
  INV_X1    g023(.A(G148gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT3), .B1(new_n226_), .B2(KEYINPUT87), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n226_), .A2(KEYINPUT87), .A3(KEYINPUT3), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n220_), .B(new_n221_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n220_), .A2(KEYINPUT1), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n220_), .A2(KEYINPUT1), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n231_), .A2(KEYINPUT86), .A3(new_n232_), .A4(new_n221_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n226_), .A2(new_n222_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n233_), .B(new_n234_), .C1(KEYINPUT86), .C2(new_n231_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT29), .ZN(new_n237_));
  INV_X1    g036(.A(G233gat), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n238_), .A2(KEYINPUT89), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(KEYINPUT89), .ZN(new_n240_));
  OAI21_X1  g039(.A(G228gat), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n202_), .B1(new_n219_), .B2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n217_), .B(KEYINPUT92), .ZN(new_n244_));
  INV_X1    g043(.A(new_n242_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(KEYINPUT93), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n217_), .B(KEYINPUT94), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n237_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n241_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G78gat), .B(G106gat), .Z(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n253_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n247_), .A2(new_n251_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n236_), .A2(KEYINPUT29), .ZN(new_n258_));
  XOR2_X1   g057(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G22gat), .B(G50gat), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n236_), .A2(KEYINPUT29), .A3(new_n259_), .ZN(new_n264_));
  OR3_X1    g063(.A1(new_n261_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT95), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n263_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n266_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n257_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n254_), .A2(new_n269_), .A3(new_n256_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G127gat), .B(G134gat), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n274_), .A2(KEYINPUT85), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(KEYINPUT85), .ZN(new_n276_));
  XOR2_X1   g075(.A(G113gat), .B(G120gat), .Z(new_n277_));
  OR3_X1    g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n277_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n280_), .B(KEYINPUT31), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G71gat), .B(G99gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(G43gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G227gat), .A2(G233gat), .ZN(new_n285_));
  INV_X1    g084(.A(G15gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n284_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT84), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT25), .ZN(new_n290_));
  INV_X1    g089(.A(G183gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT78), .B(G183gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n292_), .B1(new_n293_), .B2(new_n290_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(G190gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(KEYINPUT24), .A3(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n296_), .A2(KEYINPUT79), .A3(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n297_), .A2(KEYINPUT24), .ZN(new_n301_));
  INV_X1    g100(.A(G190gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT23), .B1(new_n291_), .B2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT80), .ZN(new_n304_));
  OR3_X1    g103(.A1(new_n291_), .A2(new_n302_), .A3(KEYINPUT23), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n300_), .A2(new_n301_), .A3(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(KEYINPUT79), .B1(new_n296_), .B2(new_n299_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT22), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(G169gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(G176gat), .B1(new_n311_), .B2(KEYINPUT82), .ZN(new_n312_));
  XOR2_X1   g111(.A(KEYINPUT81), .B(G169gat), .Z(new_n313_));
  OAI221_X1 g112(.A(new_n312_), .B1(KEYINPUT82), .B2(new_n311_), .C1(new_n313_), .C2(new_n310_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(new_n303_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n293_), .A2(new_n302_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n298_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n309_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n309_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n289_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n322_), .A2(new_n289_), .A3(new_n323_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n288_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n288_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n282_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n326_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(new_n324_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n328_), .B(new_n281_), .C1(new_n332_), .C2(new_n288_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n273_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G1gat), .B(G29gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G85gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G225gat), .A2(G233gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n280_), .A2(new_n236_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT100), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n280_), .A2(new_n236_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n346_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n342_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n343_), .A2(KEYINPUT4), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n348_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n350_), .B1(new_n351_), .B2(KEYINPUT4), .ZN(new_n352_));
  AOI211_X1 g151(.A(new_n340_), .B(new_n349_), .C1(new_n352_), .C2(new_n342_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(KEYINPUT4), .ZN(new_n354_));
  INV_X1    g153(.A(new_n350_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n342_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n349_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n339_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n353_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT27), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT25), .B(G183gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n295_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n299_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT97), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(new_n301_), .A3(new_n315_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n217_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n306_), .B1(G183gat), .B2(G190gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G169gat), .ZN(new_n368_));
  INV_X1    g167(.A(G176gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n298_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT98), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n365_), .A2(new_n366_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT99), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT19), .Z(new_n378_));
  NAND2_X1  g177(.A1(new_n319_), .A2(new_n244_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n376_), .A2(KEYINPUT20), .A3(new_n378_), .A4(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT18), .ZN(new_n382_));
  XOR2_X1   g181(.A(G64gat), .B(G92gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n378_), .B(KEYINPUT96), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n319_), .A2(new_n244_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n365_), .A2(new_n373_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT20), .B1(new_n387_), .B2(new_n366_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n385_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n380_), .A2(new_n384_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n384_), .B1(new_n380_), .B2(new_n389_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n360_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n380_), .A2(new_n384_), .A3(new_n389_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT20), .ZN(new_n394_));
  INV_X1    g193(.A(new_n248_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n394_), .B1(new_n395_), .B2(new_n387_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n378_), .B1(new_n396_), .B2(new_n379_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n386_), .A2(new_n388_), .A3(new_n385_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n393_), .B(KEYINPUT27), .C1(new_n399_), .C2(new_n384_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n359_), .A2(new_n392_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n335_), .A2(KEYINPUT101), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT101), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n330_), .A2(new_n333_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n271_), .A2(new_n272_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n359_), .A2(new_n392_), .A3(new_n400_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n403_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n384_), .A2(KEYINPUT32), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n380_), .A2(new_n389_), .A3(new_n409_), .ZN(new_n410_));
  OAI221_X1 g209(.A(new_n410_), .B1(new_n399_), .B2(new_n409_), .C1(new_n353_), .C2(new_n358_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n349_), .B1(new_n352_), .B2(new_n342_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT33), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n339_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n412_), .B2(new_n339_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n390_), .A2(new_n391_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n352_), .A2(new_n341_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n339_), .B1(new_n351_), .B2(new_n342_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n411_), .B(new_n405_), .C1(new_n416_), .C2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n404_), .B1(new_n407_), .B2(new_n273_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n402_), .A2(new_n408_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G29gat), .B(G36gat), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n425_), .A2(KEYINPUT69), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(KEYINPUT69), .ZN(new_n427_));
  XOR2_X1   g226(.A(G43gat), .B(G50gat), .Z(new_n428_));
  OR3_X1    g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n428_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT15), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT74), .B(G8gat), .ZN(new_n433_));
  INV_X1    g232(.A(G1gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT14), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G15gat), .B(G22gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G1gat), .B(G8gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n435_), .A2(new_n436_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n437_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n432_), .A2(new_n438_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n438_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n431_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G229gat), .A2(G233gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT76), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n431_), .B(new_n443_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n445_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n442_), .A2(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G113gat), .B(G141gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT77), .ZN(new_n453_));
  XOR2_X1   g252(.A(G169gat), .B(G197gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n451_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n424_), .A2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G127gat), .B(G155gat), .Z(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT16), .ZN(new_n460_));
  XOR2_X1   g259(.A(G183gat), .B(G211gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT17), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G231gat), .A2(G233gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n443_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G57gat), .B(G64gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT11), .ZN(new_n468_));
  XOR2_X1   g267(.A(G71gat), .B(G78gat), .Z(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n468_), .A2(new_n469_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n467_), .A2(KEYINPUT11), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n466_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n466_), .A2(new_n473_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT17), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n464_), .B1(new_n476_), .B2(new_n462_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT75), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n478_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n477_), .B(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT37), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NOR3_X1   g282(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(KEYINPUT66), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT66), .ZN(new_n491_));
  AND3_X1   g290(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n485_), .A2(new_n490_), .A3(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(G85gat), .A2(G92gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(G85gat), .A2(G92gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT8), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n501_));
  INV_X1    g300(.A(G99gat), .ZN(new_n502_));
  INV_X1    g301(.A(G106gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n504_), .A2(new_n488_), .A3(new_n489_), .A4(new_n482_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT65), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n496_), .A2(new_n497_), .A3(KEYINPUT8), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n506_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n500_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n496_), .A2(KEYINPUT9), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT64), .B(G92gat), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n513_), .A2(G85gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n512_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT10), .B(G99gat), .Z(new_n518_));
  AOI211_X1 g317(.A(new_n493_), .B(new_n492_), .C1(new_n518_), .C2(new_n503_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n511_), .A2(new_n431_), .A3(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT70), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n505_), .A2(new_n507_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT65), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT8), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n527_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n520_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT35), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G232gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT34), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n432_), .A2(new_n529_), .B1(new_n530_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n522_), .A2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n533_), .A2(new_n530_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(KEYINPUT71), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT71), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n536_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n535_), .A2(new_n539_), .A3(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n522_), .A2(new_n534_), .A3(new_n540_), .A4(new_n536_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G190gat), .B(G218gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT72), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G134gat), .B(G162gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT36), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n543_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n481_), .B1(new_n550_), .B2(KEYINPUT73), .ZN(new_n551_));
  INV_X1    g350(.A(new_n548_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n552_), .A2(KEYINPUT36), .ZN(new_n553_));
  AOI211_X1 g352(.A(new_n538_), .B(new_n541_), .C1(new_n522_), .C2(new_n534_), .ZN(new_n554_));
  AND4_X1   g353(.A1(new_n540_), .A2(new_n522_), .A3(new_n534_), .A4(new_n536_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n553_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n550_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n551_), .A2(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n556_), .B(new_n550_), .C1(KEYINPUT73), .C2(new_n481_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n480_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n473_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n511_), .A2(new_n562_), .A3(new_n520_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n529_), .A2(KEYINPUT12), .A3(new_n473_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT67), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT67), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n529_), .A2(new_n567_), .A3(KEYINPUT12), .A4(new_n473_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n564_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT68), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n562_), .B1(new_n511_), .B2(new_n520_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n570_), .B1(new_n571_), .B2(KEYINPUT12), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n529_), .A2(new_n473_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(KEYINPUT68), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G230gat), .A2(G233gat), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n569_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  OAI211_X1 g377(.A(G230gat), .B(G233gat), .C1(new_n564_), .C2(new_n571_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G120gat), .B(G148gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT5), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G176gat), .B(G204gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n582_), .B(new_n583_), .Z(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n584_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n578_), .A2(new_n579_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT13), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n585_), .A2(KEYINPUT13), .A3(new_n587_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n561_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n458_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT102), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n359_), .A2(G1gat), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT103), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT103), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n595_), .A2(new_n599_), .A3(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n598_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n557_), .B(KEYINPUT105), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n424_), .A2(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n592_), .A2(new_n457_), .A3(new_n480_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G1gat), .B1(new_n610_), .B2(new_n359_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n604_), .A2(new_n605_), .A3(new_n611_), .ZN(G1324gat));
  AND2_X1   g411(.A1(new_n392_), .A2(new_n400_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n609_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(G8gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT39), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(new_n618_), .A3(G8gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n595_), .A2(new_n614_), .A3(new_n433_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n622_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1325gat));
  AOI21_X1  g425(.A(new_n286_), .B1(new_n609_), .B2(new_n404_), .ZN(new_n627_));
  XOR2_X1   g426(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n628_));
  OR2_X1    g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n628_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n404_), .A2(new_n286_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n629_), .B(new_n630_), .C1(new_n594_), .C2(new_n631_), .ZN(G1326gat));
  OAI21_X1  g431(.A(G22gat), .B1(new_n610_), .B2(new_n405_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT42), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n405_), .A2(G22gat), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n594_), .B2(new_n635_), .ZN(G1327gat));
  INV_X1    g435(.A(new_n480_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n592_), .A2(new_n637_), .A3(new_n557_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n458_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(G29gat), .ZN(new_n640_));
  INV_X1    g439(.A(new_n359_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n639_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT110), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT109), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n592_), .A2(new_n457_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n480_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n558_), .A2(new_n559_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT108), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT43), .B1(new_n424_), .B2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n423_), .A2(new_n422_), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT101), .B1(new_n335_), .B2(new_n401_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n406_), .A2(new_n407_), .A3(new_n403_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n651_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n558_), .A2(new_n559_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n654_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n646_), .B1(new_n650_), .B2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n644_), .B1(new_n658_), .B2(KEYINPUT44), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n656_), .A2(new_n655_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n402_), .A2(new_n408_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n662_), .B2(new_n651_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n654_), .A2(new_n648_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(KEYINPUT43), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT109), .B(new_n660_), .C1(new_n665_), .C2(new_n646_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n659_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n359_), .B1(new_n658_), .B2(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n643_), .B1(new_n669_), .B2(G29gat), .ZN(new_n670_));
  AOI211_X1 g469(.A(KEYINPUT110), .B(new_n640_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n642_), .B1(new_n670_), .B2(new_n671_), .ZN(G1328gat));
  INV_X1    g471(.A(KEYINPUT111), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n613_), .B1(new_n658_), .B2(KEYINPUT44), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n667_), .B2(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n458_), .A2(new_n676_), .A3(new_n614_), .A4(new_n638_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n679_), .A2(KEYINPUT45), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(KEYINPUT45), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n680_), .A2(new_n681_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n675_), .B1(new_n678_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n675_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n650_), .A2(new_n657_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n646_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(KEYINPUT44), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n614_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n659_), .B2(new_n666_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n685_), .B(new_n682_), .C1(new_n690_), .C2(new_n676_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n684_), .A2(new_n691_), .ZN(G1329gat));
  XNOR2_X1  g491(.A(KEYINPUT112), .B(G43gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n639_), .B2(new_n404_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n404_), .A2(G43gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n658_), .B2(KEYINPUT44), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n667_), .B2(new_n696_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g497(.A(G50gat), .B1(new_n639_), .B2(new_n273_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n688_), .A2(G50gat), .A3(new_n273_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(new_n667_), .ZN(G1331gat));
  INV_X1    g500(.A(new_n592_), .ZN(new_n702_));
  NOR4_X1   g501(.A1(new_n424_), .A2(new_n456_), .A3(new_n702_), .A4(new_n561_), .ZN(new_n703_));
  INV_X1    g502(.A(G57gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n704_), .A3(new_n641_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n592_), .A2(new_n457_), .ZN(new_n706_));
  NOR4_X1   g505(.A1(new_n424_), .A2(new_n480_), .A3(new_n606_), .A4(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(new_n641_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n708_), .B2(new_n704_), .ZN(G1332gat));
  INV_X1    g508(.A(G64gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n707_), .B2(new_n614_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n703_), .A2(new_n710_), .A3(new_n614_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1333gat));
  INV_X1    g514(.A(G71gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n707_), .B2(new_n404_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT49), .Z(new_n718_));
  NAND3_X1  g517(.A1(new_n703_), .A2(new_n716_), .A3(new_n404_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1334gat));
  INV_X1    g519(.A(G78gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n707_), .B2(new_n273_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT50), .Z(new_n723_));
  NAND3_X1  g522(.A1(new_n703_), .A2(new_n721_), .A3(new_n273_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1335gat));
  NOR2_X1   g524(.A1(new_n424_), .A2(new_n456_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n702_), .A2(new_n637_), .A3(new_n557_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(G85gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n730_), .A3(new_n641_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n706_), .A2(new_n637_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n686_), .A2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(new_n641_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n731_), .B1(new_n734_), .B2(new_n730_), .ZN(G1336gat));
  AOI21_X1  g534(.A(G92gat), .B1(new_n729_), .B2(new_n614_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n614_), .A2(new_n513_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n733_), .B2(new_n737_), .ZN(G1337gat));
  AND2_X1   g537(.A1(new_n733_), .A2(new_n404_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n404_), .A2(new_n518_), .ZN(new_n740_));
  OAI22_X1  g539(.A1(new_n739_), .A2(new_n502_), .B1(new_n728_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g541(.A1(new_n729_), .A2(new_n503_), .A3(new_n273_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n655_), .B1(new_n654_), .B2(new_n648_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n273_), .B(new_n732_), .C1(new_n744_), .C2(new_n663_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n503_), .B1(new_n745_), .B2(KEYINPUT114), .ZN(new_n746_));
  XNOR2_X1  g545(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n686_), .A2(new_n748_), .A3(new_n273_), .A4(new_n732_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n746_), .A2(new_n747_), .A3(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n747_), .B1(new_n746_), .B2(new_n749_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n743_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n743_), .B(new_n753_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1339gat));
  NAND2_X1  g556(.A1(new_n613_), .A2(new_n641_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n758_), .A2(new_n406_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n578_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n569_), .A2(new_n576_), .A3(KEYINPUT55), .ZN(new_n763_));
  NAND3_X1  g562(.A1(KEYINPUT118), .A2(G230gat), .A3(G233gat), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n569_), .A2(new_n576_), .A3(KEYINPUT55), .A4(new_n764_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n762_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n584_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT56), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(KEYINPUT56), .A3(new_n584_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n444_), .A2(new_n446_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n442_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n455_), .B1(new_n449_), .B2(new_n446_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n451_), .A2(new_n455_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n587_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT121), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(new_n587_), .A3(KEYINPUT121), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n771_), .A2(new_n772_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n656_), .B1(new_n781_), .B2(KEYINPUT58), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n780_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n768_), .A2(KEYINPUT56), .A3(new_n584_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT56), .B1(new_n768_), .B2(new_n584_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n783_), .B(KEYINPUT58), .C1(new_n784_), .C2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n588_), .A2(new_n776_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n771_), .A2(new_n790_), .A3(new_n772_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n456_), .A2(new_n587_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n785_), .B2(KEYINPUT119), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n789_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n557_), .A2(KEYINPUT57), .ZN(new_n795_));
  OAI22_X1  g594(.A1(new_n782_), .A2(new_n787_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n784_), .A2(new_n785_), .A3(KEYINPUT119), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n769_), .A2(KEYINPUT119), .A3(new_n770_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n792_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n788_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n798_), .B1(new_n803_), .B2(new_n557_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n480_), .B1(new_n796_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n560_), .A2(new_n457_), .A3(new_n702_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n807_), .A2(KEYINPUT54), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n560_), .A2(new_n457_), .A3(new_n702_), .A4(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n805_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT122), .ZN(new_n815_));
  INV_X1    g614(.A(new_n557_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n797_), .B1(new_n794_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n795_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n803_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n783_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n656_), .A3(new_n786_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n817_), .A2(new_n819_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n812_), .B1(new_n824_), .B2(new_n480_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT122), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n760_), .B1(new_n815_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(G113gat), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n456_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n814_), .A2(new_n831_), .A3(new_n832_), .A4(new_n759_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n759_), .A2(new_n832_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT123), .B1(new_n825_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n456_), .B(new_n836_), .C1(new_n828_), .C2(new_n832_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n830_), .B1(new_n838_), .B2(new_n829_), .ZN(G1340gat));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n702_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n828_), .B(new_n841_), .C1(KEYINPUT60), .C2(new_n840_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n592_), .B(new_n836_), .C1(new_n828_), .C2(new_n832_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n844_), .B2(new_n840_), .ZN(G1341gat));
  INV_X1    g644(.A(G127gat), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n480_), .A2(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n836_), .B(new_n847_), .C1(new_n828_), .C2(new_n832_), .ZN(new_n848_));
  AOI211_X1 g647(.A(KEYINPUT122), .B(new_n812_), .C1(new_n824_), .C2(new_n480_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n826_), .B1(new_n805_), .B2(new_n813_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n637_), .B(new_n759_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n846_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n851_), .B2(new_n846_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n848_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT125), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT125), .B(new_n848_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1342gat));
  AOI21_X1  g658(.A(G134gat), .B1(new_n828_), .B2(new_n606_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT126), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n861_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n828_), .A2(new_n832_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n864_), .B1(new_n835_), .B2(new_n833_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n656_), .A2(G134gat), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n862_), .A2(new_n863_), .B1(new_n865_), .B2(new_n866_), .ZN(G1343gat));
  NOR2_X1   g666(.A1(new_n404_), .A2(new_n405_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n815_), .B2(new_n827_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n758_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n457_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n224_), .ZN(G1344gat));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n702_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n225_), .ZN(G1345gat));
  AND2_X1   g675(.A1(new_n870_), .A2(new_n871_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n637_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT61), .B(G155gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  AND3_X1   g679(.A1(new_n877_), .A2(G162gat), .A3(new_n648_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G162gat), .B1(new_n877_), .B2(new_n606_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1347gat));
  NOR3_X1   g682(.A1(new_n406_), .A2(new_n613_), .A3(new_n641_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n814_), .A2(new_n884_), .ZN(new_n885_));
  OR3_X1    g684(.A1(new_n885_), .A2(KEYINPUT127), .A3(new_n457_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT127), .B1(new_n885_), .B2(new_n457_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(G169gat), .A3(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n885_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n368_), .A3(new_n456_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n888_), .A2(new_n889_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n890_), .A2(new_n892_), .A3(new_n893_), .ZN(G1348gat));
  AOI21_X1  g693(.A(G176gat), .B1(new_n891_), .B2(new_n592_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n273_), .B1(new_n815_), .B2(new_n827_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n613_), .A2(new_n641_), .ZN(new_n897_));
  AND4_X1   g696(.A1(G176gat), .A2(new_n897_), .A3(new_n404_), .A4(new_n592_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n895_), .B1(new_n896_), .B2(new_n898_), .ZN(G1349gat));
  NOR3_X1   g698(.A1(new_n885_), .A2(new_n361_), .A3(new_n480_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n896_), .A2(new_n404_), .A3(new_n637_), .A4(new_n897_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n293_), .ZN(G1350gat));
  OAI21_X1  g701(.A(G190gat), .B1(new_n885_), .B2(new_n647_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n606_), .A2(new_n295_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n885_), .B2(new_n904_), .ZN(G1351gat));
  NAND2_X1  g704(.A1(new_n870_), .A2(new_n897_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n457_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n207_), .ZN(G1352gat));
  NOR2_X1   g707(.A1(new_n906_), .A2(new_n702_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(new_n203_), .ZN(G1353gat));
  XNOR2_X1  g709(.A(KEYINPUT63), .B(G211gat), .ZN(new_n911_));
  OR2_X1    g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n870_), .A2(new_n637_), .A3(new_n897_), .ZN(new_n913_));
  MUX2_X1   g712(.A(new_n911_), .B(new_n912_), .S(new_n913_), .Z(G1354gat));
  OAI21_X1  g713(.A(G218gat), .B1(new_n906_), .B2(new_n647_), .ZN(new_n915_));
  INV_X1    g714(.A(G218gat), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n606_), .A2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n906_), .B2(new_n917_), .ZN(G1355gat));
endmodule


