//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT9), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT9), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n203_), .A2(new_n206_), .A3(new_n208_), .A4(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT8), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n207_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n215_), .B(new_n216_), .C1(new_n218_), .C2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n221_));
  AND3_X1   g020(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT65), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n221_), .B(new_n217_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NOR3_X1   g025(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n220_), .A2(new_n224_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n213_), .B1(new_n229_), .B2(new_n202_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n202_), .A2(new_n213_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(new_n208_), .B2(new_n228_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n212_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(KEYINPUT66), .B(new_n212_), .C1(new_n230_), .C2(new_n232_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G71gat), .B(G78gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G57gat), .A2(G64gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT11), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G57gat), .A2(G64gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT11), .B1(new_n244_), .B2(new_n239_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n238_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n237_), .B(KEYINPUT11), .C1(new_n239_), .C2(new_n244_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n247_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n235_), .A2(new_n236_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT12), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n235_), .A2(new_n236_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n252_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G230gat), .A2(G233gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n246_), .A2(new_n248_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n247_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(KEYINPUT69), .A3(new_n249_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n261_), .A2(new_n233_), .A3(new_n265_), .A4(KEYINPUT12), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n256_), .A2(new_n258_), .A3(new_n259_), .A4(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n258_), .A2(new_n254_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(new_n259_), .ZN(new_n269_));
  XOR2_X1   g068(.A(KEYINPUT5), .B(G176gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT70), .B(G204gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G120gat), .B(G148gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n269_), .A2(new_n274_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT13), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n276_), .A2(KEYINPUT13), .A3(new_n277_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(KEYINPUT71), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G113gat), .B(G141gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G169gat), .B(G197gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G1gat), .B(G8gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT77), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G15gat), .ZN(new_n291_));
  INV_X1    g090(.A(G22gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G15gat), .A2(G22gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G1gat), .A2(G8gat), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n293_), .A2(new_n294_), .B1(KEYINPUT14), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n290_), .B(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(KEYINPUT72), .B(KEYINPUT73), .Z(new_n298_));
  XNOR2_X1  g097(.A(G43gat), .B(G50gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G43gat), .B(G50gat), .Z(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G29gat), .B(G36gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n300_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n297_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT15), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n300_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n305_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n307_), .A2(KEYINPUT15), .A3(new_n308_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n310_), .B1(new_n297_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G229gat), .A2(G233gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n297_), .B(new_n309_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n318_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT82), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(KEYINPUT81), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n324_), .B1(new_n323_), .B2(KEYINPUT81), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n287_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(new_n286_), .A3(new_n325_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n281_), .A2(new_n280_), .A3(KEYINPUT71), .ZN(new_n333_));
  NOR3_X1   g132(.A1(new_n283_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G127gat), .B(G134gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G113gat), .B(G120gat), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT89), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n336_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT88), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT31), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT87), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT83), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT24), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(G169gat), .B2(G176gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT25), .B(G183gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT26), .B(G190gat), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n347_), .A2(new_n349_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n352_), .A2(KEYINPUT84), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n347_), .A2(KEYINPUT24), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(G183gat), .B2(G190gat), .ZN(new_n356_));
  INV_X1    g155(.A(G183gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(KEYINPUT23), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n356_), .B1(G190gat), .B2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n354_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n352_), .A2(KEYINPUT84), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n353_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n356_), .B(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n358_), .A2(G190gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(G183gat), .B2(G190gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT85), .B(G176gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT22), .B(G169gat), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n368_), .A2(new_n369_), .B1(G169gat), .B2(G176gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n362_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373_));
  INV_X1    g172(.A(G71gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n375_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n362_), .B2(new_n371_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n345_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G15gat), .B(G43gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT30), .B(G99gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n381_), .B(new_n382_), .Z(new_n383_));
  OAI211_X1 g182(.A(new_n344_), .B(KEYINPUT87), .C1(new_n376_), .C2(new_n378_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n380_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(new_n210_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT18), .B(G64gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G226gat), .A2(G233gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT19), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G197gat), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n397_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT90), .ZN(new_n399_));
  INV_X1    g198(.A(G204gat), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(G197gat), .B2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(G197gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n398_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(G211gat), .B(G218gat), .Z(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(KEYINPUT21), .A3(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT92), .ZN(new_n406_));
  OR3_X1    g205(.A1(new_n403_), .A2(KEYINPUT91), .A3(KEYINPUT21), .ZN(new_n407_));
  XOR2_X1   g206(.A(G197gat), .B(G204gat), .Z(new_n408_));
  AOI21_X1  g207(.A(new_n404_), .B1(KEYINPUT21), .B2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT91), .B1(new_n403_), .B2(KEYINPUT21), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n407_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n406_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n346_), .A2(new_n348_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n366_), .A2(new_n352_), .A3(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G183gat), .A2(G190gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n370_), .B1(new_n359_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n412_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT20), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n419_), .A2(KEYINPUT98), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(KEYINPUT98), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT99), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n422_), .A2(new_n423_), .B1(new_n372_), .B2(new_n412_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n396_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n419_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(new_n372_), .B2(new_n412_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n428_), .A2(new_n395_), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT32), .B(new_n393_), .C1(new_n426_), .C2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT100), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G225gat), .A2(G233gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT4), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G155gat), .A2(G162gat), .ZN(new_n435_));
  OR2_X1    g234(.A1(G155gat), .A2(G162gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G141gat), .A2(G148gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT3), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G141gat), .A2(G148gat), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT2), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n435_), .B(new_n436_), .C1(new_n439_), .C2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n437_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n435_), .A2(KEYINPUT1), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n436_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n435_), .A2(KEYINPUT1), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n444_), .B(new_n440_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n443_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n342_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n337_), .A2(new_n340_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n443_), .A2(new_n451_), .A3(new_n448_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n434_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT4), .B1(new_n342_), .B2(new_n449_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n433_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(new_n432_), .A3(new_n452_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G1gat), .B(G29gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(G85gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT0), .B(G57gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n459_), .B(new_n460_), .Z(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n431_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n455_), .A2(new_n456_), .A3(new_n461_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n464_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n372_), .A2(new_n412_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n467_), .A2(new_n418_), .A3(KEYINPUT20), .A4(new_n396_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n372_), .A2(new_n412_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n396_), .B1(new_n470_), .B2(new_n427_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT32), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n472_), .B1(new_n473_), .B2(new_n392_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n430_), .A2(new_n465_), .A3(new_n466_), .A4(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n392_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT97), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n428_), .A2(new_n395_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n393_), .A3(new_n468_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n472_), .A2(KEYINPUT97), .A3(new_n393_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n432_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n450_), .A2(new_n433_), .A3(new_n452_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n462_), .A3(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n464_), .B(KEYINPUT33), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n388_), .B1(new_n475_), .B2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n449_), .A2(KEYINPUT29), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n489_), .B(KEYINPUT28), .Z(new_n490_));
  XNOR2_X1  g289(.A(G22gat), .B(G50gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n449_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT94), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n412_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G228gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G78gat), .B(G106gat), .Z(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n449_), .B2(KEYINPUT29), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n412_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n500_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n501_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n498_), .B1(new_n496_), .B2(new_n412_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n503_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n492_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n504_), .A2(KEYINPUT95), .A3(new_n508_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n492_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT95), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n500_), .A2(new_n512_), .A3(new_n501_), .A4(new_n503_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT96), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT96), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n510_), .A2(new_n516_), .A3(new_n511_), .A4(new_n513_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n509_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n488_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n388_), .ZN(new_n520_));
  AOI211_X1 g319(.A(new_n509_), .B(new_n387_), .C1(new_n515_), .C2(new_n517_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT27), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n480_), .A2(new_n523_), .A3(new_n481_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT101), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n480_), .A2(new_n481_), .A3(KEYINPUT101), .A4(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n465_), .A2(new_n466_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n392_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(KEYINPUT27), .A3(new_n479_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n528_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n519_), .B1(new_n522_), .B2(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n334_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G190gat), .B(G218gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G134gat), .B(G162gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT36), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n539_), .B(KEYINPUT34), .Z(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n316_), .A2(new_n233_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n309_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n543_), .B2(new_n257_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT35), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n541_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n257_), .A2(new_n543_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n542_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n547_), .A2(new_n548_), .A3(KEYINPUT74), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n540_), .A2(KEYINPUT35), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n546_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n544_), .A2(KEYINPUT74), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n547_), .A2(new_n548_), .A3(new_n545_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n540_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n550_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n552_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n538_), .B1(new_n551_), .B2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n549_), .B1(new_n546_), .B2(new_n550_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n537_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(KEYINPUT36), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n554_), .A2(new_n552_), .A3(new_n555_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n558_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n252_), .B(new_n564_), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(new_n297_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G127gat), .B(G155gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(G211gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT16), .B(G183gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n570_), .A2(KEYINPUT17), .ZN(new_n571_));
  XOR2_X1   g370(.A(KEYINPUT69), .B(KEYINPUT78), .Z(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(KEYINPUT17), .A3(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n566_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n566_), .A2(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n534_), .A2(new_n563_), .A3(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(G1gat), .B1(new_n578_), .B2(new_n529_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT102), .Z(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT75), .B(KEYINPUT37), .Z(new_n581_));
  NAND3_X1  g380(.A1(new_n557_), .A2(new_n562_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT76), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n563_), .A2(KEYINPUT37), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT76), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n557_), .A2(new_n585_), .A3(new_n562_), .A4(new_n581_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n583_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n577_), .B(KEYINPUT79), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT80), .Z(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n534_), .ZN(new_n591_));
  OR3_X1    g390(.A1(new_n591_), .A2(G1gat), .A3(new_n529_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(KEYINPUT103), .A2(KEYINPUT38), .ZN(new_n593_));
  AND2_X1   g392(.A1(KEYINPUT103), .A2(KEYINPUT38), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n592_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n580_), .B(new_n595_), .C1(new_n593_), .C2(new_n592_), .ZN(G1324gat));
  NAND2_X1  g395(.A1(new_n528_), .A2(new_n531_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n591_), .A2(G8gat), .A3(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT104), .ZN(new_n600_));
  OAI21_X1  g399(.A(G8gat), .B1(new_n578_), .B2(new_n598_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT39), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT40), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(new_n602_), .A3(KEYINPUT40), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(G1325gat));
  OAI21_X1  g406(.A(G15gat), .B1(new_n578_), .B2(new_n387_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT41), .Z(new_n609_));
  INV_X1    g408(.A(new_n591_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n291_), .A3(new_n388_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(G1326gat));
  OAI21_X1  g411(.A(G22gat), .B1(new_n578_), .B2(new_n518_), .ZN(new_n613_));
  XOR2_X1   g412(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n518_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n610_), .A2(new_n292_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(G1327gat));
  NOR2_X1   g417(.A1(new_n588_), .A2(new_n563_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n534_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n529_), .ZN(new_n622_));
  AOI21_X1  g421(.A(G29gat), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n588_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n518_), .B(new_n388_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n528_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n626_));
  AOI22_X1  g425(.A1(new_n625_), .A2(new_n626_), .B1(new_n518_), .B2(new_n488_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n627_), .A2(KEYINPUT43), .A3(new_n587_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT43), .ZN(new_n629_));
  INV_X1    g428(.A(new_n587_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n533_), .B2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n334_), .B(new_n624_), .C1(new_n628_), .C2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT44), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT43), .B1(new_n627_), .B2(new_n587_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n533_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n637_), .A2(KEYINPUT44), .A3(new_n334_), .A4(new_n624_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n634_), .A2(G29gat), .A3(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n623_), .B1(new_n639_), .B2(new_n622_), .ZN(G1328gat));
  NAND3_X1  g439(.A1(new_n634_), .A2(new_n597_), .A3(new_n638_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G36gat), .ZN(new_n642_));
  INV_X1    g441(.A(G36gat), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n534_), .A2(new_n597_), .A3(new_n643_), .A4(new_n619_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT45), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT46), .B1(new_n646_), .B2(KEYINPUT106), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT46), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n648_), .B(new_n649_), .C1(new_n642_), .C2(new_n645_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n647_), .A2(new_n650_), .ZN(G1329gat));
  NOR3_X1   g450(.A1(new_n620_), .A2(G43gat), .A3(new_n387_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n634_), .A2(new_n388_), .A3(new_n638_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n653_), .B2(G43gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT47), .ZN(G1330gat));
  AND4_X1   g454(.A1(G50gat), .A2(new_n634_), .A3(new_n616_), .A4(new_n638_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G50gat), .B1(new_n621_), .B2(new_n616_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1331gat));
  OR2_X1    g457(.A1(new_n283_), .A2(new_n333_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n660_), .A2(new_n331_), .A3(new_n627_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n563_), .A3(new_n588_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT108), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n663_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n664_), .A2(G57gat), .A3(new_n622_), .A4(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n661_), .A2(new_n590_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n622_), .ZN(new_n668_));
  INV_X1    g467(.A(G57gat), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n668_), .A2(KEYINPUT107), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT107), .B1(new_n668_), .B2(new_n669_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n666_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT109), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT109), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n666_), .B(new_n674_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1332gat));
  INV_X1    g475(.A(G64gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n667_), .A2(new_n677_), .A3(new_n597_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n664_), .A2(new_n597_), .A3(new_n665_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT48), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(new_n680_), .A3(G64gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n679_), .B2(G64gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(G1333gat));
  NOR2_X1   g482(.A1(new_n387_), .A2(G71gat), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT110), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n667_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n664_), .A2(new_n388_), .A3(new_n665_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT49), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n687_), .A2(new_n688_), .A3(G71gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n687_), .B2(G71gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(G1334gat));
  INV_X1    g490(.A(G78gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n667_), .A2(new_n692_), .A3(new_n616_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n664_), .A2(new_n616_), .A3(new_n665_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT50), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(new_n695_), .A3(G78gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n694_), .B2(G78gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(G1335gat));
  AND2_X1   g497(.A1(new_n661_), .A2(new_n619_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G85gat), .B1(new_n699_), .B2(new_n622_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT111), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n660_), .A2(new_n331_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n637_), .A2(new_n624_), .A3(new_n702_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n703_), .A2(KEYINPUT112), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(KEYINPUT112), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n209_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n701_), .B1(new_n622_), .B2(new_n706_), .ZN(G1336gat));
  NAND3_X1  g506(.A1(new_n699_), .A2(new_n210_), .A3(new_n597_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n598_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n210_), .ZN(G1337gat));
  OAI21_X1  g509(.A(G99gat), .B1(new_n703_), .B2(new_n387_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n699_), .A2(new_n204_), .A3(new_n388_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n711_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n714_), .B(new_n715_), .Z(G1338gat));
  NAND4_X1  g515(.A1(new_n637_), .A2(new_n616_), .A3(new_n624_), .A4(new_n702_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT114), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT52), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n717_), .A2(G106gat), .A3(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n718_), .A2(KEYINPUT52), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n699_), .A2(new_n205_), .A3(new_n616_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n721_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n717_), .A2(G106gat), .A3(new_n724_), .A4(new_n719_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n722_), .A2(new_n723_), .A3(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(G1339gat));
  INV_X1    g527(.A(KEYINPUT55), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n267_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n253_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n731_));
  AND4_X1   g530(.A1(KEYINPUT12), .A2(new_n261_), .A3(new_n265_), .A4(new_n233_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n733_), .A2(KEYINPUT55), .A3(new_n259_), .A4(new_n256_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT117), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n256_), .A2(new_n258_), .A3(new_n266_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n259_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  AOI211_X1 g538(.A(KEYINPUT117), .B(new_n259_), .C1(new_n733_), .C2(new_n256_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n735_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n274_), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT56), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n737_), .A2(new_n738_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT117), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n737_), .A2(new_n736_), .A3(new_n738_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n745_), .A2(new_n746_), .A3(new_n730_), .A4(new_n734_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT56), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n274_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n743_), .A2(new_n331_), .A3(new_n276_), .A4(new_n749_), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n317_), .A2(new_n318_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n320_), .A2(new_n321_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n287_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n323_), .A2(new_n286_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n278_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n750_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n563_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT57), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT57), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n757_), .A2(new_n760_), .A3(new_n563_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n747_), .A2(new_n748_), .A3(new_n274_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n748_), .B1(new_n747_), .B2(new_n274_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n275_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n765_), .A2(KEYINPUT118), .A3(KEYINPUT58), .A4(new_n755_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n743_), .A2(new_n276_), .A3(new_n755_), .A4(new_n749_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT58), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n769_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n766_), .A2(new_n770_), .A3(new_n630_), .A4(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n577_), .B1(new_n762_), .B2(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n587_), .A2(new_n332_), .A3(new_n282_), .A4(new_n588_), .ZN(new_n774_));
  XOR2_X1   g573(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(new_n774_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT119), .B1(new_n773_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n630_), .A2(new_n771_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n766_), .A2(new_n770_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n760_), .B1(new_n757_), .B2(new_n563_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n563_), .ZN(new_n783_));
  AOI211_X1 g582(.A(KEYINPUT57), .B(new_n783_), .C1(new_n750_), .C2(new_n756_), .ZN(new_n784_));
  OAI22_X1  g583(.A1(new_n780_), .A2(new_n781_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n577_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n778_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n787_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n597_), .A2(new_n529_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n779_), .A2(new_n790_), .A3(new_n521_), .A4(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n521_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n785_), .A2(new_n624_), .ZN(new_n794_));
  AOI211_X1 g593(.A(KEYINPUT59), .B(new_n793_), .C1(new_n794_), .C2(new_n788_), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n792_), .A2(KEYINPUT59), .B1(new_n795_), .B2(KEYINPUT120), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n795_), .A2(KEYINPUT120), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n796_), .A2(G113gat), .A3(new_n797_), .A4(new_n331_), .ZN(new_n798_));
  INV_X1    g597(.A(G113gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n792_), .B2(new_n332_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1340gat));
  NAND3_X1  g600(.A1(new_n796_), .A2(new_n659_), .A3(new_n797_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(G120gat), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT60), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n804_), .A2(G120gat), .ZN(new_n805_));
  AOI21_X1  g604(.A(G120gat), .B1(new_n659_), .B2(new_n804_), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n806_), .B(KEYINPUT121), .Z(new_n807_));
  OR3_X1    g606(.A1(new_n792_), .A2(new_n805_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n803_), .A2(new_n808_), .ZN(G1341gat));
  NAND4_X1  g608(.A1(new_n796_), .A2(G127gat), .A3(new_n797_), .A4(new_n577_), .ZN(new_n810_));
  INV_X1    g609(.A(G127gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n792_), .B2(new_n624_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1342gat));
  XNOR2_X1  g612(.A(KEYINPUT122), .B(G134gat), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n796_), .A2(new_n630_), .A3(new_n797_), .A4(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(G134gat), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n792_), .B2(new_n563_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1343gat));
  NAND4_X1  g617(.A1(new_n779_), .A2(new_n790_), .A3(new_n520_), .A4(new_n791_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT123), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n819_), .A2(new_n820_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n331_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(G141gat), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n773_), .A2(KEYINPUT119), .A3(new_n778_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n789_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n827_), .A2(KEYINPUT123), .A3(new_n520_), .A4(new_n791_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n819_), .A2(new_n820_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(G141gat), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n331_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n824_), .A2(new_n832_), .ZN(G1344gat));
  OAI21_X1  g632(.A(new_n659_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(G148gat), .ZN(new_n835_));
  INV_X1    g634(.A(G148gat), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n830_), .A2(new_n836_), .A3(new_n659_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(G1345gat));
  XNOR2_X1  g637(.A(KEYINPUT61), .B(G155gat), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n830_), .B2(new_n588_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n839_), .ZN(new_n841_));
  AOI211_X1 g640(.A(new_n624_), .B(new_n841_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1346gat));
  AOI21_X1  g642(.A(G162gat), .B1(new_n830_), .B2(new_n783_), .ZN(new_n844_));
  INV_X1    g643(.A(G162gat), .ZN(new_n845_));
  AOI211_X1 g644(.A(new_n845_), .B(new_n587_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1347gat));
  INV_X1    g646(.A(G169gat), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n794_), .A2(new_n788_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n598_), .A2(new_n622_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n388_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n849_), .A2(new_n518_), .A3(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n332_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  OR4_X1    g657(.A1(new_n848_), .A2(new_n854_), .A3(new_n855_), .A4(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n854_), .A2(new_n369_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n856_), .B(new_n857_), .C1(new_n854_), .C2(new_n848_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(G1348gat));
  AND3_X1   g661(.A1(new_n852_), .A2(G176gat), .A3(new_n659_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n827_), .A2(new_n518_), .A3(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n368_), .B1(new_n853_), .B2(new_n660_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1349gat));
  NOR3_X1   g665(.A1(new_n853_), .A2(new_n350_), .A3(new_n786_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n827_), .A2(new_n518_), .A3(new_n588_), .A4(new_n852_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n357_), .ZN(G1350gat));
  OAI21_X1  g668(.A(G190gat), .B1(new_n853_), .B2(new_n587_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n849_), .A2(new_n351_), .A3(new_n518_), .A4(new_n852_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n563_), .ZN(G1351gat));
  NAND3_X1  g671(.A1(new_n827_), .A2(new_n520_), .A3(new_n850_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n332_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(new_n397_), .ZN(G1352gat));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n660_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n400_), .ZN(G1353gat));
  NAND2_X1  g676(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n577_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n873_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT125), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n880_), .B(new_n882_), .ZN(G1354gat));
  XOR2_X1   g682(.A(KEYINPUT126), .B(G218gat), .Z(new_n884_));
  NOR3_X1   g683(.A1(new_n873_), .A2(new_n587_), .A3(new_n884_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n873_), .A2(new_n563_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n884_), .ZN(G1355gat));
endmodule


