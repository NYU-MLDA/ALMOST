//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_;
  INV_X1    g000(.A(G183gat), .ZN(new_n202_));
  OAI21_X1  g001(.A(KEYINPUT25), .B1(new_n202_), .B2(KEYINPUT78), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT25), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(G183gat), .ZN(new_n206_));
  AND3_X1   g005(.A1(KEYINPUT79), .A2(KEYINPUT26), .A3(G190gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT26), .B1(KEYINPUT79), .B2(G190gat), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n203_), .B(new_n206_), .C1(new_n207_), .C2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n217_), .A2(KEYINPUT24), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n209_), .A2(new_n214_), .A3(new_n218_), .A4(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(G169gat), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n212_), .B(new_n213_), .C1(G183gat), .C2(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G211gat), .B(G218gat), .Z(new_n226_));
  INV_X1    g025(.A(G197gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(G204gat), .ZN(new_n228_));
  INV_X1    g027(.A(G204gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(G197gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n226_), .B(KEYINPUT21), .C1(new_n228_), .C2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT21), .B1(new_n228_), .B2(new_n230_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(G197gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(G204gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT21), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G211gat), .B(G218gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n232_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n221_), .A2(new_n225_), .A3(new_n231_), .A4(new_n238_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n239_), .A2(KEYINPUT88), .A3(KEYINPUT20), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT88), .B1(new_n239_), .B2(KEYINPUT20), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n217_), .A2(new_n219_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT25), .B(G183gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT26), .B(G190gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n244_), .A2(new_n214_), .A3(new_n247_), .A4(new_n248_), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n249_), .A2(new_n225_), .B1(new_n231_), .B2(new_n238_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n240_), .A2(new_n241_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT19), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT87), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT90), .B1(new_n251_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n221_), .A2(new_n225_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n238_), .A2(new_n231_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n249_), .A2(new_n225_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n258_), .B(KEYINPUT20), .C1(new_n259_), .C2(new_n257_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n260_), .A2(new_n253_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n241_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n250_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n239_), .A2(KEYINPUT88), .A3(KEYINPUT20), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT90), .ZN(new_n266_));
  INV_X1    g065(.A(new_n254_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n255_), .A2(new_n261_), .A3(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G8gat), .B(G36gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G64gat), .B(G92gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n274_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n255_), .A2(new_n268_), .A3(new_n261_), .A4(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(KEYINPUT92), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT27), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n255_), .A2(new_n268_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT92), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n261_), .A4(new_n276_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n278_), .A2(new_n279_), .A3(new_n282_), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n251_), .A2(new_n254_), .B1(new_n253_), .B2(new_n260_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n277_), .B(KEYINPUT27), .C1(new_n276_), .C2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n257_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT84), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT84), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(G155gat), .A3(G162gat), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n288_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n287_), .B1(new_n293_), .B2(KEYINPUT85), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n291_), .B1(G155gat), .B2(G162gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n289_), .A2(KEYINPUT84), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT1), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT85), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n290_), .A2(new_n292_), .A3(new_n288_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n294_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n302_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n308_), .A2(new_n310_), .A3(new_n311_), .A4(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n290_), .A2(new_n292_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n287_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n306_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n286_), .B1(new_n318_), .B2(KEYINPUT29), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n316_), .B1(new_n301_), .B2(new_n305_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n321_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G228gat), .A2(G233gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n286_), .B2(KEYINPUT86), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n324_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT28), .B1(new_n318_), .B2(KEYINPUT29), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n329_), .B1(new_n330_), .B2(new_n323_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n319_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G22gat), .B(G50gat), .ZN(new_n333_));
  INV_X1    g132(.A(G106gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G78gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n327_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n319_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n330_), .A2(new_n323_), .A3(new_n329_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n332_), .A2(new_n336_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n336_), .B1(new_n332_), .B2(new_n340_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n283_), .A2(new_n285_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT98), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT83), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT30), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n256_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G99gat), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n350_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G227gat), .A2(G233gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n353_), .B(G15gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(G71gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT80), .B(G43gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n351_), .A2(new_n352_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n357_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n347_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n349_), .B(new_n350_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n357_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(KEYINPUT83), .A3(new_n358_), .ZN(new_n365_));
  INV_X1    g164(.A(G127gat), .ZN(new_n366_));
  INV_X1    g165(.A(G134gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G127gat), .A2(G134gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(G113gat), .ZN(new_n371_));
  INV_X1    g170(.A(G120gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G113gat), .A2(G120gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n370_), .A2(new_n375_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n368_), .A2(new_n373_), .A3(new_n369_), .A4(new_n374_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT81), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT81), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n382_), .B(new_n383_), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n361_), .A2(new_n365_), .A3(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n364_), .A2(KEYINPUT83), .A3(new_n358_), .A4(new_n384_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G1gat), .B(G29gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G57gat), .B(G85gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n382_), .B1(new_n306_), .B2(new_n317_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n378_), .ZN(new_n397_));
  AOI211_X1 g196(.A(new_n397_), .B(new_n316_), .C1(new_n301_), .C2(new_n305_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT4), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n320_), .B2(new_n382_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n395_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n320_), .A2(new_n378_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n382_), .B2(new_n320_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n395_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n394_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT96), .ZN(new_n408_));
  INV_X1    g207(.A(new_n406_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n399_), .A2(new_n401_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n409_), .B(new_n393_), .C1(new_n410_), .C2(new_n395_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT96), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n412_), .B(new_n394_), .C1(new_n402_), .C2(new_n406_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n408_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT97), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n408_), .A2(KEYINPUT97), .A3(new_n411_), .A4(new_n413_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n388_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n345_), .A2(new_n346_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n346_), .B1(new_n345_), .B2(new_n418_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n278_), .A2(new_n282_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n394_), .B1(new_n404_), .B2(new_n395_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT95), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT94), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n411_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT33), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n411_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n421_), .A2(new_n424_), .A3(new_n427_), .A4(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n336_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n340_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n338_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n341_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n276_), .A2(KEYINPUT32), .ZN(new_n436_));
  MUX2_X1   g235(.A(new_n284_), .B(new_n269_), .S(new_n436_), .Z(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n414_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n430_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n388_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n283_), .A2(new_n285_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n416_), .A2(new_n417_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n344_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  OAI22_X1  g242(.A1(new_n419_), .A2(new_n420_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G190gat), .B(G218gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G134gat), .B(G162gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT36), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(KEYINPUT10), .B(G99gat), .Z(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n334_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT6), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT9), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(G85gat), .A3(G92gat), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n453_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G85gat), .B(G92gat), .Z(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT9), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT7), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n462_), .A2(KEYINPUT64), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT64), .ZN(new_n464_));
  OAI22_X1  g263(.A1(new_n464_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n462_), .A2(new_n350_), .A3(new_n334_), .A4(KEYINPUT64), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n455_), .A2(new_n463_), .A3(new_n465_), .A4(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n467_), .A2(new_n459_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n468_), .B1(new_n467_), .B2(new_n459_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n461_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G29gat), .B(G36gat), .ZN(new_n472_));
  INV_X1    g271(.A(G43gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G50gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n472_), .B(G43gat), .ZN(new_n476_));
  INV_X1    g275(.A(G50gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n471_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n481_));
  INV_X1    g280(.A(new_n471_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n475_), .A2(new_n478_), .A3(KEYINPUT15), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT15), .B1(new_n475_), .B2(new_n478_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n480_), .B(new_n481_), .C1(new_n482_), .C2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G232gat), .A2(G233gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n487_), .B(KEYINPUT34), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n485_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n471_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(KEYINPUT71), .A3(new_n480_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n488_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n481_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n489_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n492_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n451_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n489_), .A2(new_n494_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n492_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n449_), .A2(KEYINPUT36), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n489_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n444_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT100), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n444_), .A2(KEYINPUT100), .A3(new_n504_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510_));
  INV_X1    g309(.A(G1gat), .ZN(new_n511_));
  INV_X1    g310(.A(G8gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT14), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G1gat), .B(G8gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G231gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G71gat), .B(G78gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n518_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G183gat), .B(G211gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G127gat), .B(G155gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT17), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n525_), .A2(new_n531_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n530_), .A2(KEYINPUT17), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n525_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n479_), .A2(new_n516_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n490_), .B2(new_n516_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n479_), .B(new_n516_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(G229gat), .A3(G233gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n215_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(new_n227_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n543_), .A2(new_n546_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT69), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT12), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n552_), .A2(KEYINPUT68), .ZN(new_n553_));
  INV_X1    g352(.A(new_n524_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n553_), .B1(new_n471_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n524_), .B(new_n461_), .C1(new_n470_), .C2(new_n469_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G230gat), .A2(G233gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT68), .B(KEYINPUT12), .Z(new_n559_));
  NAND3_X1  g358(.A1(new_n471_), .A2(new_n554_), .A3(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .A4(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n471_), .A2(new_n554_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT66), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n482_), .A2(new_n565_), .A3(new_n524_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n557_), .A2(KEYINPUT66), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n564_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT67), .ZN(new_n570_));
  INV_X1    g369(.A(new_n558_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT67), .B1(new_n568_), .B2(new_n558_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n562_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT5), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(G176gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n229_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n574_), .A2(new_n579_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT13), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n574_), .A2(new_n579_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT13), .B1(new_n585_), .B2(new_n580_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n551_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n583_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(KEYINPUT13), .A3(new_n580_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(KEYINPUT69), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n550_), .B1(new_n587_), .B2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n509_), .A2(new_n536_), .A3(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G1gat), .B1(new_n592_), .B2(new_n442_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT75), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n451_), .A2(KEYINPUT74), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n451_), .A2(KEYINPUT74), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n595_), .B(new_n596_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n503_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n594_), .B1(new_n598_), .B2(KEYINPUT37), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT37), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n497_), .A2(new_n503_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n535_), .B(KEYINPUT77), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n601_), .A2(KEYINPUT75), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n602_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(new_n591_), .A3(new_n444_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n442_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n511_), .A3(new_n610_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n611_), .A2(KEYINPUT99), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT38), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(KEYINPUT99), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n612_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n613_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n593_), .B1(new_n615_), .B2(new_n616_), .ZN(G1324gat));
  INV_X1    g416(.A(KEYINPUT40), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n619_));
  INV_X1    g418(.A(new_n441_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n509_), .A2(new_n536_), .A3(new_n591_), .A4(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(G8gat), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT39), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n621_), .A2(new_n624_), .A3(G8gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n609_), .A2(new_n512_), .A3(new_n620_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n619_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n621_), .A2(new_n624_), .A3(G8gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n624_), .B1(new_n621_), .B2(G8gat), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n619_), .B(new_n627_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n618_), .B1(new_n628_), .B2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n627_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT101), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(KEYINPUT40), .A3(new_n631_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(G1325gat));
  OR3_X1    g436(.A1(new_n608_), .A2(G15gat), .A3(new_n388_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G15gat), .B1(new_n592_), .B2(new_n388_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT41), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n639_), .A2(new_n640_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n638_), .B1(new_n641_), .B2(new_n642_), .ZN(G1326gat));
  OR3_X1    g442(.A1(new_n608_), .A2(G22gat), .A3(new_n344_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n592_), .A2(new_n344_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G22gat), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT103), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n648_), .A3(G22gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n647_), .A2(new_n649_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n644_), .B1(new_n652_), .B2(new_n653_), .ZN(G1327gat));
  NOR2_X1   g453(.A1(new_n504_), .A2(new_n603_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n591_), .A2(new_n444_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n610_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n604_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n444_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n444_), .A2(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT43), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n444_), .A2(KEYINPUT104), .A3(new_n658_), .A4(new_n660_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n663_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n603_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n591_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(KEYINPUT44), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G29gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT44), .B1(new_n667_), .B2(new_n669_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n657_), .B1(new_n673_), .B2(new_n610_), .ZN(G1328gat));
  NAND2_X1  g473(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(G36gat), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n441_), .B(KEYINPUT105), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n656_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT106), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n656_), .A2(new_n683_), .A3(new_n679_), .A4(new_n680_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n682_), .A2(KEYINPUT45), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT45), .B1(new_n682_), .B2(new_n684_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n672_), .A2(new_n441_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n679_), .B1(new_n689_), .B2(new_n670_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n675_), .B(new_n678_), .C1(new_n688_), .C2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n670_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G36gat), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n693_), .A2(new_n687_), .A3(new_n676_), .A4(new_n677_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1329gat));
  INV_X1    g494(.A(new_n388_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n656_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n473_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n670_), .A2(G43gat), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700_));
  NOR4_X1   g499(.A1(new_n699_), .A2(new_n672_), .A3(new_n700_), .A4(new_n388_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n670_), .A2(G43gat), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n667_), .A2(new_n669_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n388_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT108), .B1(new_n702_), .B2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n698_), .B1(new_n701_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT47), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n709_), .B(new_n698_), .C1(new_n701_), .C2(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n656_), .B2(new_n435_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n672_), .A2(new_n477_), .A3(new_n344_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n670_), .ZN(G1331gat));
  INV_X1    g513(.A(G57gat), .ZN(new_n715_));
  INV_X1    g514(.A(new_n590_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT69), .B1(new_n588_), .B2(new_n589_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n549_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n718_), .A2(new_n444_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n607_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT109), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n715_), .B1(new_n721_), .B2(new_n442_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n509_), .A2(new_n603_), .A3(new_n718_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(G57gat), .A3(new_n610_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT110), .Z(G1332gat));
  INV_X1    g525(.A(new_n680_), .ZN(new_n727_));
  OR3_X1    g526(.A1(new_n720_), .A2(G64gat), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n723_), .A2(new_n680_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(G64gat), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(KEYINPUT48), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(KEYINPUT48), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(G1333gat));
  OR3_X1    g532(.A1(new_n720_), .A2(G71gat), .A3(new_n388_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n723_), .A2(new_n696_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G71gat), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(KEYINPUT49), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(KEYINPUT49), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1334gat));
  OR3_X1    g538(.A1(new_n720_), .A2(G78gat), .A3(new_n344_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n723_), .A2(new_n435_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G78gat), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(KEYINPUT50), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(KEYINPUT50), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1335gat));
  NAND2_X1  g544(.A1(new_n719_), .A2(new_n655_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT111), .ZN(new_n747_));
  AOI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n610_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n667_), .A2(new_n668_), .A3(new_n718_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n610_), .A2(G85gat), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT112), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n748_), .B1(new_n750_), .B2(new_n752_), .ZN(G1336gat));
  INV_X1    g552(.A(G92gat), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n749_), .A2(new_n754_), .A3(new_n727_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n747_), .A2(new_n620_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(new_n754_), .ZN(G1337gat));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n746_), .B(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(new_n388_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT113), .B1(new_n760_), .B2(new_n452_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G99gat), .B1(new_n749_), .B2(new_n388_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT51), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n765_), .A3(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1338gat));
  NAND3_X1  g566(.A1(new_n747_), .A2(new_n334_), .A3(new_n435_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n667_), .A2(new_n435_), .A3(new_n668_), .A4(new_n718_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G106gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G106gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n588_), .A2(new_n589_), .A3(new_n550_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n775_), .B(KEYINPUT54), .C1(new_n606_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n584_), .A2(new_n586_), .A3(new_n549_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n659_), .A3(new_n603_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n775_), .B1(new_n780_), .B2(KEYINPUT54), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(KEYINPUT54), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n778_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n541_), .A2(new_n539_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n538_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n546_), .B(new_n784_), .C1(new_n785_), .C2(new_n539_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n547_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n562_), .A2(new_n788_), .A3(KEYINPUT55), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n555_), .B1(new_n564_), .B2(new_n559_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n566_), .A2(new_n567_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n571_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT116), .B1(new_n561_), .B2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n789_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n561_), .A2(new_n794_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT115), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n561_), .A2(new_n799_), .A3(new_n794_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n578_), .B1(new_n796_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n787_), .B1(new_n802_), .B2(KEYINPUT56), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n803_), .B(new_n580_), .C1(KEYINPUT56), .C2(new_n802_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT58), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n660_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n790_), .A2(KEYINPUT55), .A3(new_n557_), .A4(new_n558_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n808_), .A2(KEYINPUT116), .B1(new_n792_), .B2(new_n571_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n809_), .A2(new_n789_), .A3(new_n798_), .A4(new_n800_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT117), .B1(new_n810_), .B2(new_n578_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n580_), .B1(new_n811_), .B2(KEYINPUT56), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n802_), .A2(new_n813_), .A3(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n549_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n807_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n802_), .A2(new_n813_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n581_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n550_), .B1(new_n811_), .B2(KEYINPUT56), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(KEYINPUT118), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n547_), .B(new_n786_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n816_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n504_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n824_), .B1(new_n823_), .B2(new_n504_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n806_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n783_), .B1(new_n828_), .B2(new_n535_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n610_), .A2(new_n345_), .A3(new_n696_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT59), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  OR3_X1    g630(.A1(new_n778_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n823_), .A2(new_n504_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT57), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n834_), .A2(new_n825_), .B1(new_n660_), .B2(new_n805_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n832_), .B1(new_n835_), .B2(new_n603_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  INV_X1    g636(.A(new_n830_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n831_), .A2(new_n839_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n840_), .A2(new_n371_), .A3(new_n550_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT119), .B1(new_n829_), .B2(new_n830_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n832_), .B1(new_n835_), .B2(new_n536_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n838_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n842_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(G113gat), .B1(new_n846_), .B2(new_n549_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n841_), .A2(new_n847_), .ZN(G1340gat));
  NOR2_X1   g647(.A1(new_n716_), .A2(new_n717_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n372_), .B1(new_n850_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n846_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n372_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G120gat), .B1(new_n840_), .B2(new_n850_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1341gat));
  NOR3_X1   g653(.A1(new_n840_), .A2(new_n366_), .A3(new_n535_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n829_), .A2(KEYINPUT119), .A3(new_n830_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n844_), .B1(new_n843_), .B2(new_n838_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n603_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n366_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n668_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT120), .B1(new_n861_), .B2(G127gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n855_), .B1(new_n860_), .B2(new_n862_), .ZN(G1342gat));
  NOR3_X1   g662(.A1(new_n840_), .A2(new_n367_), .A3(new_n659_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n504_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n367_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n504_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT121), .B1(new_n869_), .B2(G134gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n864_), .B1(new_n868_), .B2(new_n870_), .ZN(G1343gat));
  NOR2_X1   g670(.A1(new_n829_), .A2(new_n442_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n696_), .A2(new_n344_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n680_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n550_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT122), .B(G141gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1344gat));
  NAND3_X1  g678(.A1(new_n872_), .A2(new_n849_), .A3(new_n875_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g680(.A1(new_n876_), .A2(new_n668_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT61), .B(G155gat), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT123), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n882_), .B(new_n884_), .ZN(G1346gat));
  INV_X1    g684(.A(G162gat), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n876_), .A2(new_n886_), .A3(new_n659_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n872_), .A2(new_n865_), .A3(new_n875_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n886_), .B2(new_n888_), .ZN(G1347gat));
  INV_X1    g688(.A(KEYINPUT22), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n680_), .A2(new_n344_), .A3(new_n418_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n836_), .A2(new_n890_), .A3(new_n549_), .A4(new_n892_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(G169gat), .ZN(new_n896_));
  INV_X1    g695(.A(new_n836_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n897_), .A2(new_n550_), .A3(new_n891_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n894_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n215_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n896_), .B1(new_n900_), .B2(new_n895_), .ZN(G1348gat));
  NOR2_X1   g700(.A1(new_n897_), .A2(new_n891_), .ZN(new_n902_));
  AOI21_X1  g701(.A(G176gat), .B1(new_n902_), .B2(new_n849_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n829_), .A2(new_n891_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n850_), .A2(new_n216_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(G1349gat));
  AOI21_X1  g705(.A(G183gat), .B1(new_n904_), .B2(new_n603_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n535_), .A2(new_n245_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n902_), .B2(new_n908_), .ZN(G1350gat));
  NAND3_X1  g708(.A1(new_n902_), .A2(new_n865_), .A3(new_n246_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n897_), .A2(new_n659_), .A3(new_n891_), .ZN(new_n911_));
  INV_X1    g710(.A(G190gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(G1351gat));
  NOR2_X1   g712(.A1(new_n874_), .A2(new_n610_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n914_), .A2(KEYINPUT125), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n843_), .A2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n727_), .B1(KEYINPUT125), .B2(new_n914_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n916_), .A2(new_n549_), .A3(new_n917_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g718(.A1(new_n916_), .A2(new_n849_), .A3(new_n917_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g720(.A(KEYINPUT63), .B(G211gat), .ZN(new_n922_));
  OR2_X1    g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n916_), .A2(new_n536_), .A3(new_n917_), .ZN(new_n924_));
  MUX2_X1   g723(.A(new_n922_), .B(new_n923_), .S(new_n924_), .Z(G1354gat));
  NAND2_X1  g724(.A1(new_n660_), .A2(G218gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT126), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n843_), .A2(new_n917_), .A3(new_n915_), .A4(new_n927_), .ZN(new_n928_));
  AND4_X1   g727(.A1(new_n865_), .A2(new_n843_), .A3(new_n917_), .A4(new_n915_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(G218gat), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(KEYINPUT127), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n932_), .B(new_n928_), .C1(new_n929_), .C2(G218gat), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n933_), .ZN(G1355gat));
endmodule


