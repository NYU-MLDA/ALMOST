//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n966_, new_n967_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1001_, new_n1002_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1024_, new_n1025_,
    new_n1026_, new_n1028_, new_n1029_, new_n1031_, new_n1032_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT103), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT19), .ZN(new_n205_));
  AND3_X1   g004(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT22), .B(G169gat), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(new_n211_), .A3(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT26), .B(G190gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT25), .B(G183gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n211_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n213_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n218_), .A2(new_n208_), .A3(new_n221_), .A4(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n215_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G197gat), .ZN(new_n227_));
  INV_X1    g026(.A(G204gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G197gat), .A2(G204gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT21), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT91), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n229_), .A2(KEYINPUT21), .A3(new_n230_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n234_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n238_), .A2(KEYINPUT21), .A3(new_n229_), .A4(new_n230_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT20), .B1(new_n226_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G183gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT25), .B1(new_n242_), .B2(KEYINPUT79), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT79), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(G183gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n216_), .A2(new_n243_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT80), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n216_), .A2(KEYINPUT80), .A3(new_n243_), .A4(new_n246_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G183gat), .A2(G190gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT23), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n224_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n211_), .A2(KEYINPUT24), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(new_n219_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n249_), .A2(new_n250_), .A3(new_n258_), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n208_), .A2(new_n209_), .B1(G169gat), .B2(G176gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT81), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n223_), .A2(KEYINPUT22), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT22), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(G169gat), .ZN(new_n265_));
  AND4_X1   g064(.A1(new_n261_), .A2(new_n263_), .A3(new_n265_), .A4(new_n213_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n260_), .B1(new_n262_), .B2(new_n266_), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n259_), .A2(new_n267_), .B1(new_n239_), .B2(new_n237_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n205_), .B1(new_n241_), .B2(new_n268_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n237_), .A2(new_n239_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(new_n267_), .A3(new_n259_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT20), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n226_), .B2(new_n240_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n269_), .B1(new_n205_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT32), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G8gat), .B(G36gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n277_), .B(KEYINPUT96), .Z(new_n278_));
  XOR2_X1   g077(.A(G64gat), .B(G92gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n278_), .A2(new_n279_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n278_), .A2(new_n279_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n281_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n276_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n275_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT101), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT101), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n275_), .A2(new_n287_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n274_), .A2(new_n205_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n260_), .A2(new_n214_), .B1(new_n258_), .B2(new_n218_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n272_), .B1(new_n270_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n259_), .A2(new_n267_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n240_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n205_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n292_), .A2(new_n298_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n289_), .B(new_n291_), .C1(new_n299_), .C2(new_n287_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G1gat), .B(G29gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT0), .ZN(new_n302_));
  INV_X1    g101(.A(G57gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(G85gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT4), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310_));
  OR2_X1    g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT88), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT87), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT87), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT88), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n311_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n311_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n310_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G141gat), .A2(G148gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT2), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT3), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT3), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(G141gat), .B2(G148gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n321_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n310_), .A2(KEYINPUT1), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT1), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(G155gat), .A3(G162gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n314_), .A2(KEYINPUT88), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n312_), .A2(KEYINPUT87), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n331_), .B1(new_n335_), .B2(new_n316_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n320_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n337_), .A2(new_n322_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  OAI22_X1  g138(.A1(new_n319_), .A2(new_n327_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G134gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G127gat), .ZN(new_n342_));
  INV_X1    g141(.A(G127gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G134gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT84), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n342_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n345_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n347_));
  OAI21_X1  g146(.A(G113gat), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n343_), .A2(G134gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n341_), .A2(G127gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT84), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G113gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n342_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n348_), .A2(G120gat), .A3(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(G120gat), .B1(new_n348_), .B2(new_n354_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n340_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G120gat), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n346_), .A2(new_n347_), .A3(G113gat), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n352_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n348_), .A2(new_n354_), .A3(G120gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n331_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n338_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n335_), .A2(new_n316_), .B1(G155gat), .B2(G162gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n321_), .A2(new_n326_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n361_), .A2(new_n362_), .A3(new_n365_), .A4(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT98), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n357_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n355_), .A2(new_n356_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n364_), .A2(new_n338_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(KEYINPUT98), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n309_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT99), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n357_), .B2(KEYINPUT4), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n361_), .A2(new_n362_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n378_), .A2(KEYINPUT99), .A3(new_n309_), .A4(new_n340_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n308_), .B1(new_n375_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n371_), .A2(new_n374_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n307_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n306_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n381_), .A2(new_n306_), .A3(new_n384_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n300_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT100), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n389_), .B(new_n306_), .C1(new_n383_), .C2(new_n307_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n382_), .A2(KEYINPUT4), .ZN(new_n391_));
  INV_X1    g190(.A(new_n380_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n307_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n307_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n306_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT100), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n390_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n241_), .A2(new_n268_), .A3(new_n205_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n297_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n283_), .A2(new_n286_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT97), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n283_), .A2(new_n286_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT97), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n299_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(new_n401_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n402_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n397_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n381_), .A2(new_n384_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT33), .B1(new_n409_), .B2(new_n395_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n385_), .A2(KEYINPUT33), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n388_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G43gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(G15gat), .ZN(new_n418_));
  INV_X1    g217(.A(G15gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(G43gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT82), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n416_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G71gat), .B(G99gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n419_), .A2(G43gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n417_), .A2(G15gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT82), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n415_), .A3(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n424_), .A2(new_n425_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n425_), .B1(new_n424_), .B2(new_n430_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n414_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n295_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n425_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n422_), .A2(new_n423_), .A3(new_n416_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n415_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n424_), .A2(new_n430_), .A3(new_n425_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(KEYINPUT83), .A3(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n259_), .A2(new_n267_), .A3(KEYINPUT30), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n433_), .A2(new_n435_), .A3(new_n441_), .A4(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT83), .B1(new_n439_), .B2(new_n440_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n442_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT30), .B1(new_n259_), .B2(new_n267_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n444_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT85), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n443_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT86), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT31), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n443_), .A2(new_n447_), .A3(new_n448_), .A4(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n450_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n451_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n378_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n450_), .A2(new_n453_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT31), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n450_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n372_), .A3(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n456_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT89), .B1(new_n373_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n340_), .A2(new_n464_), .A3(KEYINPUT29), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(G233gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT90), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(G228gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(G228gat), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n467_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n270_), .A2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n474_));
  NAND2_X1  g273(.A1(new_n340_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n240_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n466_), .A2(new_n473_), .B1(new_n472_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G78gat), .B(G106gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  AOI211_X1 g279(.A(KEYINPUT89), .B(new_n462_), .C1(new_n365_), .C2(new_n368_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n464_), .B1(new_n340_), .B2(KEYINPUT29), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n473_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n476_), .A2(new_n472_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n480_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G22gat), .B(G50gat), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT28), .B1(new_n373_), .B2(new_n462_), .ZN(new_n490_));
  AND4_X1   g289(.A1(KEYINPUT28), .A2(new_n365_), .A3(new_n368_), .A4(new_n462_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n489_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n373_), .A2(KEYINPUT28), .A3(new_n462_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT28), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(new_n340_), .B2(KEYINPUT29), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n495_), .A3(new_n488_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT93), .ZN(new_n498_));
  AOI211_X1 g297(.A(KEYINPUT94), .B(new_n497_), .C1(new_n498_), .C2(new_n485_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT94), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n485_), .A2(new_n498_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n497_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n487_), .B1(new_n499_), .B2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT93), .B1(new_n477_), .B2(new_n479_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT94), .B1(new_n505_), .B2(new_n497_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n480_), .A2(new_n486_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n501_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n461_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n413_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n387_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n513_), .A2(new_n385_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n402_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT27), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n403_), .A2(new_n275_), .A3(KEYINPUT102), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT102), .B1(new_n403_), .B2(new_n275_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT27), .B(new_n406_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n514_), .A2(new_n517_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n456_), .A2(new_n460_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n510_), .A2(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n504_), .A2(new_n509_), .A3(new_n456_), .A4(new_n460_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n521_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n512_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT37), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT6), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT7), .ZN(new_n531_));
  INV_X1    g330(.A(G99gat), .ZN(new_n532_));
  INV_X1    g331(.A(G106gat), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n536_));
  AND4_X1   g335(.A1(new_n530_), .A2(new_n534_), .A3(new_n535_), .A4(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT65), .ZN(new_n538_));
  AND2_X1   g337(.A1(G85gat), .A2(G92gat), .ZN(new_n539_));
  NOR2_X1   g338(.A1(G85gat), .A2(G92gat), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(G92gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n305_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G85gat), .A2(G92gat), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(KEYINPUT65), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT8), .B1(new_n537_), .B2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n534_), .A2(new_n530_), .A3(new_n535_), .A4(new_n536_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT8), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n541_), .A4(new_n545_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT66), .ZN(new_n552_));
  OR2_X1    g351(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n533_), .A3(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n543_), .A2(KEYINPUT9), .A3(new_n544_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT9), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(G85gat), .A3(G92gat), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n530_), .A2(new_n559_), .A3(new_n535_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT64), .B1(new_n557_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n560_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT64), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n562_), .A2(new_n563_), .A3(new_n555_), .A4(new_n556_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n551_), .A2(new_n552_), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n552_), .B1(new_n551_), .B2(new_n565_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G29gat), .B(G36gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G43gat), .B(G50gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT34), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n571_), .B(KEYINPUT15), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n551_), .A2(new_n565_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n576_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n578_), .A2(new_n579_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n572_), .A2(new_n577_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT74), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(new_n579_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT72), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT72), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n578_), .A2(new_n579_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n571_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n566_), .A2(new_n567_), .A3(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n574_), .B(new_n580_), .C1(new_n588_), .C2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT74), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n572_), .A2(new_n581_), .A3(new_n592_), .A4(new_n577_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n583_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(new_n341_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT73), .ZN(new_n597_));
  INV_X1    g396(.A(G162gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n599_), .A2(new_n600_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n594_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n594_), .B2(new_n602_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n527_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n583_), .A2(new_n591_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n606_), .A2(new_n600_), .A3(new_n599_), .A4(new_n593_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n594_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(KEYINPUT37), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT75), .B(G15gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(G22gat), .ZN(new_n612_));
  INV_X1    g411(.A(G1gat), .ZN(new_n613_));
  INV_X1    g412(.A(G8gat), .ZN(new_n614_));
  OAI21_X1  g413(.A(KEYINPUT14), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(G1gat), .B(G8gat), .Z(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n612_), .A2(new_n617_), .A3(new_n615_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G57gat), .B(G64gat), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT11), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT67), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT67), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n627_), .A3(KEYINPUT11), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n624_), .A2(KEYINPUT11), .ZN(new_n630_));
  XOR2_X1   g429(.A(G71gat), .B(G78gat), .Z(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n626_), .A2(new_n630_), .A3(new_n631_), .A4(new_n628_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n623_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n623_), .A2(new_n636_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G127gat), .B(G155gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT16), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(new_n242_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(G211gat), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT17), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n643_), .A2(new_n644_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n639_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT76), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n637_), .B(new_n638_), .C1(new_n644_), .C2(new_n643_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n648_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n526_), .A2(new_n610_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT13), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT70), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n579_), .A2(new_n635_), .A3(KEYINPUT12), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n635_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT12), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n658_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(G230gat), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n467_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n568_), .B2(new_n636_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n579_), .A2(KEYINPUT66), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n551_), .A2(new_n565_), .A3(new_n552_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n666_), .A3(new_n636_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n659_), .A2(new_n667_), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n661_), .A2(new_n664_), .B1(new_n668_), .B2(new_n663_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(G120gat), .B(G148gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(new_n228_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(KEYINPUT5), .B(G176gat), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n671_), .B(new_n672_), .Z(new_n673_));
  NAND2_X1  g472(.A1(new_n669_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n566_), .A2(new_n567_), .A3(new_n635_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n636_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n663_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n657_), .B1(new_n677_), .B2(KEYINPUT12), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n667_), .B1(new_n662_), .B2(new_n467_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT68), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT68), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n669_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n673_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n675_), .B1(new_n686_), .B2(KEYINPUT69), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT69), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n682_), .A2(new_n684_), .A3(new_n688_), .A4(new_n685_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n656_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n685_), .B1(new_n669_), .B2(new_n683_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n661_), .A2(new_n664_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n692_), .A2(new_n683_), .A3(new_n678_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT69), .B1(new_n691_), .B2(new_n693_), .ZN(new_n694_));
  AND4_X1   g493(.A1(new_n656_), .A2(new_n694_), .A3(new_n689_), .A4(new_n674_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n655_), .B1(new_n690_), .B2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n694_), .A2(new_n689_), .A3(new_n674_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT70), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n694_), .A2(new_n656_), .A3(new_n689_), .A4(new_n674_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(KEYINPUT13), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n621_), .A2(new_n589_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT77), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n619_), .A2(new_n620_), .A3(new_n571_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n701_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n621_), .A2(KEYINPUT77), .A3(new_n589_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n704_), .A2(G229gat), .A3(G233gat), .A4(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n621_), .A2(new_n578_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(G229gat), .A2(G233gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n703_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(G169gat), .B(G197gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(G141gat), .ZN(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT78), .B(G113gat), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n712_), .B(new_n713_), .Z(new_n714_));
  NAND2_X1  g513(.A1(new_n710_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n714_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n706_), .A2(new_n709_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n696_), .A2(new_n700_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n654_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n514_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n721_), .A2(new_n613_), .A3(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n202_), .A2(KEYINPUT103), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n203_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n603_), .A2(new_n604_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n652_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n650_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n521_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n524_), .ZN(new_n732_));
  AOI22_X1  g531(.A1(new_n509_), .A2(new_n504_), .B1(new_n456_), .B2(new_n460_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n397_), .B(new_n407_), .C1(new_n385_), .C2(KEYINPUT33), .ZN(new_n735_));
  INV_X1    g534(.A(new_n412_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n461_), .B(new_n510_), .C1(new_n737_), .C2(new_n388_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n730_), .B1(new_n734_), .B2(new_n738_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n739_), .A2(new_n696_), .A3(new_n700_), .A4(new_n718_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G1gat), .B1(new_n740_), .B2(new_n514_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n725_), .B(new_n741_), .C1(new_n203_), .C2(new_n723_), .ZN(G1324gat));
  INV_X1    g541(.A(KEYINPUT40), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n517_), .A2(new_n520_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n653_), .A2(new_n726_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n512_), .B2(new_n525_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n719_), .A2(new_n745_), .A3(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT39), .B1(new_n748_), .B2(new_n614_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT104), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(KEYINPUT39), .C1(new_n748_), .C2(new_n614_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT39), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n753_), .B(G8gat), .C1(new_n740_), .C2(new_n745_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT105), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n720_), .A2(new_n744_), .A3(new_n739_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n753_), .A4(G8gat), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n750_), .A2(new_n752_), .A3(new_n755_), .A4(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n721_), .A2(new_n614_), .A3(new_n744_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n759_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n743_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n759_), .A2(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT106), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n759_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(KEYINPUT40), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n764_), .A2(new_n768_), .ZN(G1325gat));
  OAI21_X1  g568(.A(G15gat), .B1(new_n740_), .B2(new_n461_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT41), .Z(new_n771_));
  NAND3_X1  g570(.A1(new_n721_), .A2(new_n419_), .A3(new_n522_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1326gat));
  OAI21_X1  g572(.A(G22gat), .B1(new_n740_), .B2(new_n510_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT42), .ZN(new_n775_));
  INV_X1    g574(.A(G22gat), .ZN(new_n776_));
  INV_X1    g575(.A(new_n510_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n721_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n775_), .A2(new_n778_), .ZN(G1327gat));
  INV_X1    g578(.A(G29gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n610_), .B1(new_n512_), .B2(new_n525_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n729_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT43), .B(new_n610_), .C1(new_n512_), .C2(new_n525_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(new_n720_), .A3(new_n784_), .ZN(new_n785_));
  XOR2_X1   g584(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n783_), .A2(new_n720_), .A3(KEYINPUT44), .A4(new_n784_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n722_), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n780_), .B1(new_n789_), .B2(KEYINPUT108), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(KEYINPUT108), .B2(new_n789_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n526_), .A2(new_n727_), .A3(new_n729_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n720_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(new_n780_), .A3(new_n722_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n791_), .A2(new_n795_), .ZN(G1328gat));
  AOI21_X1  g595(.A(new_n745_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n788_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(G36gat), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n745_), .A2(G36gat), .ZN(new_n801_));
  XOR2_X1   g600(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n802_));
  NAND3_X1  g601(.A1(new_n794_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n802_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n801_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n793_), .B2(new_n805_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n799_), .A2(new_n800_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(G36gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n797_), .B2(new_n788_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n803_), .A2(new_n806_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT110), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n808_), .A2(new_n812_), .A3(KEYINPUT46), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT46), .B1(new_n808_), .B2(new_n812_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1329gat));
  NAND4_X1  g614(.A1(new_n787_), .A2(G43gat), .A3(new_n522_), .A4(new_n788_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n417_), .B1(new_n793_), .B2(new_n461_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g618(.A(G50gat), .B1(new_n794_), .B2(new_n777_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n787_), .A2(G50gat), .A3(new_n777_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(new_n788_), .ZN(G1331gat));
  AOI21_X1  g621(.A(new_n718_), .B1(new_n696_), .B2(new_n700_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n654_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(new_n303_), .A3(new_n722_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n739_), .ZN(new_n826_));
  OAI21_X1  g625(.A(G57gat), .B1(new_n826_), .B2(new_n514_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1332gat));
  OAI21_X1  g627(.A(G64gat), .B1(new_n826_), .B2(new_n745_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT48), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n745_), .A2(G64gat), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT111), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n824_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(G1333gat));
  INV_X1    g633(.A(G71gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n824_), .A2(new_n835_), .A3(new_n522_), .ZN(new_n836_));
  OAI21_X1  g635(.A(G71gat), .B1(new_n826_), .B2(new_n461_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n837_), .A2(new_n838_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n836_), .B1(new_n839_), .B2(new_n840_), .ZN(G1334gat));
  OAI21_X1  g640(.A(G78gat), .B1(new_n826_), .B2(new_n510_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT50), .ZN(new_n843_));
  INV_X1    g642(.A(G78gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n824_), .A2(new_n844_), .A3(new_n777_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1335gat));
  NAND2_X1  g645(.A1(new_n792_), .A2(new_n823_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(new_n305_), .A3(new_n722_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n783_), .A2(new_n784_), .A3(new_n823_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G85gat), .B1(new_n850_), .B2(new_n514_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1336gat));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n848_), .A2(new_n744_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n542_), .ZN(new_n855_));
  AOI211_X1 g654(.A(KEYINPUT113), .B(G92gat), .C1(new_n848_), .C2(new_n744_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n744_), .A2(G92gat), .ZN(new_n857_));
  OAI22_X1  g656(.A1(new_n855_), .A2(new_n856_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n858_));
  XOR2_X1   g657(.A(new_n858_), .B(KEYINPUT114), .Z(G1337gat));
  OAI21_X1  g658(.A(G99gat), .B1(new_n850_), .B2(new_n461_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n522_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n847_), .B2(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g662(.A1(new_n783_), .A2(new_n777_), .A3(new_n784_), .A4(new_n823_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n864_), .A2(new_n865_), .A3(G106gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n864_), .B2(G106gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n510_), .A2(G106gat), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI22_X1  g668(.A1(new_n866_), .A2(new_n867_), .B1(new_n847_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT115), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n872_));
  OAI221_X1 g671(.A(new_n872_), .B1(new_n847_), .B2(new_n869_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n871_), .A2(KEYINPUT53), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT53), .B1(new_n871_), .B2(new_n873_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1339gat));
  NOR3_X1   g675(.A1(new_n610_), .A2(new_n718_), .A3(new_n653_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n696_), .A3(new_n700_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n703_), .A2(G229gat), .A3(G233gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n716_), .B1(new_n881_), .B2(new_n707_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n704_), .A2(new_n705_), .A3(new_n708_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n717_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n690_), .B2(new_n695_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n667_), .B(new_n657_), .C1(new_n677_), .C2(KEYINPUT12), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n661_), .A2(KEYINPUT117), .A3(new_n667_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n890_), .A2(new_n891_), .A3(new_n663_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT55), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n692_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n661_), .A2(KEYINPUT55), .A3(new_n664_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n685_), .B1(new_n892_), .B2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT56), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n679_), .A2(new_n680_), .A3(new_n893_), .ZN(new_n900_));
  AOI21_X1  g699(.A(KEYINPUT55), .B1(new_n661_), .B2(new_n664_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n890_), .A2(new_n891_), .A3(new_n663_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n904_), .A2(KEYINPUT56), .A3(new_n685_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n899_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n718_), .A2(new_n674_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT116), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n718_), .A2(KEYINPUT116), .A3(new_n674_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n906_), .A2(new_n909_), .A3(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n726_), .B1(new_n887_), .B2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT118), .B1(new_n912_), .B2(KEYINPUT57), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n675_), .A2(new_n885_), .ZN(new_n914_));
  AOI21_X1  g713(.A(KEYINPUT56), .B1(new_n904_), .B2(new_n685_), .ZN(new_n915_));
  AOI211_X1 g714(.A(new_n898_), .B(new_n673_), .C1(new_n902_), .C2(new_n903_), .ZN(new_n916_));
  OAI211_X1 g715(.A(KEYINPUT58), .B(new_n914_), .C1(new_n915_), .C2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n610_), .ZN(new_n918_));
  AOI21_X1  g717(.A(KEYINPUT58), .B1(new_n906_), .B2(new_n914_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n920_), .B1(new_n912_), .B2(KEYINPUT57), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n885_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n909_), .A2(new_n910_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n899_), .B2(new_n905_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n727_), .B1(new_n922_), .B2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT118), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT57), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n925_), .A2(new_n926_), .A3(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n913_), .A2(new_n921_), .A3(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n880_), .B1(new_n929_), .B2(new_n653_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n514_), .A2(new_n744_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n733_), .A2(new_n931_), .ZN(new_n932_));
  OAI21_X1  g731(.A(KEYINPUT59), .B1(new_n930_), .B2(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n912_), .A2(KEYINPUT57), .ZN(new_n934_));
  OAI211_X1 g733(.A(KEYINPUT57), .B(new_n727_), .C1(new_n922_), .C2(new_n924_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n906_), .A2(new_n914_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT58), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n938_), .A2(new_n610_), .A3(new_n917_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n935_), .A2(new_n939_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n653_), .B1(new_n934_), .B2(new_n940_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n878_), .B(KEYINPUT54), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n944_));
  INV_X1    g743(.A(new_n932_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n943_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n933_), .A2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n718_), .ZN(new_n948_));
  OAI21_X1  g747(.A(G113gat), .B1(new_n947_), .B2(new_n948_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n930_), .A2(new_n932_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n950_), .A2(new_n352_), .A3(new_n718_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n949_), .A2(new_n951_), .ZN(G1340gat));
  AND3_X1   g751(.A1(new_n925_), .A2(new_n926_), .A3(new_n927_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n926_), .B1(new_n925_), .B2(new_n927_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n953_), .A2(new_n954_), .A3(new_n940_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n942_), .B1(new_n955_), .B2(new_n729_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n696_), .A2(new_n700_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n957_), .B1(new_n959_), .B2(G120gat), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n956_), .A2(new_n945_), .A3(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(new_n958_), .ZN(new_n962_));
  OAI21_X1  g761(.A(G120gat), .B1(new_n962_), .B2(new_n947_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n950_), .A2(new_n957_), .A3(new_n960_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n963_), .A2(new_n964_), .ZN(G1341gat));
  OAI21_X1  g764(.A(G127gat), .B1(new_n947_), .B2(new_n653_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n950_), .A2(new_n343_), .A3(new_n729_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(new_n967_), .ZN(G1342gat));
  INV_X1    g767(.A(new_n610_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(KEYINPUT119), .B(G134gat), .ZN(new_n970_));
  NOR3_X1   g769(.A1(new_n947_), .A2(new_n969_), .A3(new_n970_), .ZN(new_n971_));
  AOI21_X1  g770(.A(G134gat), .B1(new_n950_), .B2(new_n726_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(new_n971_), .A2(new_n972_), .ZN(G1343gat));
  XNOR2_X1  g772(.A(KEYINPUT121), .B(G141gat), .ZN(new_n974_));
  INV_X1    g773(.A(new_n974_), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT120), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n732_), .A2(new_n931_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n976_), .B1(new_n930_), .B2(new_n977_), .ZN(new_n978_));
  INV_X1    g777(.A(new_n977_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(new_n954_), .A2(new_n940_), .ZN(new_n980_));
  AOI21_X1  g779(.A(new_n729_), .B1(new_n980_), .B2(new_n928_), .ZN(new_n981_));
  OAI211_X1 g780(.A(KEYINPUT120), .B(new_n979_), .C1(new_n981_), .C2(new_n880_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n978_), .A2(new_n982_), .ZN(new_n983_));
  AOI21_X1  g782(.A(new_n975_), .B1(new_n983_), .B2(new_n718_), .ZN(new_n984_));
  AOI211_X1 g783(.A(new_n948_), .B(new_n974_), .C1(new_n978_), .C2(new_n982_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n984_), .A2(new_n985_), .ZN(G1344gat));
  AOI21_X1  g785(.A(KEYINPUT120), .B1(new_n956_), .B2(new_n979_), .ZN(new_n987_));
  NOR3_X1   g786(.A1(new_n930_), .A2(new_n976_), .A3(new_n977_), .ZN(new_n988_));
  OAI21_X1  g787(.A(new_n958_), .B1(new_n987_), .B2(new_n988_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n989_), .A2(G148gat), .ZN(new_n990_));
  INV_X1    g789(.A(G148gat), .ZN(new_n991_));
  NAND3_X1  g790(.A1(new_n983_), .A2(new_n991_), .A3(new_n958_), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n990_), .A2(new_n992_), .ZN(G1345gat));
  OAI21_X1  g792(.A(new_n729_), .B1(new_n987_), .B2(new_n988_), .ZN(new_n994_));
  XNOR2_X1  g793(.A(KEYINPUT61), .B(G155gat), .ZN(new_n995_));
  XNOR2_X1  g794(.A(new_n995_), .B(KEYINPUT122), .ZN(new_n996_));
  INV_X1    g795(.A(new_n996_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n994_), .A2(new_n997_), .ZN(new_n998_));
  NAND3_X1  g797(.A1(new_n983_), .A2(new_n729_), .A3(new_n996_), .ZN(new_n999_));
  NAND2_X1  g798(.A1(new_n998_), .A2(new_n999_), .ZN(G1346gat));
  NAND3_X1  g799(.A1(new_n983_), .A2(new_n598_), .A3(new_n726_), .ZN(new_n1001_));
  AOI21_X1  g800(.A(new_n969_), .B1(new_n978_), .B2(new_n982_), .ZN(new_n1002_));
  OAI21_X1  g801(.A(new_n1001_), .B1(new_n598_), .B2(new_n1002_), .ZN(G1347gat));
  NOR2_X1   g802(.A1(new_n722_), .A2(new_n745_), .ZN(new_n1004_));
  NAND2_X1  g803(.A1(new_n1004_), .A2(new_n522_), .ZN(new_n1005_));
  XNOR2_X1  g804(.A(new_n1005_), .B(KEYINPUT123), .ZN(new_n1006_));
  NOR2_X1   g805(.A1(new_n1006_), .A2(new_n777_), .ZN(new_n1007_));
  NAND2_X1  g806(.A1(new_n943_), .A2(new_n1007_), .ZN(new_n1008_));
  INV_X1    g807(.A(new_n1008_), .ZN(new_n1009_));
  NAND2_X1  g808(.A1(new_n1009_), .A2(new_n718_), .ZN(new_n1010_));
  NAND2_X1  g809(.A1(new_n1010_), .A2(G169gat), .ZN(new_n1011_));
  INV_X1    g810(.A(KEYINPUT62), .ZN(new_n1012_));
  NAND2_X1  g811(.A1(new_n1011_), .A2(new_n1012_), .ZN(new_n1013_));
  NAND3_X1  g812(.A1(new_n1010_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n1014_));
  NAND3_X1  g813(.A1(new_n1009_), .A2(new_n718_), .A3(new_n212_), .ZN(new_n1015_));
  NAND3_X1  g814(.A1(new_n1013_), .A2(new_n1014_), .A3(new_n1015_), .ZN(G1348gat));
  AOI21_X1  g815(.A(G176gat), .B1(new_n1009_), .B2(new_n958_), .ZN(new_n1017_));
  INV_X1    g816(.A(KEYINPUT124), .ZN(new_n1018_));
  AOI21_X1  g817(.A(new_n1018_), .B1(new_n956_), .B2(new_n510_), .ZN(new_n1019_));
  NOR3_X1   g818(.A1(new_n930_), .A2(KEYINPUT124), .A3(new_n777_), .ZN(new_n1020_));
  OR2_X1    g819(.A1(new_n1019_), .A2(new_n1020_), .ZN(new_n1021_));
  NOR3_X1   g820(.A1(new_n959_), .A2(new_n1006_), .A3(new_n213_), .ZN(new_n1022_));
  AOI21_X1  g821(.A(new_n1017_), .B1(new_n1021_), .B2(new_n1022_), .ZN(G1349gat));
  NOR3_X1   g822(.A1(new_n1008_), .A2(new_n653_), .A3(new_n217_), .ZN(new_n1024_));
  NOR2_X1   g823(.A1(new_n1006_), .A2(new_n653_), .ZN(new_n1025_));
  OAI21_X1  g824(.A(new_n1025_), .B1(new_n1019_), .B2(new_n1020_), .ZN(new_n1026_));
  AOI21_X1  g825(.A(new_n1024_), .B1(new_n1026_), .B2(new_n242_), .ZN(G1350gat));
  OAI21_X1  g826(.A(G190gat), .B1(new_n1008_), .B2(new_n969_), .ZN(new_n1028_));
  NAND2_X1  g827(.A1(new_n726_), .A2(new_n216_), .ZN(new_n1029_));
  OAI21_X1  g828(.A(new_n1028_), .B1(new_n1008_), .B2(new_n1029_), .ZN(G1351gat));
  INV_X1    g829(.A(KEYINPUT125), .ZN(new_n1031_));
  NAND2_X1  g830(.A1(new_n732_), .A2(new_n1004_), .ZN(new_n1032_));
  INV_X1    g831(.A(new_n1032_), .ZN(new_n1033_));
  AOI21_X1  g832(.A(new_n1031_), .B1(new_n956_), .B2(new_n1033_), .ZN(new_n1034_));
  NOR3_X1   g833(.A1(new_n930_), .A2(KEYINPUT125), .A3(new_n1032_), .ZN(new_n1035_));
  OAI21_X1  g834(.A(new_n718_), .B1(new_n1034_), .B2(new_n1035_), .ZN(new_n1036_));
  NAND2_X1  g835(.A1(new_n1036_), .A2(G197gat), .ZN(new_n1037_));
  OAI21_X1  g836(.A(KEYINPUT125), .B1(new_n930_), .B2(new_n1032_), .ZN(new_n1038_));
  OAI211_X1 g837(.A(new_n1031_), .B(new_n1033_), .C1(new_n981_), .C2(new_n880_), .ZN(new_n1039_));
  NAND2_X1  g838(.A1(new_n1038_), .A2(new_n1039_), .ZN(new_n1040_));
  NAND3_X1  g839(.A1(new_n1040_), .A2(new_n227_), .A3(new_n718_), .ZN(new_n1041_));
  NAND2_X1  g840(.A1(new_n1037_), .A2(new_n1041_), .ZN(G1352gat));
  AOI21_X1  g841(.A(new_n959_), .B1(new_n1038_), .B2(new_n1039_), .ZN(new_n1043_));
  XOR2_X1   g842(.A(KEYINPUT126), .B(G204gat), .Z(new_n1044_));
  NAND2_X1  g843(.A1(new_n1043_), .A2(new_n1044_), .ZN(new_n1045_));
  AND2_X1   g844(.A1(new_n228_), .A2(KEYINPUT126), .ZN(new_n1046_));
  OAI21_X1  g845(.A(new_n1045_), .B1(new_n1043_), .B2(new_n1046_), .ZN(G1353gat));
  NOR2_X1   g846(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1048_));
  INV_X1    g847(.A(new_n1048_), .ZN(new_n1049_));
  AOI21_X1  g848(.A(new_n653_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1050_));
  AOI21_X1  g849(.A(new_n1049_), .B1(new_n1040_), .B2(new_n1050_), .ZN(new_n1051_));
  INV_X1    g850(.A(new_n1050_), .ZN(new_n1052_));
  AOI211_X1 g851(.A(new_n1048_), .B(new_n1052_), .C1(new_n1038_), .C2(new_n1039_), .ZN(new_n1053_));
  NOR2_X1   g852(.A1(new_n1051_), .A2(new_n1053_), .ZN(G1354gat));
  NAND2_X1  g853(.A1(new_n1040_), .A2(new_n726_), .ZN(new_n1055_));
  INV_X1    g854(.A(G218gat), .ZN(new_n1056_));
  NAND2_X1  g855(.A1(new_n610_), .A2(G218gat), .ZN(new_n1057_));
  XOR2_X1   g856(.A(new_n1057_), .B(KEYINPUT127), .Z(new_n1058_));
  AOI22_X1  g857(.A1(new_n1055_), .A2(new_n1056_), .B1(new_n1040_), .B2(new_n1058_), .ZN(G1355gat));
endmodule


