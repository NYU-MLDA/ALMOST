//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202_));
  XOR2_X1   g001(.A(G85gat), .B(G92gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT6), .ZN(new_n205_));
  NAND2_X1  g004(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n203_), .B1(new_n207_), .B2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT8), .ZN(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT10), .B(G99gat), .Z(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n216_));
  INV_X1    g015(.A(G85gat), .ZN(new_n217_));
  INV_X1    g016(.A(G92gat), .ZN(new_n218_));
  OR3_X1    g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT9), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n215_), .A2(new_n216_), .A3(new_n219_), .A4(new_n205_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n212_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(G71gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(G78gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G57gat), .B(G64gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT11), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n224_), .A2(KEYINPUT11), .ZN(new_n227_));
  OR3_X1    g026(.A1(new_n223_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(new_n226_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n221_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G230gat), .ZN(new_n232_));
  INV_X1    g031(.A(G233gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n202_), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  AOI211_X1 g035(.A(KEYINPUT68), .B(new_n234_), .C1(new_n221_), .C2(new_n230_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n212_), .A2(new_n220_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n230_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT12), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n239_), .B(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(KEYINPUT12), .A3(new_n240_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n238_), .A2(new_n243_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(KEYINPUT66), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(new_n231_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n234_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G120gat), .B(G148gat), .ZN(new_n252_));
  INV_X1    g051(.A(G204gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT5), .ZN(new_n255_));
  INV_X1    g054(.A(G176gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n251_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n247_), .A2(new_n250_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n257_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT13), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT13), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n258_), .A2(new_n264_), .A3(new_n261_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT76), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G29gat), .B(G36gat), .ZN(new_n268_));
  INV_X1    g067(.A(G43gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G50gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT15), .ZN(new_n273_));
  XOR2_X1   g072(.A(G15gat), .B(G22gat), .Z(new_n274_));
  NAND2_X1  g073(.A1(G1gat), .A2(G8gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n274_), .B1(KEYINPUT14), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT72), .ZN(new_n277_));
  XOR2_X1   g076(.A(G1gat), .B(G8gat), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n276_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n273_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n279_), .A2(new_n283_), .A3(new_n272_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G229gat), .A2(G233gat), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n267_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n286_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n284_), .B2(new_n273_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n292_), .A2(KEYINPUT76), .A3(new_n288_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n272_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n284_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(new_n286_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n284_), .A2(KEYINPUT75), .A3(new_n294_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n289_), .A3(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n290_), .A2(new_n293_), .A3(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G169gat), .B(G197gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(G141gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT77), .ZN(new_n303_));
  INV_X1    g102(.A(G113gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n300_), .A2(new_n305_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n266_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT26), .B(G190gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT78), .ZN(new_n312_));
  INV_X1    g111(.A(G183gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n312_), .B1(new_n313_), .B2(KEYINPUT25), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT25), .B(G183gat), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n311_), .B(new_n314_), .C1(new_n315_), .C2(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT23), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT79), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT23), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(G183gat), .A3(G190gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT79), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n317_), .A2(new_n322_), .A3(KEYINPUT23), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n319_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT24), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(G169gat), .B2(G176gat), .ZN(new_n326_));
  INV_X1    g125(.A(G169gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n256_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n325_), .A2(new_n327_), .A3(new_n256_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n316_), .A2(new_n324_), .A3(new_n329_), .A4(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n318_), .A2(new_n321_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n332_), .B1(G183gat), .B2(G190gat), .ZN(new_n333_));
  OR2_X1    g132(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(G176gat), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n333_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n331_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT30), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n342_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G71gat), .B(G99gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G15gat), .B(G43gat), .Z(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n343_), .A2(new_n344_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n344_), .A2(new_n349_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(G113gat), .ZN(new_n355_));
  INV_X1    g154(.A(G127gat), .ZN(new_n356_));
  INV_X1    g155(.A(G134gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G127gat), .A2(G134gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(new_n304_), .A3(new_n359_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n355_), .A2(G120gat), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(G120gat), .B1(new_n355_), .B2(new_n360_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT31), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n353_), .A2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n351_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n353_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT1), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(G155gat), .B2(G162gat), .ZN(new_n371_));
  NOR2_X1   g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n369_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(G155gat), .A3(G162gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n372_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT1), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n377_), .A3(KEYINPUT82), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n373_), .A2(new_n374_), .A3(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(G141gat), .B(G148gat), .Z(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G141gat), .A2(G148gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT2), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n382_), .B1(new_n383_), .B2(KEYINPUT83), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(KEYINPUT83), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n387_));
  OR3_X1    g186(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(KEYINPUT83), .A3(new_n383_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .A4(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n390_), .A2(new_n376_), .A3(new_n375_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n381_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n394_));
  XOR2_X1   g193(.A(new_n393_), .B(new_n394_), .Z(new_n395_));
  XNOR2_X1  g194(.A(G22gat), .B(G50gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n395_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT89), .B(G78gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(new_n214_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n392_), .B1(new_n381_), .B2(new_n391_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n253_), .A2(G197gat), .ZN(new_n402_));
  INV_X1    g201(.A(G197gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(G204gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n404_), .A3(KEYINPUT85), .ZN(new_n405_));
  OR3_X1    g204(.A1(new_n253_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(KEYINPUT21), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT21), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n403_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT86), .B1(new_n403_), .B2(G204gat), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n408_), .B(new_n402_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G211gat), .B(G218gat), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n407_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n402_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(KEYINPUT21), .A3(new_n412_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n414_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n415_), .B1(new_n414_), .B2(new_n417_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n401_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G228gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(new_n233_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT88), .B1(new_n420_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n381_), .A2(new_n391_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT29), .ZN(new_n426_));
  INV_X1    g225(.A(new_n419_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n414_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n422_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n424_), .A2(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n414_), .A2(new_n417_), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n401_), .A2(new_n422_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n400_), .B1(new_n432_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n400_), .ZN(new_n437_));
  AOI211_X1 g236(.A(new_n437_), .B(new_n434_), .C1(new_n424_), .C2(new_n431_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n398_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n420_), .A2(KEYINPUT88), .A3(new_n423_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n430_), .B1(new_n429_), .B2(new_n422_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n435_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n437_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n432_), .A2(new_n400_), .A3(new_n435_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n395_), .B(new_n396_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n439_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n368_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT27), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G64gat), .B(G92gat), .ZN(new_n450_));
  INV_X1    g249(.A(G36gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT93), .B(G8gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n452_), .A2(new_n453_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n452_), .A2(new_n453_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n455_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT19), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n324_), .B1(G183gat), .B2(G190gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT91), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n338_), .B1(new_n336_), .B2(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n465_), .B(new_n467_), .C1(new_n466_), .C2(new_n338_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n311_), .A2(new_n315_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n329_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n469_), .A2(KEYINPUT90), .A3(new_n329_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n472_), .A2(new_n332_), .A3(new_n473_), .A4(new_n330_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n433_), .B1(new_n468_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n414_), .A2(new_n417_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT20), .B1(new_n340_), .B2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n464_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(new_n468_), .A3(new_n433_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n340_), .B2(new_n476_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n464_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n479_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n462_), .A2(new_n478_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n462_), .B1(new_n478_), .B2(new_n483_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n449_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n468_), .B(new_n474_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n482_), .B1(new_n488_), .B2(new_n481_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n475_), .A2(new_n464_), .A3(new_n477_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n461_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(KEYINPUT27), .A3(new_n484_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n362_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n355_), .A2(G120gat), .A3(new_n360_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n425_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n363_), .A2(new_n381_), .A3(new_n391_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(KEYINPUT4), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G225gat), .A2(G233gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT4), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n425_), .A2(new_n501_), .A3(new_n495_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n496_), .A2(new_n499_), .A3(new_n497_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT0), .B(G57gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(G85gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(G1gat), .B(G29gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT96), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n508_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AOI211_X1 g312(.A(new_n510_), .B(new_n508_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n487_), .B(new_n492_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n448_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT97), .ZN(new_n517_));
  NOR2_X1   g316(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n509_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n518_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n503_), .A2(new_n504_), .A3(new_n508_), .A4(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n478_), .A2(new_n483_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n461_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n498_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n508_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n496_), .A2(new_n500_), .A3(new_n497_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n524_), .A2(new_n484_), .A3(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n522_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n513_), .A2(new_n514_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT32), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n461_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n478_), .B(new_n483_), .C1(new_n461_), .C2(new_n532_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT95), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT95), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n533_), .B(new_n537_), .C1(new_n490_), .C2(new_n489_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n530_), .B1(new_n531_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n439_), .A2(new_n446_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n517_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n514_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n512_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(new_n510_), .A3(new_n509_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n539_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n522_), .A2(new_n529_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(KEYINPUT97), .A3(new_n447_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT98), .B1(new_n447_), .B2(new_n515_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n531_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n487_), .A2(new_n492_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT98), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n551_), .A2(new_n541_), .A3(new_n553_), .A4(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n542_), .A2(new_n549_), .A3(new_n550_), .A4(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n368_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n516_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n245_), .A2(new_n273_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT34), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(KEYINPUT69), .B(KEYINPUT35), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n221_), .A2(new_n272_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n559_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n562_), .A2(new_n564_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n559_), .A2(new_n570_), .A3(new_n565_), .A4(new_n566_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G190gat), .B(G218gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G134gat), .ZN(new_n574_));
  INV_X1    g373(.A(G162gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT36), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT70), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT71), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n572_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n569_), .A2(new_n582_), .A3(new_n576_), .A4(new_n571_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT37), .ZN(new_n585_));
  INV_X1    g384(.A(new_n579_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n572_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n583_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n585_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n230_), .B(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(new_n284_), .Z(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT16), .B(G183gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(G211gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT73), .B(KEYINPUT17), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n593_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT74), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n597_), .B(KEYINPUT17), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n593_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n590_), .A2(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n310_), .A2(new_n558_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(G1gat), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(new_n607_), .A3(new_n531_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT38), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n266_), .A2(KEYINPUT99), .A3(new_n309_), .A4(new_n604_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n587_), .A2(new_n583_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n556_), .A2(new_n557_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n516_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n610_), .A2(new_n611_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n310_), .B2(new_n603_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n615_), .A2(KEYINPUT100), .A3(new_n617_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n551_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n609_), .B1(new_n622_), .B2(new_n607_), .ZN(G1324gat));
  OAI21_X1  g422(.A(G8gat), .B1(new_n618_), .B2(new_n553_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  OAI211_X1 g425(.A(KEYINPUT39), .B(G8gat), .C1(new_n618_), .C2(new_n553_), .ZN(new_n627_));
  INV_X1    g426(.A(G8gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n606_), .A2(new_n628_), .A3(new_n552_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT101), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(new_n627_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT102), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n626_), .A2(new_n630_), .A3(new_n633_), .A4(new_n627_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g435(.A(G15gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n606_), .A2(new_n637_), .A3(new_n368_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n557_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n639_), .A2(KEYINPUT103), .A3(new_n637_), .ZN(new_n640_));
  OAI21_X1  g439(.A(KEYINPUT103), .B1(new_n639_), .B2(new_n637_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n640_), .A2(new_n641_), .A3(KEYINPUT41), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(new_n640_), .B2(new_n641_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n638_), .B1(new_n642_), .B2(new_n643_), .ZN(G1326gat));
  INV_X1    g443(.A(G22gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n620_), .A2(new_n621_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n646_), .B2(new_n541_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT42), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n606_), .A2(new_n645_), .A3(new_n541_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1327gat));
  NOR4_X1   g449(.A1(new_n310_), .A2(new_n604_), .A3(new_n558_), .A4(new_n611_), .ZN(new_n651_));
  INV_X1    g450(.A(G29gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(new_n652_), .A3(new_n531_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n266_), .A2(new_n309_), .A3(new_n603_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  INV_X1    g456(.A(new_n590_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n614_), .B2(new_n658_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n558_), .A2(KEYINPUT43), .A3(new_n590_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n656_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n654_), .B1(new_n661_), .B2(KEYINPUT105), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT105), .B1(new_n661_), .B2(KEYINPUT104), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n614_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT43), .B1(new_n558_), .B2(new_n590_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n655_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n665_), .B(KEYINPUT44), .C1(new_n668_), .C2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n664_), .A2(new_n531_), .A3(new_n670_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n671_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT106), .B1(new_n671_), .B2(G29gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n653_), .B1(new_n672_), .B2(new_n673_), .ZN(G1328gat));
  NAND3_X1  g473(.A1(new_n651_), .A2(new_n451_), .A3(new_n552_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT45), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n552_), .B(new_n670_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n677_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT107), .B1(new_n677_), .B2(G36gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n676_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT46), .B(new_n676_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1329gat));
  OAI211_X1 g483(.A(new_n368_), .B(new_n670_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G43gat), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n651_), .A2(new_n269_), .A3(new_n368_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT108), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n686_), .A2(new_n691_), .A3(new_n688_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT47), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n691_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n694_));
  AOI211_X1 g493(.A(KEYINPUT108), .B(new_n687_), .C1(new_n685_), .C2(G43gat), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n694_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n693_), .A2(new_n697_), .ZN(G1330gat));
  NAND3_X1  g497(.A1(new_n651_), .A2(new_n271_), .A3(new_n541_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n664_), .A2(new_n541_), .A3(new_n670_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(new_n271_), .ZN(G1331gat));
  INV_X1    g500(.A(new_n266_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n558_), .A2(new_n309_), .ZN(new_n703_));
  AND4_X1   g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n604_), .A4(new_n611_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(G57gat), .A3(new_n531_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(KEYINPUT109), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n708_), .B1(new_n558_), .B2(new_n309_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n266_), .B1(new_n707_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n605_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n531_), .ZN(new_n713_));
  INV_X1    g512(.A(G57gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n706_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  AOI211_X1 g514(.A(KEYINPUT110), .B(G57gat), .C1(new_n712_), .C2(new_n531_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n705_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT111), .Z(G1332gat));
  INV_X1    g517(.A(G64gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n704_), .B2(new_n552_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT48), .Z(new_n721_));
  NAND3_X1  g520(.A1(new_n712_), .A2(new_n719_), .A3(new_n552_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1333gat));
  INV_X1    g522(.A(G71gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n704_), .B2(new_n368_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT49), .Z(new_n726_));
  NAND3_X1  g525(.A1(new_n712_), .A2(new_n724_), .A3(new_n368_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1334gat));
  INV_X1    g527(.A(G78gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n704_), .B2(new_n541_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT112), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT50), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n712_), .A2(new_n729_), .A3(new_n541_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1335gat));
  NAND2_X1  g533(.A1(new_n666_), .A2(new_n667_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n604_), .A2(new_n309_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n702_), .A3(new_n736_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n737_), .A2(new_n217_), .A3(new_n551_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n604_), .A2(new_n611_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n710_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT113), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n710_), .A2(KEYINPUT113), .A3(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n531_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n738_), .B1(new_n745_), .B2(new_n217_), .ZN(G1336gat));
  NOR3_X1   g545(.A1(new_n737_), .A2(new_n218_), .A3(new_n553_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n744_), .A2(new_n552_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n218_), .ZN(G1337gat));
  NAND3_X1  g548(.A1(new_n744_), .A2(new_n213_), .A3(new_n368_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G99gat), .B1(new_n737_), .B2(new_n557_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g552(.A1(new_n735_), .A2(new_n702_), .A3(new_n541_), .A4(new_n736_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(KEYINPUT115), .A3(G106gat), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(KEYINPUT52), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT115), .B1(new_n754_), .B2(G106gat), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n756_), .B(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n743_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT113), .B1(new_n710_), .B2(new_n739_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n214_), .B(new_n541_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n744_), .A2(KEYINPUT114), .A3(new_n214_), .A4(new_n541_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n758_), .A2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n758_), .A2(new_n765_), .A3(new_n767_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1339gat));
  NAND2_X1  g570(.A1(new_n258_), .A2(new_n309_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n246_), .A2(new_n243_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n231_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n234_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n236_), .A2(new_n237_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n238_), .A2(KEYINPUT55), .A3(new_n243_), .A4(new_n246_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT56), .B1(new_n780_), .B2(new_n260_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(KEYINPUT56), .A3(new_n260_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n772_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT119), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n297_), .A2(new_n288_), .A3(new_n298_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n305_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n292_), .A2(new_n289_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n786_), .A2(KEYINPUT118), .A3(new_n305_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n789_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n785_), .B1(new_n792_), .B2(new_n306_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n307_), .A2(KEYINPUT119), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n796_), .A2(new_n262_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n611_), .B1(new_n784_), .B2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n783_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n796_), .B(new_n258_), .C1(new_n801_), .C2(new_n781_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n782_), .A2(new_n783_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n805_), .A2(KEYINPUT58), .A3(new_n258_), .A4(new_n796_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(new_n806_), .A3(new_n658_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n309_), .B(new_n258_), .C1(new_n801_), .C2(new_n781_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n796_), .A2(new_n262_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n799_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n611_), .A3(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n800_), .A2(new_n807_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n603_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n815_));
  INV_X1    g614(.A(new_n309_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n266_), .A2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n815_), .B1(new_n817_), .B2(new_n605_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n815_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n711_), .A2(new_n816_), .A3(new_n266_), .A4(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n814_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n448_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n551_), .A2(new_n552_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT121), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n823_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n823_), .A2(KEYINPUT59), .A3(new_n827_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n830_), .A2(KEYINPUT122), .A3(new_n831_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n834_), .A2(G113gat), .A3(new_n309_), .A4(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n304_), .B1(new_n828_), .B2(new_n816_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1340gat));
  INV_X1    g637(.A(new_n828_), .ZN(new_n839_));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n266_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n839_), .B(new_n841_), .C1(KEYINPUT60), .C2(new_n840_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n266_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n840_), .ZN(G1341gat));
  NAND4_X1  g643(.A1(new_n834_), .A2(G127gat), .A3(new_n604_), .A4(new_n835_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n356_), .B1(new_n828_), .B2(new_n603_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1342gat));
  NAND4_X1  g646(.A1(new_n834_), .A2(G134gat), .A3(new_n658_), .A4(new_n835_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n357_), .B1(new_n828_), .B2(new_n611_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1343gat));
  AOI21_X1  g649(.A(new_n821_), .B1(new_n813_), .B2(new_n603_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n368_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n852_), .A2(new_n825_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n541_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n816_), .ZN(new_n855_));
  INV_X1    g654(.A(G141gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1344gat));
  NOR2_X1   g656(.A1(new_n854_), .A2(new_n266_), .ZN(new_n858_));
  INV_X1    g657(.A(G148gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1345gat));
  NOR2_X1   g659(.A1(new_n854_), .A2(new_n603_), .ZN(new_n861_));
  XOR2_X1   g660(.A(KEYINPUT61), .B(G155gat), .Z(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1346gat));
  AND2_X1   g662(.A1(new_n853_), .A2(new_n541_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n611_), .ZN(new_n865_));
  AOI21_X1  g664(.A(G162gat), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n590_), .A2(new_n575_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT123), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n864_), .B2(new_n868_), .ZN(G1347gat));
  NOR2_X1   g668(.A1(new_n553_), .A2(new_n531_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n811_), .B1(new_n810_), .B2(new_n611_), .ZN(new_n871_));
  AOI211_X1 g670(.A(new_n865_), .B(new_n799_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n604_), .B1(new_n873_), .B2(new_n807_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n824_), .B(new_n870_), .C1(new_n874_), .C2(new_n821_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT124), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n448_), .B1(new_n814_), .B2(new_n822_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(new_n878_), .A3(new_n870_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n334_), .A2(new_n335_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n309_), .A3(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(G169gat), .B1(new_n875_), .B2(new_n816_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n883_), .A2(KEYINPUT62), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(KEYINPUT62), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n882_), .B1(new_n884_), .B2(new_n885_), .ZN(G1348gat));
  NAND3_X1  g685(.A1(new_n880_), .A2(new_n256_), .A3(new_n702_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G176gat), .B1(new_n875_), .B2(new_n266_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1349gat));
  INV_X1    g688(.A(new_n315_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n878_), .B1(new_n877_), .B2(new_n870_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n870_), .ZN(new_n892_));
  NOR4_X1   g691(.A1(new_n851_), .A2(KEYINPUT124), .A3(new_n448_), .A4(new_n892_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n604_), .B(new_n890_), .C1(new_n891_), .C2(new_n893_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n894_), .A2(KEYINPUT125), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(KEYINPUT125), .ZN(new_n896_));
  INV_X1    g695(.A(new_n875_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G183gat), .B1(new_n897_), .B2(new_n604_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n895_), .A2(new_n896_), .A3(new_n898_), .ZN(G1350gat));
  OAI211_X1 g698(.A(new_n865_), .B(new_n311_), .C1(new_n891_), .C2(new_n893_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n590_), .B1(new_n876_), .B2(new_n879_), .ZN(new_n901_));
  INV_X1    g700(.A(G190gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT126), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n900_), .B(KEYINPUT126), .C1(new_n901_), .C2(new_n902_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1351gat));
  NAND3_X1  g706(.A1(new_n852_), .A2(new_n541_), .A3(new_n870_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT127), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n852_), .A2(new_n910_), .A3(new_n541_), .A4(new_n870_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n816_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n403_), .ZN(G1352gat));
  AOI21_X1  g712(.A(new_n266_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n253_), .ZN(G1353gat));
  XNOR2_X1  g714(.A(KEYINPUT63), .B(G211gat), .ZN(new_n916_));
  AOI211_X1 g715(.A(new_n603_), .B(new_n916_), .C1(new_n909_), .C2(new_n911_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n909_), .A2(new_n911_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n604_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n917_), .B1(new_n919_), .B2(new_n920_), .ZN(G1354gat));
  NAND2_X1  g720(.A1(new_n918_), .A2(new_n865_), .ZN(new_n922_));
  INV_X1    g721(.A(G218gat), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n924_));
  AOI22_X1  g723(.A1(new_n922_), .A2(new_n923_), .B1(new_n924_), .B2(new_n658_), .ZN(G1355gat));
endmodule


