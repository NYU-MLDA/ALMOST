//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT71), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G57gat), .B(G64gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT68), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G71gat), .B(G78gat), .Z(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n210_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n211_));
  INV_X1    g010(.A(G64gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G57gat), .ZN(new_n213_));
  INV_X1    g012(.A(G57gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G64gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(new_n205_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n204_), .A2(KEYINPUT67), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT11), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n208_), .A2(new_n211_), .A3(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n209_), .B1(new_n219_), .B2(KEYINPUT11), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n220_), .B1(new_n219_), .B2(KEYINPUT11), .ZN(new_n224_));
  AOI211_X1 g023(.A(KEYINPUT68), .B(new_n207_), .C1(new_n217_), .C2(new_n218_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n223_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G99gat), .A2(G106gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT6), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT6), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(G99gat), .A3(G106gat), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G99gat), .A2(G106gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  OAI22_X1  g036(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n229_), .B1(new_n234_), .B2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(KEYINPUT10), .B(G99gat), .Z(new_n243_));
  INV_X1    g042(.A(G106gat), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n243_), .A2(new_n244_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n228_), .B1(new_n227_), .B2(KEYINPUT9), .ZN(new_n246_));
  NOR3_X1   g045(.A1(new_n227_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G85gat), .A2(G92gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT9), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n246_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n245_), .A2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT66), .B(KEYINPUT8), .Z(new_n254_));
  OAI211_X1 g053(.A(new_n229_), .B(new_n254_), .C1(new_n234_), .C2(new_n239_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n242_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n222_), .A2(new_n226_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT12), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G230gat), .A2(G233gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT12), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n257_), .A2(new_n258_), .A3(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n256_), .B1(new_n222_), .B2(new_n226_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n260_), .A2(new_n261_), .A3(new_n263_), .A4(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n267_), .A3(new_n257_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n261_), .B1(new_n264_), .B2(KEYINPUT69), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G120gat), .B(G148gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT5), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G176gat), .B(G204gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n266_), .A2(new_n270_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n275_), .B1(new_n266_), .B2(new_n270_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n203_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n266_), .A2(new_n270_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n274_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n266_), .A2(new_n270_), .A3(new_n275_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(KEYINPUT71), .A3(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n278_), .A2(new_n282_), .A3(KEYINPUT13), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT13), .B1(new_n278_), .B2(new_n282_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n202_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n278_), .A2(new_n282_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT13), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n278_), .A2(new_n282_), .A3(KEYINPUT13), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(KEYINPUT72), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G229gat), .A2(G233gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G29gat), .B(G36gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G43gat), .B(G50gat), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G15gat), .B(G22gat), .ZN(new_n300_));
  INV_X1    g099(.A(G1gat), .ZN(new_n301_));
  INV_X1    g100(.A(G8gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT14), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT78), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT78), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n300_), .A2(new_n306_), .A3(new_n303_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT79), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G1gat), .B(G8gat), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n308_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(new_n307_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT79), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n311_), .B1(new_n316_), .B2(new_n309_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n299_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n312_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n316_), .A2(new_n311_), .A3(new_n309_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n298_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n318_), .A2(KEYINPUT82), .A3(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT82), .B1(new_n318_), .B2(new_n321_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n293_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n321_), .A2(new_n292_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT15), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n298_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n296_), .A2(KEYINPUT15), .A3(new_n297_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n324_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G113gat), .B(G141gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G169gat), .B(G197gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT84), .B1(new_n332_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT84), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n324_), .A2(new_n338_), .A3(new_n331_), .A4(new_n335_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n332_), .A2(KEYINPUT83), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT83), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n324_), .A2(new_n342_), .A3(new_n331_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n336_), .A3(new_n343_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n291_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G71gat), .B(G99gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(G43gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT30), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT25), .B(G183gat), .ZN(new_n350_));
  INV_X1    g149(.A(G190gat), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT26), .B1(new_n351_), .B2(KEYINPUT85), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n351_), .A2(KEYINPUT26), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n350_), .B(new_n352_), .C1(new_n353_), .C2(KEYINPUT85), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G183gat), .A2(G190gat), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(G169gat), .ZN(new_n362_));
  INV_X1    g161(.A(G176gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OR3_X1    g163(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n354_), .A2(new_n359_), .A3(new_n364_), .A4(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n357_), .B(new_n358_), .C1(G183gat), .C2(G190gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT22), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n367_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n349_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n349_), .A2(new_n372_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G227gat), .A2(G233gat), .ZN(new_n376_));
  INV_X1    g175(.A(G15gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n373_), .A2(new_n378_), .A3(new_n374_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT31), .ZN(new_n384_));
  INV_X1    g183(.A(G134gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G127gat), .ZN(new_n386_));
  INV_X1    g185(.A(G127gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G134gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G120gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G113gat), .ZN(new_n391_));
  INV_X1    g190(.A(G113gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G120gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n386_), .A2(new_n388_), .A3(new_n391_), .A4(new_n393_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT87), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n395_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n401_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n395_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n404_), .A3(new_n399_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT31), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n380_), .A2(new_n381_), .A3(new_n407_), .A4(new_n382_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n384_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n406_), .B1(new_n384_), .B2(new_n408_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(G85gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT0), .B(G57gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G225gat), .A2(G233gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418_));
  NOR2_X1   g217(.A1(G155gat), .A2(G162gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT89), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT89), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n421_), .B1(G155gat), .B2(G162gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G155gat), .A2(G162gat), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n420_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G141gat), .A2(G148gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT2), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n428_));
  INV_X1    g227(.A(G141gat), .ZN(new_n429_));
  INV_X1    g228(.A(G148gat), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n429_), .B(new_n430_), .C1(KEYINPUT90), .C2(KEYINPUT3), .ZN(new_n431_));
  NAND2_X1  g230(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n427_), .B(new_n428_), .C1(new_n431_), .C2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT91), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(KEYINPUT91), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n424_), .B1(new_n434_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n423_), .A2(KEYINPUT1), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT1), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(G155gat), .A3(G162gat), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n420_), .A2(new_n422_), .A3(new_n441_), .A4(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G141gat), .A2(G148gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n446_), .A2(new_n425_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n440_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT92), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT92), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n440_), .A2(new_n451_), .A3(new_n448_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n450_), .A2(new_n452_), .A3(new_n405_), .A4(new_n402_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n427_), .A2(new_n428_), .ZN(new_n454_));
  OR2_X1    g253(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(new_n432_), .A3(new_n445_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n454_), .A2(new_n456_), .A3(new_n437_), .A4(new_n438_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n457_), .A2(new_n424_), .B1(new_n444_), .B2(new_n447_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT100), .ZN(new_n459_));
  INV_X1    g258(.A(new_n396_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n459_), .B1(new_n404_), .B2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n395_), .A2(KEYINPUT100), .A3(new_n396_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n418_), .B1(new_n453_), .B2(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n440_), .A2(new_n451_), .A3(new_n448_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n451_), .B1(new_n440_), .B2(new_n448_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT4), .B1(new_n467_), .B2(new_n406_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n417_), .B1(new_n464_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n453_), .A2(new_n463_), .A3(new_n416_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT101), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT101), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n453_), .A2(new_n473_), .A3(new_n416_), .A4(new_n463_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n415_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n415_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n469_), .A2(new_n472_), .A3(new_n474_), .A4(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(G204gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(KEYINPUT95), .A3(G197gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(G197gat), .ZN(new_n483_));
  INV_X1    g282(.A(G197gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(G204gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(KEYINPUT21), .B(new_n482_), .C1(new_n486_), .C2(KEYINPUT95), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n483_), .A2(new_n485_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT21), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G211gat), .B(G218gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n487_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n488_), .A2(new_n489_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n491_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT29), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n496_), .B1(new_n458_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G233gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT94), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(G228gat), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(G228gat), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n499_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G78gat), .B(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n465_), .A2(new_n466_), .A3(new_n497_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n494_), .B1(new_n489_), .B2(new_n488_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n509_), .A2(new_n487_), .B1(new_n494_), .B2(new_n493_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n510_), .A2(new_n504_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n505_), .B(new_n507_), .C1(new_n508_), .C2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT96), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n497_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G22gat), .B(G50gat), .Z(new_n519_));
  OAI211_X1 g318(.A(new_n497_), .B(new_n516_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n519_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n514_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n505_), .B1(new_n508_), .B2(new_n511_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n506_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n512_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n519_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n450_), .A2(new_n452_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n516_), .B1(new_n529_), .B2(new_n497_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n520_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n528_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n534_), .A2(KEYINPUT96), .A3(new_n512_), .A4(new_n525_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n527_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT20), .ZN(new_n537_));
  INV_X1    g336(.A(new_n371_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT26), .B(G190gat), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n539_), .A2(KEYINPUT97), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(KEYINPUT97), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n350_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n364_), .A2(new_n359_), .A3(new_n365_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n538_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n537_), .B1(new_n544_), .B2(new_n510_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n372_), .A2(new_n496_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT98), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G226gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT19), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n372_), .A2(new_n496_), .A3(KEYINPUT98), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n545_), .A2(new_n548_), .A3(new_n551_), .A4(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G8gat), .B(G36gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G64gat), .B(G92gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n366_), .A2(new_n492_), .A3(new_n495_), .A4(new_n371_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n559_), .B(KEYINPUT20), .C1(new_n544_), .C2(new_n510_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n550_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n553_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n560_), .A2(new_n550_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n545_), .A2(new_n548_), .A3(new_n552_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n550_), .B2(new_n564_), .ZN(new_n565_));
  OAI211_X1 g364(.A(KEYINPUT27), .B(new_n562_), .C1(new_n565_), .C2(new_n558_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT27), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n553_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n558_), .B1(new_n553_), .B2(new_n561_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n411_), .A2(new_n480_), .A3(new_n536_), .A4(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n527_), .A2(new_n535_), .A3(new_n570_), .A4(new_n566_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(new_n479_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n558_), .A2(KEYINPUT32), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n553_), .A2(new_n561_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n575_), .B1(new_n576_), .B2(KEYINPUT104), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n564_), .A2(new_n550_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n563_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n578_), .A2(new_n579_), .A3(KEYINPUT32), .A4(new_n558_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n553_), .A2(KEYINPUT104), .A3(new_n561_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n577_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n472_), .A2(new_n474_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n477_), .B1(new_n583_), .B2(new_n469_), .ZN(new_n584_));
  AND4_X1   g383(.A1(new_n469_), .A2(new_n472_), .A3(new_n474_), .A4(new_n477_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n582_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT33), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n478_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n568_), .A2(new_n569_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n453_), .A2(new_n463_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n415_), .B1(new_n590_), .B2(new_n416_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT103), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n416_), .B1(new_n464_), .B2(new_n468_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT103), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n594_), .B(new_n415_), .C1(new_n590_), .C2(new_n416_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n592_), .A2(new_n593_), .A3(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(new_n589_), .A3(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n415_), .A2(new_n587_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n469_), .A2(new_n472_), .A3(new_n474_), .A4(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT102), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT102), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n583_), .A2(new_n601_), .A3(new_n469_), .A4(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n586_), .B1(new_n597_), .B2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n574_), .B1(new_n604_), .B2(new_n536_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n572_), .B1(new_n605_), .B2(new_n411_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n346_), .A2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(G127gat), .B(G155gat), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT16), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT17), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT80), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n615_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n319_), .A2(KEYINPUT80), .A3(new_n320_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n614_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n616_), .A2(new_n614_), .A3(new_n617_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n619_), .A2(new_n222_), .A3(new_n226_), .A4(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n222_), .A2(new_n226_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n620_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n622_), .B1(new_n623_), .B2(new_n618_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n613_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT81), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n611_), .A2(new_n612_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n621_), .A2(new_n624_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n625_), .A2(KEYINPUT81), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT34), .Z(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT73), .B(KEYINPUT35), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n242_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(new_n329_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n634_), .A2(new_n635_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT74), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n242_), .A2(new_n253_), .A3(new_n255_), .A4(new_n298_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n636_), .B1(new_n638_), .B2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n256_), .A2(new_n328_), .A3(new_n327_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n636_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n644_), .A2(new_n645_), .A3(new_n641_), .A4(new_n640_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(G190gat), .B(G218gat), .Z(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT75), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G134gat), .B(G162gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT36), .Z(new_n652_));
  NAND2_X1  g451(.A1(new_n647_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT76), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT37), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n651_), .A2(KEYINPUT36), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n643_), .A2(new_n646_), .A3(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n647_), .A2(new_n652_), .A3(KEYINPUT76), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n655_), .A2(new_n656_), .A3(new_n658_), .A4(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n653_), .A2(new_n658_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT37), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT77), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT77), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(new_n665_), .A3(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n632_), .A2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n607_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n301_), .A3(new_n479_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT38), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n655_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n411_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n536_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n596_), .A2(new_n589_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n677_), .A2(new_n588_), .A3(new_n600_), .A4(new_n602_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n676_), .B1(new_n678_), .B2(new_n586_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n679_), .B2(new_n574_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n674_), .B1(new_n680_), .B2(new_n572_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n346_), .A2(new_n631_), .A3(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G1gat), .B1(new_n682_), .B2(new_n480_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n670_), .A2(new_n671_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n672_), .A2(new_n683_), .A3(new_n684_), .ZN(G1324gat));
  INV_X1    g484(.A(new_n571_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n669_), .A2(new_n302_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT39), .ZN(new_n688_));
  INV_X1    g487(.A(new_n682_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n686_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n690_), .B2(G8gat), .ZN(new_n691_));
  AOI211_X1 g490(.A(KEYINPUT39), .B(new_n302_), .C1(new_n689_), .C2(new_n686_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n687_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g493(.A(G15gat), .B1(new_n682_), .B2(new_n675_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT41), .Z(new_n696_));
  NAND3_X1  g495(.A1(new_n669_), .A2(new_n377_), .A3(new_n411_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1326gat));
  OAI21_X1  g497(.A(G22gat), .B1(new_n682_), .B2(new_n536_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT42), .ZN(new_n700_));
  INV_X1    g499(.A(G22gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n669_), .A2(new_n701_), .A3(new_n676_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1327gat));
  NOR2_X1   g502(.A1(new_n631_), .A2(new_n673_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n607_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G29gat), .B1(new_n706_), .B2(new_n479_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n345_), .ZN(new_n708_));
  AND4_X1   g507(.A1(new_n632_), .A2(new_n285_), .A3(new_n290_), .A4(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n660_), .A2(new_n665_), .A3(new_n662_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n665_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n711_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT105), .B1(new_n664_), .B2(new_n666_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n710_), .B1(new_n606_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n667_), .A2(new_n710_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n680_), .B2(new_n572_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n709_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n720_), .A2(KEYINPUT106), .A3(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n709_), .B(KEYINPUT44), .C1(new_n717_), .C2(new_n719_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n479_), .A2(G29gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n707_), .B1(new_n728_), .B2(new_n729_), .ZN(G1328gat));
  NOR2_X1   g529(.A1(new_n571_), .A2(G36gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n607_), .A2(new_n704_), .A3(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n727_), .A2(new_n686_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n720_), .A2(KEYINPUT106), .A3(new_n721_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT106), .B1(new_n720_), .B2(new_n721_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n735_), .B(new_n736_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G36gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n736_), .B1(new_n726_), .B2(new_n735_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n734_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI211_X1 g543(.A(KEYINPUT46), .B(new_n734_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1329gat));
  INV_X1    g545(.A(G43gat), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n675_), .A2(new_n747_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n727_), .B(new_n748_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT109), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n726_), .A2(new_n751_), .A3(new_n727_), .A4(new_n748_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n747_), .B1(new_n705_), .B2(new_n675_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT47), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n750_), .A2(new_n752_), .A3(new_n756_), .A4(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1330gat));
  AOI21_X1  g557(.A(G50gat), .B1(new_n706_), .B2(new_n676_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n676_), .A2(G50gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n728_), .B2(new_n760_), .ZN(G1331gat));
  NAND4_X1  g560(.A1(new_n681_), .A2(new_n631_), .A3(new_n291_), .A4(new_n345_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n762_), .A2(new_n214_), .A3(new_n480_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n606_), .A2(new_n345_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT111), .Z(new_n766_));
  NAND2_X1  g565(.A1(new_n291_), .A2(new_n668_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT110), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n764_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n772_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(KEYINPUT113), .A3(new_n770_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n775_), .A3(new_n479_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n763_), .B1(new_n776_), .B2(new_n214_), .ZN(G1332gat));
  NOR2_X1   g576(.A1(new_n771_), .A2(new_n772_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n212_), .A3(new_n686_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G64gat), .B1(new_n762_), .B2(new_n571_), .ZN(new_n780_));
  XOR2_X1   g579(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(G1333gat));
  INV_X1    g582(.A(G71gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n778_), .A2(new_n784_), .A3(new_n411_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G71gat), .B1(new_n762_), .B2(new_n675_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT49), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1334gat));
  INV_X1    g587(.A(G78gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n778_), .A2(new_n789_), .A3(new_n676_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G78gat), .B1(new_n762_), .B2(new_n536_), .ZN(new_n791_));
  XOR2_X1   g590(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(G1335gat));
  OR2_X1    g593(.A1(new_n717_), .A2(new_n719_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n291_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n796_), .A2(new_n631_), .A3(new_n708_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(G85gat), .B1(new_n798_), .B2(new_n480_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n291_), .A2(new_n704_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n766_), .A2(new_n800_), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n480_), .A2(G85gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n799_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n803_), .B(KEYINPUT116), .Z(G1336gat));
  INV_X1    g603(.A(new_n801_), .ZN(new_n805_));
  AOI21_X1  g604(.A(G92gat), .B1(new_n805_), .B2(new_n686_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n798_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n686_), .A2(G92gat), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n808_), .B(KEYINPUT117), .Z(new_n809_));
  AOI21_X1  g608(.A(new_n806_), .B1(new_n807_), .B2(new_n809_), .ZN(G1337gat));
  OAI21_X1  g609(.A(G99gat), .B1(new_n798_), .B2(new_n675_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n411_), .A2(new_n243_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n801_), .B2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g613(.A1(new_n805_), .A2(new_n244_), .A3(new_n676_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n795_), .A2(new_n676_), .A3(new_n797_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n816_), .A2(new_n817_), .A3(G106gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n816_), .B2(G106gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n815_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g620(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n264_), .B1(new_n259_), .B2(KEYINPUT12), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n261_), .B1(new_n823_), .B2(new_n263_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n266_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n823_), .A2(KEYINPUT55), .A3(new_n261_), .A4(new_n263_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n275_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n321_), .A2(new_n293_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n336_), .B1(new_n831_), .B2(new_n330_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n322_), .A2(new_n323_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n292_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n830_), .A2(new_n835_), .A3(new_n281_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n828_), .A2(new_n829_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n822_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n828_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT56), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n276_), .B(new_n834_), .C1(new_n337_), .C2(new_n339_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n822_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n840_), .A2(new_n841_), .A3(new_n842_), .A4(new_n830_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n838_), .A2(new_n667_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n839_), .A2(new_n845_), .A3(KEYINPUT56), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n276_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n829_), .B1(new_n828_), .B2(KEYINPUT118), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n835_), .A2(new_n282_), .A3(new_n278_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n674_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n844_), .B1(new_n851_), .B2(KEYINPUT57), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n853_), .B(new_n674_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n632_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n711_), .A2(new_n712_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n631_), .A2(new_n345_), .A3(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n283_), .A2(new_n284_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n857_), .A2(new_n858_), .A3(KEYINPUT54), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n855_), .A2(new_n863_), .ZN(new_n864_));
  NOR4_X1   g663(.A1(new_n675_), .A2(new_n480_), .A3(new_n676_), .A4(new_n686_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT59), .ZN(new_n867_));
  OAI21_X1  g666(.A(G113gat), .B1(new_n867_), .B2(new_n345_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n866_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n869_), .A2(new_n392_), .A3(new_n708_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1340gat));
  OAI21_X1  g670(.A(G120gat), .B1(new_n867_), .B2(new_n796_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n390_), .B1(new_n796_), .B2(KEYINPUT60), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n869_), .B(new_n873_), .C1(KEYINPUT60), .C2(new_n390_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(G1341gat));
  OAI21_X1  g674(.A(G127gat), .B1(new_n867_), .B2(new_n632_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n869_), .A2(new_n387_), .A3(new_n631_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1342gat));
  OAI21_X1  g677(.A(G134gat), .B1(new_n867_), .B2(new_n856_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n869_), .A2(new_n385_), .A3(new_n674_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1343gat));
  NOR2_X1   g680(.A1(new_n861_), .A2(new_n862_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n849_), .A2(new_n850_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n673_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n853_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n851_), .A2(KEYINPUT57), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(new_n886_), .A3(new_n844_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n882_), .B1(new_n887_), .B2(new_n632_), .ZN(new_n888_));
  NOR4_X1   g687(.A1(new_n888_), .A2(new_n480_), .A3(new_n573_), .A4(new_n411_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n708_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n291_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT120), .B(G148gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1345gat));
  NAND2_X1  g693(.A1(new_n889_), .A2(new_n631_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1346gat));
  AOI21_X1  g696(.A(G162gat), .B1(new_n889_), .B2(new_n674_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n716_), .A2(G162gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(KEYINPUT121), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n898_), .B1(new_n889_), .B2(new_n900_), .ZN(G1347gat));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n902_));
  NOR4_X1   g701(.A1(new_n675_), .A2(new_n479_), .A3(new_n676_), .A4(new_n571_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n864_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n345_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n902_), .B1(new_n905_), .B2(new_n369_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(G169gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n362_), .B1(new_n905_), .B2(new_n902_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n906_), .B2(new_n908_), .ZN(G1348gat));
  NOR2_X1   g708(.A1(new_n904_), .A2(new_n796_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n363_), .A2(KEYINPUT122), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n363_), .A2(KEYINPUT122), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n913_), .B1(new_n910_), .B2(new_n912_), .ZN(G1349gat));
  NOR2_X1   g713(.A1(new_n904_), .A2(new_n632_), .ZN(new_n915_));
  MUX2_X1   g714(.A(G183gat), .B(new_n350_), .S(new_n915_), .Z(G1350gat));
  OR2_X1    g715(.A1(new_n540_), .A2(new_n541_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n864_), .A2(new_n674_), .A3(new_n917_), .A4(new_n903_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n904_), .A2(new_n856_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n351_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  OAI211_X1 g721(.A(KEYINPUT123), .B(new_n918_), .C1(new_n919_), .C2(new_n351_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1351gat));
  NOR3_X1   g723(.A1(new_n411_), .A2(new_n479_), .A3(new_n536_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n926_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n927_), .A2(new_n686_), .A3(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(KEYINPUT125), .B1(new_n864_), .B2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932_));
  AOI211_X1 g731(.A(new_n932_), .B(new_n929_), .C1(new_n855_), .C2(new_n863_), .ZN(new_n933_));
  OAI211_X1 g732(.A(G197gat), .B(new_n708_), .C1(new_n931_), .C2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(KEYINPUT126), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n931_), .A2(new_n933_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n484_), .B1(new_n936_), .B2(new_n345_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n932_), .B1(new_n888_), .B2(new_n929_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n864_), .A2(KEYINPUT125), .A3(new_n930_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n940_), .A2(new_n941_), .A3(G197gat), .A4(new_n708_), .ZN(new_n942_));
  AND3_X1   g741(.A1(new_n935_), .A2(new_n937_), .A3(new_n942_), .ZN(G1352gat));
  NAND2_X1  g742(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n940_), .A2(new_n291_), .A3(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n936_), .A2(new_n796_), .ZN(new_n946_));
  XOR2_X1   g745(.A(KEYINPUT127), .B(G204gat), .Z(new_n947_));
  OAI21_X1  g746(.A(new_n945_), .B1(new_n946_), .B2(new_n947_), .ZN(G1353gat));
  AOI211_X1 g747(.A(KEYINPUT63), .B(G211gat), .C1(new_n940_), .C2(new_n631_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(KEYINPUT63), .B(G211gat), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n936_), .A2(new_n632_), .A3(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n949_), .A2(new_n951_), .ZN(G1354gat));
  OAI21_X1  g751(.A(G218gat), .B1(new_n936_), .B2(new_n856_), .ZN(new_n953_));
  OR2_X1    g752(.A1(new_n673_), .A2(G218gat), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n936_), .B2(new_n954_), .ZN(G1355gat));
endmodule


