//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n959_, new_n960_,
    new_n961_, new_n963_, new_n964_, new_n965_, new_n967_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT81), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT82), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT23), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  OR3_X1    g014(.A1(new_n215_), .A2(KEYINPUT80), .A3(KEYINPUT26), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(KEYINPUT79), .A3(G183gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT26), .B1(new_n215_), .B2(KEYINPUT80), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n217_), .A2(G183gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(G183gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n214_), .B1(new_n220_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT83), .B(G176gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT22), .B(G169gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n203_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT84), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n231_), .B1(new_n232_), .B2(new_n208_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n229_), .A2(KEYINPUT84), .ZN(new_n237_));
  OAI22_X1  g036(.A1(new_n207_), .A2(new_n226_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G227gat), .A2(G233gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(G15gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n238_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G71gat), .B(G99gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT86), .B(G43gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n245_), .B(new_n246_), .Z(new_n247_));
  NOR2_X1   g046(.A1(new_n241_), .A2(new_n242_), .ZN(new_n248_));
  NOR3_X1   g047(.A1(new_n244_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT87), .ZN(new_n252_));
  XOR2_X1   g051(.A(G113gat), .B(G120gat), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT87), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n251_), .B(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(new_n253_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT88), .B1(new_n255_), .B2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT88), .B1(new_n257_), .B2(new_n253_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT31), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT89), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n247_), .B1(new_n244_), .B2(new_n248_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n250_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(KEYINPUT89), .ZN(new_n268_));
  INV_X1    g067(.A(new_n247_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n241_), .A2(new_n242_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(new_n243_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n268_), .B1(new_n249_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(G141gat), .A2(G148gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G155gat), .A2(G162gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT90), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT1), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n275_), .B(new_n276_), .C1(new_n279_), .C2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT2), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n284_), .B(new_n285_), .C1(new_n275_), .C2(KEYINPUT3), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n275_), .A2(KEYINPUT3), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT91), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT91), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n275_), .A2(new_n289_), .A3(KEYINPUT3), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n286_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n277_), .B(KEYINPUT90), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n280_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n282_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(KEYINPUT29), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT28), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G228gat), .A2(G233gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G211gat), .B(G218gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT95), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT93), .B(G197gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G204gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(G197gat), .B2(G204gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT21), .ZN(new_n304_));
  NOR3_X1   g103(.A1(new_n300_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G204gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n306_), .A2(G197gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n306_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n307_), .B1(new_n308_), .B2(KEYINPUT94), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT94), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n301_), .A2(new_n310_), .A3(new_n306_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n304_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n298_), .B(KEYINPUT95), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n314_), .B1(new_n304_), .B2(new_n303_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n305_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n297_), .B1(new_n316_), .B2(KEYINPUT92), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n296_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G106gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n303_), .A2(new_n304_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n300_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n303_), .A2(new_n304_), .ZN(new_n322_));
  OAI22_X1  g121(.A1(new_n321_), .A2(new_n312_), .B1(new_n322_), .B2(new_n300_), .ZN(new_n323_));
  INV_X1    g122(.A(G78gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n294_), .A2(KEYINPUT29), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n324_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n319_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(G106gat), .A3(new_n326_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G22gat), .B(G50gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n329_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n318_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(new_n331_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n332_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n318_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n329_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n336_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT18), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G64gat), .B(G92gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n238_), .A2(new_n323_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT26), .B(G190gat), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n217_), .A2(G183gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n349_), .A3(new_n223_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n204_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n202_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT97), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n214_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(KEYINPUT97), .A3(new_n352_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT98), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n228_), .B(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n227_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n203_), .B1(new_n234_), .B2(new_n233_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n357_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n316_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT19), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT20), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n347_), .A2(new_n365_), .A3(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n367_), .B(KEYINPUT96), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n205_), .B(KEYINPUT82), .ZN(new_n373_));
  INV_X1    g172(.A(new_n237_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n229_), .A2(KEYINPUT84), .B1(new_n234_), .B2(new_n233_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n373_), .A2(new_n225_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n316_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n368_), .B1(new_n323_), .B2(new_n363_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n372_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n346_), .B1(new_n370_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT20), .B1(new_n364_), .B2(new_n316_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n238_), .A2(new_n323_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n371_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n346_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n347_), .A2(new_n365_), .A3(new_n369_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n380_), .A2(new_n386_), .A3(KEYINPUT99), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT99), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n388_), .B(new_n346_), .C1(new_n370_), .C2(new_n379_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n259_), .A2(new_n294_), .A3(new_n261_), .ZN(new_n391_));
  OAI221_X1 g190(.A(new_n282_), .B1(new_n291_), .B2(new_n293_), .C1(new_n255_), .C2(new_n258_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(KEYINPUT4), .A3(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT100), .B(KEYINPUT4), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n259_), .A2(new_n294_), .A3(new_n261_), .A4(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n398_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT101), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G85gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT0), .B(G57gat), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n405_), .B(new_n406_), .Z(new_n407_));
  NAND4_X1  g206(.A1(new_n402_), .A2(new_n403_), .A3(KEYINPUT33), .A4(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n397_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n409_), .B2(new_n400_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT101), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n393_), .A2(new_n397_), .A3(new_n395_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n391_), .A2(new_n398_), .A3(new_n392_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n407_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n410_), .A2(new_n411_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n390_), .A2(new_n408_), .A3(new_n412_), .A4(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n384_), .A2(KEYINPUT32), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n370_), .A2(new_n379_), .A3(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(KEYINPUT102), .B(KEYINPUT20), .Z(new_n421_));
  NAND3_X1  g220(.A1(new_n347_), .A2(new_n365_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n367_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n377_), .A2(new_n378_), .A3(new_n372_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n420_), .B1(new_n425_), .B2(new_n419_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n399_), .A2(new_n401_), .A3(KEYINPUT103), .A4(new_n415_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n399_), .A2(new_n401_), .A3(new_n415_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT103), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(new_n410_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n426_), .A2(new_n427_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n342_), .B1(new_n418_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n427_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(new_n341_), .A3(new_n336_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n387_), .A2(new_n435_), .A3(new_n389_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n425_), .A2(new_n346_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(KEYINPUT27), .A3(new_n386_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n434_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n274_), .B1(new_n432_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(KEYINPUT104), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT104), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n436_), .A2(new_n443_), .A3(new_n438_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n342_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n433_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n267_), .B2(new_n272_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n441_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G190gat), .B(G218gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G134gat), .B(G162gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n453_), .B(KEYINPUT36), .Z(new_n454_));
  XOR2_X1   g253(.A(G85gat), .B(G92gat), .Z(new_n455_));
  INV_X1    g254(.A(KEYINPUT64), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(KEYINPUT9), .ZN(new_n457_));
  XOR2_X1   g256(.A(KEYINPUT10), .B(G99gat), .Z(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n319_), .ZN(new_n459_));
  INV_X1    g258(.A(G85gat), .ZN(new_n460_));
  INV_X1    g259(.A(G92gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT9), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G85gat), .B(G92gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(KEYINPUT64), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT6), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G99gat), .A3(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n457_), .A2(new_n459_), .A3(new_n464_), .A4(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT8), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT65), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT7), .ZN(new_n474_));
  INV_X1    g273(.A(G99gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n319_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n466_), .A2(new_n468_), .A3(KEYINPUT65), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n473_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n471_), .B1(new_n481_), .B2(new_n455_), .ZN(new_n482_));
  AOI211_X1 g281(.A(KEYINPUT8), .B(new_n463_), .C1(new_n479_), .C2(new_n469_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n470_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT15), .ZN(new_n485_));
  INV_X1    g284(.A(G50gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(G43gat), .ZN(new_n487_));
  INV_X1    g286(.A(G43gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(G50gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G29gat), .B(G36gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(G36gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(G29gat), .ZN(new_n494_));
  INV_X1    g293(.A(G29gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(G36gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G43gat), .B(G50gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n492_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n492_), .B2(new_n499_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n485_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n500_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n497_), .A2(new_n498_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n490_), .A2(new_n491_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n492_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(KEYINPUT15), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n484_), .A2(new_n510_), .A3(KEYINPUT68), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT68), .B1(new_n484_), .B2(new_n510_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT69), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT68), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n501_), .A2(new_n502_), .A3(new_n485_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT15), .B1(new_n507_), .B2(new_n508_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n470_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n466_), .A2(new_n468_), .A3(KEYINPUT65), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT65), .B1(new_n466_), .B2(new_n468_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n519_), .A2(new_n520_), .A3(new_n478_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT8), .B1(new_n521_), .B2(new_n463_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n479_), .A2(new_n469_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(new_n471_), .A3(new_n455_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n518_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n514_), .B1(new_n517_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT69), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n484_), .A2(new_n510_), .A3(KEYINPUT68), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G232gat), .A2(G233gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT34), .Z(new_n531_));
  INV_X1    g330(.A(KEYINPUT35), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT70), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n501_), .A2(new_n502_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n525_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n513_), .A2(new_n529_), .A3(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n531_), .A2(new_n532_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT71), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(KEYINPUT71), .A3(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n511_), .A2(new_n512_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n536_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n544_), .A2(new_n538_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT72), .B1(new_n543_), .B2(new_n547_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n537_), .A2(KEYINPUT71), .A3(new_n538_), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT71), .B1(new_n537_), .B2(new_n538_), .ZN(new_n550_));
  OAI211_X1 g349(.A(KEYINPUT72), .B(new_n547_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n454_), .B1(new_n548_), .B2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n453_), .A2(KEYINPUT36), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n554_), .B(new_n547_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n450_), .A2(KEYINPUT105), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT105), .B1(new_n450_), .B2(new_n556_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G57gat), .B(G64gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n561_));
  XOR2_X1   g360(.A(G71gat), .B(G78gat), .Z(new_n562_));
  OR2_X1    g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n562_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n484_), .A2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n470_), .B(new_n566_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT12), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G230gat), .A2(G233gat), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT12), .B1(new_n484_), .B2(new_n567_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n571_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n572_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n570_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G120gat), .B(G148gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT5), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G176gat), .B(G204gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n580_), .B(new_n581_), .Z(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n575_), .A2(new_n577_), .A3(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n586_), .A2(KEYINPUT13), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(KEYINPUT13), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G15gat), .B(G22gat), .ZN(new_n591_));
  INV_X1    g390(.A(G1gat), .ZN(new_n592_));
  INV_X1    g391(.A(G8gat), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT14), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G1gat), .B(G8gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  NAND2_X1  g396(.A1(new_n535_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n598_), .B(new_n599_), .C1(new_n517_), .C2(new_n597_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n507_), .A2(new_n508_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n595_), .B(new_n596_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n604_), .A2(KEYINPUT77), .A3(new_n599_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT77), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n598_), .A2(new_n603_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n599_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n600_), .B1(new_n605_), .B2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G113gat), .B(G141gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT78), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G169gat), .B(G197gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  AND2_X1   g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n614_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n600_), .B(new_n616_), .C1(new_n605_), .C2(new_n609_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n590_), .A2(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(G127gat), .B(G155gat), .Z(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G183gat), .B(G211gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT17), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n566_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT73), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n631_), .A2(new_n632_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n602_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n631_), .A2(new_n632_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n597_), .A3(new_n633_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT17), .B1(new_n636_), .B2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n628_), .B1(new_n639_), .B2(new_n626_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT75), .B1(new_n636_), .B2(new_n638_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n640_), .B(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n621_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n559_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n447_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(G1gat), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n546_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n454_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n555_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT37), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n547_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT72), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n651_), .B1(new_n656_), .B2(new_n551_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT37), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n555_), .A2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n653_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n643_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT76), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n417_), .A2(new_n412_), .A3(new_n408_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n387_), .A2(new_n389_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n431_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n446_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n342_), .A2(new_n433_), .A3(new_n436_), .A4(new_n438_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n342_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n669_));
  AOI22_X1  g468(.A1(new_n668_), .A2(new_n274_), .B1(new_n669_), .B2(new_n448_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(new_n621_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n662_), .A2(new_n592_), .A3(new_n447_), .A4(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n672_), .A2(new_n673_), .A3(new_n649_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n672_), .B2(new_n649_), .ZN(new_n675_));
  OAI221_X1 g474(.A(new_n648_), .B1(new_n649_), .B2(new_n672_), .C1(new_n674_), .C2(new_n675_), .ZN(G1324gat));
  XNOR2_X1  g475(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT108), .ZN(new_n679_));
  INV_X1    g478(.A(new_n445_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n680_), .B(new_n645_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G8gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT39), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT39), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n681_), .A2(new_n684_), .A3(G8gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n662_), .A2(new_n593_), .A3(new_n680_), .A4(new_n671_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n679_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n681_), .A2(new_n684_), .A3(G8gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n684_), .B1(new_n681_), .B2(G8gat), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n687_), .B(new_n679_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n678_), .B1(new_n688_), .B2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT108), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(new_n691_), .A3(new_n677_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n696_), .ZN(G1325gat));
  NAND2_X1  g496(.A1(new_n662_), .A2(new_n671_), .ZN(new_n698_));
  OR3_X1    g497(.A1(new_n698_), .A2(G15gat), .A3(new_n274_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n646_), .A2(new_n273_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n700_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT41), .B1(new_n700_), .B2(G15gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n699_), .B1(new_n701_), .B2(new_n702_), .ZN(G1326gat));
  OR3_X1    g502(.A1(new_n698_), .A2(G22gat), .A3(new_n446_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n646_), .A2(new_n342_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G22gat), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(KEYINPUT42), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(KEYINPUT42), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(G1327gat));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n710_), .B1(new_n670_), .B2(new_n660_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n659_), .ZN(new_n714_));
  AOI22_X1  g513(.A1(new_n553_), .A2(new_n714_), .B1(KEYINPUT37), .B2(new_n652_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT109), .B1(new_n450_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT43), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n713_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n590_), .A2(new_n644_), .A3(new_n620_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n718_), .A2(KEYINPUT44), .A3(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G29gat), .B1(new_n725_), .B2(new_n433_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n556_), .A2(new_n643_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n671_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n447_), .A2(new_n495_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT110), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n726_), .A2(new_n731_), .ZN(G1328gat));
  INV_X1    g531(.A(KEYINPUT46), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT44), .B1(new_n718_), .B2(new_n720_), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n722_), .B(new_n719_), .C1(new_n713_), .C2(new_n717_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n493_), .B1(new_n736_), .B2(new_n680_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n728_), .A2(new_n493_), .A3(new_n680_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT45), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n733_), .B1(new_n737_), .B2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G36gat), .B1(new_n725_), .B2(new_n445_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(KEYINPUT46), .A3(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1329gat));
  AOI21_X1  g543(.A(G43gat), .B1(new_n728_), .B2(new_n273_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT111), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n274_), .A2(new_n488_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n725_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT47), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n746_), .B(new_n751_), .C1(new_n725_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1330gat));
  AOI21_X1  g552(.A(G50gat), .B1(new_n728_), .B2(new_n342_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n446_), .A2(new_n486_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n736_), .B2(new_n755_), .ZN(G1331gat));
  NOR3_X1   g555(.A1(new_n670_), .A2(new_n620_), .A3(new_n590_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n662_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(G57gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n759_), .A3(new_n447_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n590_), .A2(new_n644_), .A3(new_n620_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n559_), .A2(new_n761_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(new_n447_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n760_), .B1(new_n763_), .B2(new_n759_), .ZN(G1332gat));
  NOR2_X1   g563(.A1(new_n445_), .A2(G64gat), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT112), .Z(new_n766_));
  NAND2_X1  g565(.A1(new_n758_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n762_), .A2(new_n680_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(G64gat), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(KEYINPUT48), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(KEYINPUT48), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(G1333gat));
  INV_X1    g571(.A(G71gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n758_), .A2(new_n773_), .A3(new_n273_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n762_), .A2(new_n273_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(G71gat), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(KEYINPUT49), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(KEYINPUT49), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(G1334gat));
  NAND3_X1  g578(.A1(new_n758_), .A2(new_n324_), .A3(new_n342_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n762_), .A2(new_n342_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(G78gat), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n782_), .A2(KEYINPUT50), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(KEYINPUT50), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(G1335gat));
  NAND2_X1  g584(.A1(new_n757_), .A2(new_n727_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT113), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n460_), .A3(new_n447_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n644_), .A2(new_n589_), .A3(new_n619_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT114), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n718_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791_), .B2(new_n433_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n788_), .A2(new_n792_), .ZN(G1336gat));
  NAND3_X1  g592(.A1(new_n787_), .A2(new_n461_), .A3(new_n680_), .ZN(new_n794_));
  OAI21_X1  g593(.A(G92gat), .B1(new_n791_), .B2(new_n445_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1337gat));
  NAND3_X1  g595(.A1(new_n787_), .A2(new_n458_), .A3(new_n273_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n791_), .A2(new_n274_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(new_n475_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT51), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n797_), .B(new_n801_), .C1(new_n475_), .C2(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1338gat));
  NOR2_X1   g602(.A1(new_n716_), .A2(KEYINPUT43), .ZN(new_n804_));
  AOI211_X1 g603(.A(KEYINPUT109), .B(new_n712_), .C1(new_n450_), .C2(new_n715_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n342_), .B(new_n790_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(KEYINPUT115), .A3(G106gat), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT115), .B1(new_n806_), .B2(G106gat), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n808_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n810_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n446_), .A2(G106gat), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n787_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT53), .B1(new_n811_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n809_), .A2(new_n810_), .B1(new_n787_), .B2(new_n813_), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n809_), .A2(new_n810_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n817_), .B(new_n818_), .C1(new_n819_), .C2(new_n808_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n816_), .A2(new_n820_), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT12), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n823_), .A2(new_n576_), .A3(new_n573_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n576_), .B1(new_n823_), .B2(new_n573_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(KEYINPUT55), .B2(new_n825_), .ZN(new_n826_));
  AND4_X1   g625(.A1(KEYINPUT55), .A2(new_n571_), .A3(new_n572_), .A4(new_n574_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n582_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n585_), .A2(KEYINPUT117), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n619_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n825_), .A2(KEYINPUT55), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n575_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n827_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n584_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n835_), .A2(KEYINPUT117), .A3(new_n829_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n831_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n517_), .A2(new_n597_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n598_), .A2(new_n608_), .ZN(new_n839_));
  OAI221_X1 g638(.A(new_n614_), .B1(new_n604_), .B2(new_n608_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n617_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n837_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n556_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n841_), .A2(new_n585_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n828_), .B2(KEYINPUT56), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n835_), .A2(new_n829_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n849_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n835_), .A2(new_n829_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n828_), .A2(KEYINPUT56), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(KEYINPUT58), .A4(new_n850_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n715_), .A2(new_n853_), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n555_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n845_), .B(KEYINPUT57), .C1(new_n858_), .C2(new_n657_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n848_), .A2(new_n857_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n644_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n640_), .A2(new_n641_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n640_), .A2(new_n641_), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n864_), .A2(new_n865_), .A3(new_n619_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n590_), .A2(new_n863_), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n643_), .A2(new_n619_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT116), .B1(new_n868_), .B2(new_n589_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n862_), .B1(new_n870_), .B2(new_n660_), .ZN(new_n871_));
  AOI211_X1 g670(.A(KEYINPUT54), .B(new_n715_), .C1(new_n869_), .C2(new_n867_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n861_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n669_), .A2(new_n447_), .A3(new_n273_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(G113gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(new_n878_), .A3(new_n620_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n859_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n843_), .B1(new_n831_), .B2(new_n836_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n853_), .A2(new_n856_), .ZN(new_n883_));
  OAI22_X1  g682(.A1(new_n882_), .A2(KEYINPUT57), .B1(new_n660_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n880_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n848_), .A2(new_n857_), .A3(KEYINPUT118), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n643_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n872_), .A2(new_n871_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n874_), .A2(KEYINPUT59), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n876_), .A2(KEYINPUT59), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n892_), .A2(new_n620_), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n879_), .B1(new_n895_), .B2(new_n878_), .ZN(G1340gat));
  INV_X1    g695(.A(G120gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n590_), .B2(KEYINPUT60), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n877_), .B(new_n898_), .C1(KEYINPUT60), .C2(new_n897_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n892_), .A2(new_n589_), .A3(new_n893_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n899_), .B1(new_n901_), .B2(new_n897_), .ZN(G1341gat));
  INV_X1    g701(.A(G127gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n877_), .A2(new_n903_), .A3(new_n643_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n892_), .A2(new_n643_), .A3(new_n893_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n904_), .B1(new_n906_), .B2(new_n903_), .ZN(G1342gat));
  NOR2_X1   g706(.A1(new_n876_), .A2(new_n556_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n909_));
  OR3_X1    g708(.A1(new_n908_), .A2(new_n909_), .A3(G134gat), .ZN(new_n910_));
  XOR2_X1   g709(.A(KEYINPUT120), .B(G134gat), .Z(new_n911_));
  NAND4_X1  g710(.A1(new_n892_), .A2(new_n715_), .A3(new_n893_), .A4(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n909_), .B1(new_n908_), .B2(G134gat), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n910_), .A2(new_n912_), .A3(new_n913_), .ZN(G1343gat));
  NAND4_X1  g713(.A1(new_n445_), .A2(new_n274_), .A3(new_n342_), .A4(new_n447_), .ZN(new_n915_));
  XOR2_X1   g714(.A(new_n915_), .B(KEYINPUT121), .Z(new_n916_));
  NAND2_X1  g715(.A1(new_n873_), .A2(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n619_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT122), .B(G141gat), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1344gat));
  NOR2_X1   g719(.A1(new_n917_), .A2(new_n590_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(G148gat), .Z(G1345gat));
  OR3_X1    g721(.A1(new_n917_), .A2(KEYINPUT123), .A3(new_n644_), .ZN(new_n923_));
  OAI21_X1  g722(.A(KEYINPUT123), .B1(new_n917_), .B2(new_n644_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT61), .B(G155gat), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1346gat));
  OAI21_X1  g727(.A(G162gat), .B1(new_n917_), .B2(new_n660_), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n556_), .A2(G162gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n917_), .B2(new_n930_), .ZN(G1347gat));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n680_), .A2(new_n448_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(new_n342_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n937_), .A2(new_n619_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n932_), .B1(new_n938_), .B2(new_n211_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n359_), .ZN(new_n940_));
  OAI211_X1 g739(.A(KEYINPUT62), .B(G169gat), .C1(new_n937_), .C2(new_n619_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n939_), .A2(new_n940_), .A3(new_n941_), .ZN(G1348gat));
  AND2_X1   g741(.A1(new_n873_), .A2(new_n446_), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n935_), .A2(new_n212_), .A3(new_n590_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n589_), .B(new_n936_), .C1(new_n888_), .C2(new_n889_), .ZN(new_n946_));
  AND3_X1   g745(.A1(new_n946_), .A2(KEYINPUT125), .A3(new_n227_), .ZN(new_n947_));
  AOI21_X1  g746(.A(KEYINPUT125), .B1(new_n946_), .B2(new_n227_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n945_), .B1(new_n947_), .B2(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(KEYINPUT126), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951_));
  OAI211_X1 g750(.A(new_n951_), .B(new_n945_), .C1(new_n947_), .C2(new_n948_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n950_), .A2(new_n952_), .ZN(G1349gat));
  NOR2_X1   g752(.A1(new_n935_), .A2(new_n644_), .ZN(new_n954_));
  AOI21_X1  g753(.A(G183gat), .B1(new_n943_), .B2(new_n954_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n937_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n644_), .B1(new_n349_), .B2(new_n223_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n955_), .B1(new_n956_), .B2(new_n957_), .ZN(G1350gat));
  OAI21_X1  g757(.A(G190gat), .B1(new_n937_), .B2(new_n660_), .ZN(new_n959_));
  INV_X1    g758(.A(new_n556_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(new_n348_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n959_), .B1(new_n937_), .B2(new_n961_), .ZN(G1351gat));
  NOR3_X1   g761(.A1(new_n445_), .A2(new_n434_), .A3(new_n273_), .ZN(new_n963_));
  AND2_X1   g762(.A1(new_n873_), .A2(new_n963_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(new_n620_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g765(.A1(new_n964_), .A2(new_n589_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g767(.A1(new_n964_), .A2(new_n643_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n970_));
  AND2_X1   g769(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n971_));
  NOR3_X1   g770(.A1(new_n969_), .A2(new_n970_), .A3(new_n971_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n972_), .B1(new_n969_), .B2(new_n970_), .ZN(G1354gat));
  INV_X1    g772(.A(G218gat), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n964_), .A2(new_n974_), .A3(new_n960_), .ZN(new_n975_));
  INV_X1    g774(.A(new_n975_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n974_), .B1(new_n964_), .B2(new_n715_), .ZN(new_n977_));
  OAI21_X1  g776(.A(KEYINPUT127), .B1(new_n976_), .B2(new_n977_), .ZN(new_n978_));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979_));
  AND2_X1   g778(.A1(new_n964_), .A2(new_n715_), .ZN(new_n980_));
  OAI211_X1 g779(.A(new_n979_), .B(new_n975_), .C1(new_n980_), .C2(new_n974_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n978_), .A2(new_n981_), .ZN(G1355gat));
endmodule


