//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT64), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(KEYINPUT9), .A3(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n217_), .A2(KEYINPUT9), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n209_), .A2(new_n213_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n206_), .A2(new_n208_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT7), .ZN(new_n222_));
  INV_X1    g021(.A(G99gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n211_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n221_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228_));
  INV_X1    g027(.A(new_n217_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n216_), .A2(KEYINPUT65), .A3(new_n217_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NOR3_X1   g032(.A1(new_n227_), .A2(KEYINPUT8), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT8), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n231_), .A2(new_n232_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n209_), .A2(new_n225_), .A3(new_n224_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n235_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n220_), .B1(new_n234_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT11), .ZN(new_n240_));
  INV_X1    g039(.A(G78gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G71gat), .ZN(new_n242_));
  INV_X1    g041(.A(G71gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G78gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G57gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(G64gat), .ZN(new_n247_));
  INV_X1    g046(.A(G64gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(G57gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT66), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(G57gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n246_), .A2(G64gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  AOI211_X1 g053(.A(new_n240_), .B(new_n245_), .C1(new_n250_), .C2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n245_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n250_), .A2(new_n254_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n256_), .B1(new_n257_), .B2(KEYINPUT11), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n250_), .A2(new_n240_), .A3(new_n254_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n255_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT12), .B1(new_n239_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n239_), .A2(new_n260_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n264_));
  INV_X1    g063(.A(new_n220_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT8), .B1(new_n227_), .B2(new_n233_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n236_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n265_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n254_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n253_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT11), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(new_n259_), .A3(new_n245_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n257_), .A2(KEYINPUT11), .A3(new_n256_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n268_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n264_), .B1(new_n275_), .B2(KEYINPUT12), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT12), .ZN(new_n277_));
  NOR4_X1   g076(.A1(new_n268_), .A2(new_n274_), .A3(KEYINPUT67), .A4(new_n277_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n204_), .B(new_n263_), .C1(new_n276_), .C2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n204_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n239_), .A2(new_n260_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n280_), .B1(new_n281_), .B2(new_n275_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G120gat), .B(G148gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT5), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G176gat), .B(G204gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  XNOR2_X1  g086(.A(new_n283_), .B(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n288_), .A2(KEYINPUT13), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(KEYINPUT13), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT73), .B(G15gat), .ZN(new_n293_));
  INV_X1    g092(.A(G22gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G8gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G1gat), .B(G8gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n298_), .B(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G29gat), .B(G36gat), .Z(new_n302_));
  XOR2_X1   g101(.A(G43gat), .B(G50gat), .Z(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G29gat), .B(G36gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G43gat), .B(G50gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n301_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n298_), .B(new_n299_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT15), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n304_), .A2(KEYINPUT15), .A3(new_n307_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G229gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT75), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n309_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT76), .ZN(new_n319_));
  INV_X1    g118(.A(new_n316_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n309_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n301_), .A2(new_n308_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n320_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n309_), .A2(new_n315_), .A3(new_n324_), .A4(new_n317_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n319_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G113gat), .B(G141gat), .Z(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT77), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G169gat), .B(G197gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n319_), .A2(new_n323_), .A3(new_n325_), .A4(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n292_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G231gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n301_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(new_n260_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G127gat), .B(G155gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT16), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G183gat), .B(G211gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT17), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n343_), .A2(KEYINPUT74), .ZN(new_n344_));
  OR3_X1    g143(.A1(new_n338_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n343_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n338_), .B(new_n346_), .C1(new_n342_), .C2(new_n344_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n335_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G227gat), .A2(G233gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n350_), .B(G15gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G43gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G71gat), .B(G99gat), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n353_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(KEYINPUT82), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G183gat), .A2(G190gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n361_), .A2(KEYINPUT80), .A3(KEYINPUT23), .A4(new_n362_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n361_), .A2(KEYINPUT23), .A3(new_n362_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT23), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(G183gat), .A3(G190gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n358_), .B(new_n363_), .C1(new_n364_), .C2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT81), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n361_), .A2(new_n362_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n367_), .B(new_n366_), .C1(new_n371_), .C2(new_n365_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n358_), .A4(new_n363_), .ZN(new_n374_));
  OR3_X1    g173(.A1(KEYINPUT79), .A2(KEYINPUT22), .A3(G176gat), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT79), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G169gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n370_), .A2(new_n374_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT30), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT25), .B(G183gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT26), .B(G190gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G169gat), .ZN(new_n384_));
  INV_X1    g183(.A(G176gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G169gat), .A2(G176gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(KEYINPUT24), .A3(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n386_), .A2(KEYINPUT24), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n383_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  MUX2_X1   g189(.A(new_n359_), .B(new_n371_), .S(new_n365_), .Z(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n379_), .A2(new_n380_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n380_), .B1(new_n379_), .B2(new_n392_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n357_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n352_), .B(new_n353_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n395_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n393_), .A4(new_n356_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n396_), .A2(new_n401_), .A3(KEYINPUT83), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT84), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n393_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n405_), .B2(new_n357_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n401_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT31), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n403_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G127gat), .B(G134gat), .Z(new_n412_));
  XOR2_X1   g211(.A(G113gat), .B(G120gat), .Z(new_n413_));
  XOR2_X1   g212(.A(new_n412_), .B(new_n413_), .Z(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n410_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n408_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n407_), .B1(new_n406_), .B2(new_n401_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT31), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n403_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n414_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G226gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n390_), .A2(KEYINPUT93), .A3(new_n372_), .A4(new_n363_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT93), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n363_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n383_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n391_), .A2(new_n358_), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT22), .B(G169gat), .Z(new_n433_));
  MUX2_X1   g232(.A(new_n384_), .B(new_n433_), .S(new_n385_), .Z(new_n434_));
  AOI22_X1  g233(.A1(new_n427_), .A2(new_n431_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G197gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT90), .ZN(new_n438_));
  INV_X1    g237(.A(G204gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n439_), .B2(G197gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT89), .B(G204gat), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n437_), .B(new_n440_), .C1(new_n441_), .C2(new_n436_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G211gat), .B(G218gat), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT21), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n443_), .B1(new_n442_), .B2(KEYINPUT21), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n439_), .A2(G197gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT88), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n441_), .A2(new_n436_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n444_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n446_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT20), .B1(new_n435_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n379_), .A2(new_n392_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(new_n452_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n426_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G8gat), .B(G36gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G64gat), .B(G92gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n455_), .A2(new_n452_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n435_), .A2(new_n453_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(KEYINPUT20), .A4(new_n425_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n457_), .A2(new_n462_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT27), .ZN(new_n467_));
  INV_X1    g266(.A(new_n463_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n432_), .A2(new_n434_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n430_), .B2(new_n429_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT20), .B1(new_n470_), .B2(new_n452_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n426_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n454_), .A2(new_n456_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n472_), .B1(new_n473_), .B2(new_n426_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n462_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT100), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(KEYINPUT100), .A3(new_n475_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n467_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n457_), .A2(new_n465_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n475_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(KEYINPUT95), .A3(new_n466_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT27), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT95), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n457_), .A2(new_n485_), .A3(new_n462_), .A4(new_n465_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n483_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT101), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT101), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n483_), .A2(new_n489_), .A3(new_n484_), .A4(new_n486_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n480_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT1), .ZN(new_n494_));
  NAND3_X1  g293(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n495_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT1), .B1(new_n497_), .B2(new_n492_), .ZN(new_n498_));
  INV_X1    g297(.A(G155gat), .ZN(new_n499_));
  INV_X1    g298(.A(G162gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n496_), .A2(new_n498_), .A3(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G141gat), .B(G148gat), .Z(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OR3_X1    g303(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT2), .ZN(new_n506_));
  INV_X1    g305(.A(G141gat), .ZN(new_n507_));
  INV_X1    g306(.A(G148gat), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n506_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n505_), .A2(new_n509_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n493_), .A2(new_n495_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n504_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT86), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT4), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n504_), .A2(KEYINPUT86), .A3(new_n514_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .A4(new_n414_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G225gat), .A2(G233gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(new_n519_), .A3(new_n414_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n504_), .A2(new_n415_), .A3(new_n514_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(KEYINPUT4), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G1gat), .B(G29gat), .Z(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G57gat), .B(G85gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  NAND3_X1  g333(.A1(new_n524_), .A2(new_n525_), .A3(new_n521_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n526_), .A2(KEYINPUT96), .A3(new_n522_), .A4(new_n520_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n529_), .A2(new_n534_), .A3(new_n535_), .A4(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n535_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT96), .B1(new_n523_), .B2(new_n526_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT99), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n537_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n517_), .A2(new_n519_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT28), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  AOI221_X4 g348(.A(new_n516_), .B1(new_n512_), .B2(new_n513_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT86), .B1(new_n504_), .B2(new_n514_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n548_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT28), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G22gat), .B(G50gat), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n549_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n549_), .B2(new_n553_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT91), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n549_), .A2(new_n553_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n554_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n549_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(G233gat), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT87), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(G228gat), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(G228gat), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n564_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n452_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n550_), .A2(new_n551_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n571_), .B1(new_n572_), .B2(KEYINPUT29), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n515_), .A2(KEYINPUT29), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n570_), .B1(new_n575_), .B2(new_n452_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G78gat), .B(G106gat), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n574_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n578_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n557_), .A2(new_n563_), .A3(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n555_), .A2(new_n556_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n584_), .A2(new_n561_), .A3(new_n581_), .A4(new_n580_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n422_), .A2(new_n491_), .A3(new_n545_), .A4(new_n586_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n543_), .A2(new_n544_), .A3(new_n586_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n537_), .A2(new_n541_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n462_), .A2(KEYINPUT32), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n590_), .B1(new_n481_), .B2(KEYINPUT98), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n457_), .A2(KEYINPUT98), .A3(new_n465_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n590_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n472_), .B(new_n593_), .C1(new_n473_), .C2(new_n426_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n591_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n589_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n526_), .A2(new_n521_), .A3(new_n520_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n524_), .A2(new_n525_), .A3(new_n522_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(new_n538_), .A3(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n457_), .A2(new_n462_), .A3(new_n465_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n462_), .B1(new_n457_), .B2(new_n465_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n485_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n486_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n599_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n537_), .A2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n539_), .A2(new_n540_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(KEYINPUT33), .A3(new_n534_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n596_), .B1(new_n604_), .B2(new_n609_), .ZN(new_n610_));
  AOI22_X1  g409(.A1(new_n491_), .A2(new_n588_), .B1(new_n610_), .B2(new_n586_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n587_), .B1(new_n611_), .B2(new_n422_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT35), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT34), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI22_X1  g415(.A1(new_n268_), .A2(new_n308_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n239_), .A2(new_n314_), .A3(KEYINPUT69), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT70), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n616_), .A2(new_n613_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT69), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n312_), .A2(new_n313_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n622_), .B1(new_n268_), .B2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .A4(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n617_), .A2(new_n618_), .A3(new_n624_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n621_), .A2(new_n620_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT70), .B1(new_n616_), .B2(new_n613_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n626_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G190gat), .B(G218gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G134gat), .B(G162gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n625_), .A2(KEYINPUT36), .A3(new_n629_), .A4(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(KEYINPUT36), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n625_), .A2(new_n629_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n635_), .B2(KEYINPUT71), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT71), .ZN(new_n637_));
  INV_X1    g436(.A(new_n634_), .ZN(new_n638_));
  AOI211_X1 g437(.A(new_n637_), .B(new_n638_), .C1(new_n625_), .C2(new_n629_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n633_), .B1(new_n636_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n349_), .A2(new_n612_), .A3(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT103), .Z(new_n644_));
  INV_X1    g443(.A(new_n545_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n202_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT104), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n291_), .B(KEYINPUT68), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n640_), .A2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n633_), .B(new_n650_), .C1(new_n636_), .C2(new_n639_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n348_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n649_), .A2(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n612_), .A2(new_n334_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n202_), .A3(new_n645_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT38), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n647_), .A2(new_n663_), .ZN(G1324gat));
  INV_X1    g463(.A(new_n491_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n661_), .A2(new_n296_), .A3(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G8gat), .B1(new_n643_), .B2(new_n491_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n667_), .A2(KEYINPUT105), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(KEYINPUT105), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n669_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n666_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(KEYINPUT40), .B(new_n666_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1325gat));
  NAND2_X1  g476(.A1(new_n644_), .A2(new_n422_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G15gat), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT107), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n681_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n422_), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n660_), .A2(G15gat), .A3(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(new_n683_), .A3(new_n685_), .ZN(G1326gat));
  XOR2_X1   g485(.A(new_n586_), .B(KEYINPUT108), .Z(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n294_), .B1(new_n644_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n661_), .A2(new_n294_), .A3(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1327gat));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n694_), .B1(new_n642_), .B2(new_n656_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n640_), .B(KEYINPUT102), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(KEYINPUT110), .A3(new_n348_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n291_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n659_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(G29gat), .B1(new_n701_), .B2(new_n645_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n335_), .A2(new_n656_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n488_), .A2(new_n490_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n480_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n588_), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n610_), .A2(new_n586_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n422_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n705_), .A2(new_n586_), .A3(new_n706_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n415_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n419_), .A2(new_n414_), .A3(new_n420_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n545_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n710_), .A2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n704_), .B(new_n654_), .C1(new_n709_), .C2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n612_), .B2(new_n654_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n703_), .B1(new_n716_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT44), .B(new_n703_), .C1(new_n716_), .C2(new_n719_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n645_), .A2(G29gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n702_), .B1(new_n724_), .B2(new_n725_), .ZN(G1328gat));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n491_), .A2(G36gat), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n700_), .B2(new_n729_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n659_), .A2(new_n699_), .A3(KEYINPUT45), .A4(new_n728_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n722_), .A2(new_n665_), .A3(new_n723_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(G36gat), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n735_), .A2(new_n736_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n734_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n737_), .A2(new_n740_), .ZN(G1329gat));
  NAND4_X1  g540(.A1(new_n722_), .A2(G43gat), .A3(new_n422_), .A4(new_n723_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n700_), .A2(new_n684_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(G43gat), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g544(.A(new_n586_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n724_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G50gat), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n687_), .A2(G50gat), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT112), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n700_), .B2(new_n750_), .ZN(G1331gat));
  NOR3_X1   g550(.A1(new_n648_), .A2(new_n348_), .A3(new_n334_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n752_), .A2(new_n612_), .A3(new_n642_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G57gat), .B1(new_n753_), .B2(new_n545_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n334_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n612_), .A2(new_n755_), .ZN(new_n756_));
  OR3_X1    g555(.A1(new_n756_), .A2(new_n292_), .A3(new_n657_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n645_), .A2(new_n246_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1332gat));
  OAI21_X1  g558(.A(G64gat), .B1(new_n753_), .B2(new_n491_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT48), .ZN(new_n761_));
  INV_X1    g560(.A(new_n757_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n248_), .A3(new_n665_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1333gat));
  OAI21_X1  g563(.A(G71gat), .B1(new_n753_), .B2(new_n684_), .ZN(new_n765_));
  XOR2_X1   g564(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n762_), .A2(new_n243_), .A3(new_n422_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1334gat));
  OAI21_X1  g568(.A(G78gat), .B1(new_n753_), .B2(new_n687_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n687_), .A2(G78gat), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT115), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n772_), .B1(new_n757_), .B2(new_n774_), .ZN(G1335gat));
  NAND3_X1  g574(.A1(new_n291_), .A2(new_n348_), .A3(new_n755_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT116), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n716_), .B2(new_n719_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G85gat), .B1(new_n778_), .B2(new_n545_), .ZN(new_n779_));
  OR3_X1    g578(.A1(new_n756_), .A2(new_n698_), .A3(new_n648_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n645_), .A2(new_n214_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(G1336gat));
  OAI21_X1  g581(.A(G92gat), .B1(new_n778_), .B2(new_n491_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n665_), .A2(new_n215_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n780_), .B2(new_n784_), .ZN(G1337gat));
  OAI21_X1  g584(.A(G99gat), .B1(new_n778_), .B2(new_n684_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n422_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n780_), .B2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g588(.A(new_n746_), .B(new_n777_), .C1(new_n716_), .C2(new_n719_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(new_n791_), .A3(G106gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n790_), .B2(G106gat), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n746_), .A2(new_n211_), .ZN(new_n794_));
  OAI22_X1  g593(.A1(new_n792_), .A2(new_n793_), .B1(new_n780_), .B2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n317_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n309_), .A2(new_n315_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n798_), .B(new_n330_), .C1(new_n799_), .C2(new_n317_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n333_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n288_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n287_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n283_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n279_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n263_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n280_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT67), .B1(new_n262_), .B2(new_n277_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n275_), .A2(new_n264_), .A3(KEYINPUT12), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n811_), .A2(KEYINPUT55), .A3(new_n204_), .A4(new_n263_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n806_), .A2(new_n808_), .A3(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n287_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n334_), .B(new_n804_), .C1(new_n814_), .C2(KEYINPUT117), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n287_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(KEYINPUT117), .A3(new_n814_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n802_), .B1(new_n816_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n797_), .B1(new_n821_), .B2(new_n696_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT118), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n288_), .A2(new_n801_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n287_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n287_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n824_), .B1(new_n828_), .B2(new_n815_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(KEYINPUT57), .A3(new_n642_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT120), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n829_), .A2(new_n832_), .A3(KEYINPUT57), .A4(new_n642_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT119), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n819_), .A2(new_n814_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n801_), .B1(new_n283_), .B2(new_n803_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n838_), .B(new_n836_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n654_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n834_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n348_), .B1(new_n823_), .B2(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n292_), .A2(new_n656_), .A3(new_n755_), .A4(new_n655_), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(KEYINPUT54), .Z(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n844_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n684_), .A2(new_n545_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n710_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n849_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(G113gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n334_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n852_), .A2(KEYINPUT59), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n822_), .A2(new_n842_), .A3(KEYINPUT121), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT57), .B1(new_n829_), .B2(new_n642_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n654_), .A2(new_n841_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n839_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n859_), .B1(new_n860_), .B2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n834_), .A2(new_n858_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n348_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n846_), .B1(new_n865_), .B2(KEYINPUT122), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n864_), .A2(new_n867_), .A3(new_n348_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n857_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  INV_X1    g669(.A(new_n852_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n848_), .B2(new_n871_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n869_), .A2(new_n872_), .A3(new_n755_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n855_), .B1(new_n873_), .B2(new_n854_), .ZN(G1340gat));
  INV_X1    g673(.A(G120gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n292_), .B2(KEYINPUT60), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n853_), .B(new_n876_), .C1(KEYINPUT60), .C2(new_n875_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n869_), .A2(new_n872_), .A3(new_n648_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n875_), .ZN(G1341gat));
  XNOR2_X1  g678(.A(new_n860_), .B(KEYINPUT118), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n862_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n656_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n656_), .B(new_n871_), .C1(new_n882_), .C2(new_n846_), .ZN(new_n883_));
  INV_X1    g682(.A(G127gat), .ZN(new_n884_));
  AOI21_X1  g683(.A(KEYINPUT123), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n883_), .A2(KEYINPUT123), .A3(new_n884_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n869_), .A2(new_n872_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n348_), .A2(new_n884_), .ZN(new_n888_));
  AOI211_X1 g687(.A(new_n885_), .B(new_n886_), .C1(new_n887_), .C2(new_n888_), .ZN(G1342gat));
  INV_X1    g688(.A(G134gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n853_), .A2(new_n890_), .A3(new_n696_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n869_), .A2(new_n872_), .A3(new_n655_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n890_), .ZN(G1343gat));
  AOI21_X1  g692(.A(new_n422_), .B1(new_n844_), .B2(new_n847_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n665_), .A2(new_n545_), .A3(new_n586_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n755_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n507_), .ZN(G1344gat));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n648_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n508_), .ZN(G1345gat));
  NOR2_X1   g699(.A1(new_n896_), .A2(new_n348_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT61), .B(G155gat), .Z(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  NOR3_X1   g702(.A1(new_n896_), .A2(new_n500_), .A3(new_n655_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n500_), .B1(new_n896_), .B2(new_n642_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  OAI211_X1 g706(.A(KEYINPUT124), .B(new_n500_), .C1(new_n896_), .C2(new_n642_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n904_), .B1(new_n907_), .B2(new_n908_), .ZN(G1347gat));
  NAND2_X1  g708(.A1(new_n865_), .A2(KEYINPUT122), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n910_), .A2(new_n847_), .A3(new_n868_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n713_), .A2(new_n491_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n911_), .A2(new_n334_), .A3(new_n687_), .A4(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G169gat), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n913_), .A2(new_n433_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n915_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n913_), .A2(G169gat), .A3(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n916_), .A2(new_n917_), .A3(new_n919_), .ZN(G1348gat));
  AOI21_X1  g719(.A(new_n688_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(new_n291_), .A3(new_n912_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n849_), .A2(new_n746_), .ZN(new_n923_));
  NOR4_X1   g722(.A1(new_n648_), .A2(new_n385_), .A3(new_n491_), .A4(new_n713_), .ZN(new_n924_));
  AOI22_X1  g723(.A1(new_n922_), .A2(new_n385_), .B1(new_n923_), .B2(new_n924_), .ZN(G1349gat));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n656_), .A3(new_n912_), .ZN(new_n926_));
  INV_X1    g725(.A(G183gat), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n713_), .A2(new_n491_), .A3(new_n381_), .A4(new_n348_), .ZN(new_n928_));
  AOI22_X1  g727(.A1(new_n926_), .A2(new_n927_), .B1(new_n921_), .B2(new_n928_), .ZN(G1350gat));
  NAND2_X1  g728(.A1(new_n921_), .A2(new_n912_), .ZN(new_n930_));
  OAI21_X1  g729(.A(G190gat), .B1(new_n930_), .B2(new_n655_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n696_), .A2(new_n382_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n930_), .B2(new_n932_), .ZN(G1351gat));
  NOR3_X1   g732(.A1(new_n491_), .A2(new_n645_), .A3(new_n586_), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n684_), .B(new_n934_), .C1(new_n882_), .C2(new_n846_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(new_n755_), .ZN(new_n936_));
  OR2_X1    g735(.A1(new_n436_), .A2(KEYINPUT126), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n436_), .A2(KEYINPUT126), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n939_), .B1(new_n936_), .B2(new_n938_), .ZN(G1352gat));
  NOR2_X1   g739(.A1(new_n935_), .A2(new_n648_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(G204gat), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n942_), .B1(new_n441_), .B2(new_n941_), .ZN(G1353gat));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n348_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n894_), .A2(new_n945_), .A3(new_n934_), .A4(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(G211gat), .ZN(new_n948_));
  INV_X1    g747(.A(new_n946_), .ZN(new_n949_));
  OAI21_X1  g748(.A(KEYINPUT127), .B1(new_n935_), .B2(new_n949_), .ZN(new_n950_));
  AND4_X1   g749(.A1(new_n944_), .A2(new_n947_), .A3(new_n948_), .A4(new_n950_), .ZN(new_n951_));
  AOI22_X1  g750(.A1(new_n947_), .A2(new_n950_), .B1(new_n944_), .B2(new_n948_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1354gat));
  OAI21_X1  g752(.A(G218gat), .B1(new_n935_), .B2(new_n655_), .ZN(new_n954_));
  OR2_X1    g753(.A1(new_n642_), .A2(G218gat), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n935_), .B2(new_n955_), .ZN(G1355gat));
endmodule


