//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n948_,
    new_n949_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n958_, new_n959_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_, new_n968_;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  OR2_X1    g003(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n205_));
  INV_X1    g004(.A(G204gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT21), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n209_), .B1(G197gat), .B2(G204gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n204_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n206_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G197gat), .A2(G204gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n209_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n212_), .A2(new_n213_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n203_), .A2(new_n209_), .ZN(new_n216_));
  AOI22_X1  g015(.A1(new_n211_), .A2(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT84), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT2), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n218_), .A2(KEYINPUT84), .A3(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n220_), .A2(new_n222_), .A3(new_n225_), .A4(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G155gat), .B(G162gat), .Z(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n223_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n232_), .A2(new_n218_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n217_), .B1(new_n236_), .B2(KEYINPUT29), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G228gat), .A2(G233gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G22gat), .B(G50gat), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n227_), .A2(new_n228_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT28), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT29), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n243_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n241_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n247_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n241_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n245_), .A3(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G78gat), .B(G106gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n248_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n253_), .A2(KEYINPUT86), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n240_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n250_), .B1(new_n249_), .B2(new_n245_), .ZN(new_n259_));
  NOR3_X1   g058(.A1(new_n246_), .A2(new_n247_), .A3(new_n241_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n239_), .B(new_n254_), .C1(new_n261_), .C2(new_n256_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G227gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(G15gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n267_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT26), .B(G190gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT25), .B(G183gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT23), .ZN(new_n276_));
  NAND3_X1  g075(.A1(KEYINPUT80), .A2(G183gat), .A3(G190gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT80), .B1(G183gat), .B2(G190gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n276_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT81), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT79), .B(KEYINPUT23), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n280_), .A2(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT80), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT23), .B1(new_n286_), .B2(new_n277_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT81), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n275_), .B1(new_n284_), .B2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(G169gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n286_), .A2(KEYINPUT23), .A3(new_n277_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n294_));
  INV_X1    g093(.A(G183gat), .ZN(new_n295_));
  INV_X1    g094(.A(G190gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n292_), .B1(new_n294_), .B2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n266_), .B1(new_n289_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT83), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n294_), .A2(new_n297_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n291_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT24), .ZN(new_n303_));
  INV_X1    g102(.A(G169gat), .ZN(new_n304_));
  INV_X1    g103(.A(G176gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n270_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n306_), .B1(new_n307_), .B2(new_n268_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n283_), .A2(new_n282_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(new_n287_), .B2(KEYINPUT81), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n280_), .A2(new_n281_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n309_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n302_), .A2(new_n313_), .A3(new_n265_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n299_), .A2(new_n300_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n300_), .B1(new_n299_), .B2(new_n314_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G71gat), .B(G99gat), .ZN(new_n318_));
  INV_X1    g117(.A(G43gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n316_), .A2(new_n317_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n299_), .A2(new_n314_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT83), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n322_), .B1(new_n326_), .B2(new_n315_), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n324_), .A2(new_n327_), .A3(KEYINPUT31), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT31), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n323_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n326_), .A2(new_n322_), .A3(new_n315_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G127gat), .B(G134gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(G113gat), .B(G120gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n328_), .A2(new_n332_), .A3(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT31), .B1(new_n324_), .B2(new_n327_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n330_), .A2(new_n331_), .A3(new_n329_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n335_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n263_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n336_), .B1(new_n328_), .B2(new_n332_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n263_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n338_), .A2(new_n335_), .A3(new_n339_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT27), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT88), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n273_), .A2(KEYINPUT89), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n273_), .A2(KEYINPUT89), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n272_), .A3(new_n354_), .ZN(new_n355_));
  AND4_X1   g154(.A1(KEYINPUT90), .A2(new_n355_), .A3(new_n294_), .A4(new_n271_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n294_), .A2(new_n271_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT90), .B1(new_n357_), .B2(new_n355_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n297_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n291_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n217_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n302_), .A2(new_n313_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n217_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT20), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n352_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n364_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT91), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n355_), .A2(new_n294_), .A3(new_n271_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT90), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n357_), .A2(KEYINPUT90), .A3(new_n355_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n371_), .A2(new_n361_), .A3(new_n217_), .A4(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n359_), .A2(KEYINPUT91), .A3(new_n217_), .A4(new_n361_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n350_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n376_), .A2(KEYINPUT20), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G8gat), .B(G36gat), .Z(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G64gat), .B(G92gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n366_), .A2(new_n378_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n366_), .B2(new_n378_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n347_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n383_), .ZN(new_n387_));
  XOR2_X1   g186(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n388_));
  NAND2_X1  g187(.A1(new_n369_), .A2(new_n217_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n284_), .A2(new_n288_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n292_), .B1(new_n390_), .B2(new_n297_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n388_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT98), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n392_), .A2(new_n393_), .B1(new_n364_), .B2(new_n363_), .ZN(new_n394_));
  OAI211_X1 g193(.A(KEYINPUT98), .B(new_n388_), .C1(new_n389_), .C2(new_n391_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n376_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n362_), .A2(new_n365_), .A3(new_n352_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n387_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n366_), .A2(new_n378_), .A3(new_n383_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(KEYINPUT27), .A3(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G85gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT0), .B(G57gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n336_), .B1(new_n236_), .B2(KEYINPUT93), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT93), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n242_), .A2(new_n407_), .A3(new_n335_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT4), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n336_), .A2(new_n242_), .A3(KEYINPUT4), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n405_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n405_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n404_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n415_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n404_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n411_), .B1(new_n409_), .B2(KEYINPUT4), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n417_), .B(new_n418_), .C1(new_n419_), .C2(new_n405_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n416_), .A2(new_n420_), .A3(KEYINPUT99), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n417_), .B1(new_n419_), .B2(new_n405_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT99), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n404_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n386_), .A2(new_n400_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n366_), .A2(new_n378_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n387_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n422_), .B(new_n404_), .C1(KEYINPUT94), .C2(KEYINPUT33), .ZN(new_n429_));
  NOR2_X1   g228(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n416_), .A2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n428_), .A2(new_n429_), .A3(new_n431_), .A4(new_n399_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n419_), .A2(new_n405_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n406_), .A2(KEYINPUT95), .A3(new_n408_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT95), .B1(new_n406_), .B2(new_n408_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n414_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(new_n436_), .A3(new_n418_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT96), .ZN(new_n438_));
  OAI211_X1 g237(.A(KEYINPUT32), .B(new_n383_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n383_), .A2(KEYINPUT32), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n366_), .A2(new_n378_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  OAI22_X1  g241(.A1(new_n432_), .A2(new_n438_), .B1(new_n442_), .B2(new_n425_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n263_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n346_), .A2(new_n426_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G113gat), .B(G141gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G169gat), .B(G197gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n446_), .B(new_n447_), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G15gat), .B(G22gat), .ZN(new_n450_));
  INV_X1    g249(.A(G1gat), .ZN(new_n451_));
  OR2_X1    g250(.A1(KEYINPUT71), .A2(G8gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(KEYINPUT71), .A2(G8gat), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT14), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n450_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G1gat), .B(G8gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n450_), .B(new_n457_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G29gat), .B(G36gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G43gat), .B(G50gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n463_), .A2(new_n464_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT15), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n463_), .A2(new_n464_), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT15), .B1(new_n470_), .B2(new_n465_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n462_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G229gat), .A2(G233gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT77), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT76), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n470_), .A2(new_n465_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n461_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n476_), .B1(new_n461_), .B2(new_n477_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n473_), .B(new_n475_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT78), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n461_), .A2(new_n477_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n461_), .A2(new_n477_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT76), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n461_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n482_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  OAI22_X1  g285(.A1(new_n480_), .A2(new_n481_), .B1(new_n486_), .B2(new_n474_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n480_), .A2(new_n481_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n449_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n478_), .A2(new_n479_), .ZN(new_n490_));
  OAI211_X1 g289(.A(G229gat), .B(G233gat), .C1(new_n490_), .C2(new_n482_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n480_), .A2(new_n481_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n484_), .A2(new_n485_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n493_), .A2(KEYINPUT78), .A3(new_n473_), .A4(new_n475_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n491_), .A2(new_n492_), .A3(new_n494_), .A4(new_n448_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n489_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n202_), .B1(new_n445_), .B2(new_n497_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n337_), .A2(new_n340_), .A3(new_n263_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n343_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n426_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n443_), .A2(new_n444_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(KEYINPUT100), .A3(new_n496_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G57gat), .B(G64gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G71gat), .B(G78gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(KEYINPUT11), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(KEYINPUT11), .ZN(new_n509_));
  INV_X1    g308(.A(new_n507_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n506_), .A2(KEYINPUT11), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n508_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G231gat), .A2(G233gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n461_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n513_), .B(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n462_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT72), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G127gat), .B(G155gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT16), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G183gat), .B(G211gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT73), .B(KEYINPUT17), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT74), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n519_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n516_), .A2(KEYINPUT72), .A3(new_n518_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n523_), .B(KEYINPUT17), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n518_), .B2(new_n516_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT75), .B1(new_n530_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT75), .ZN(new_n535_));
  AOI211_X1 g334(.A(new_n535_), .B(new_n532_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT65), .ZN(new_n538_));
  INV_X1    g337(.A(G99gat), .ZN(new_n539_));
  INV_X1    g338(.A(G106gat), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT7), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT65), .B1(G99gat), .B2(G106gat), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n545_));
  NOR2_X1   g344(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n546_));
  OAI211_X1 g345(.A(G99gat), .B(G106gat), .C1(new_n545_), .C2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n548_));
  OR2_X1    g347(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G99gat), .A2(G106gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n544_), .A2(new_n547_), .A3(new_n548_), .A4(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554_));
  NOR2_X1   g353(.A1(G85gat), .A2(G92gat), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT8), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n558_));
  NOR2_X1   g357(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n558_), .A2(new_n559_), .A3(G106gat), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT6), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n550_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n555_), .B1(new_n554_), .B2(KEYINPUT9), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT64), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT9), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n568_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n566_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n553_), .A2(new_n557_), .B1(new_n565_), .B2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n554_), .A2(new_n555_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n543_), .A2(new_n542_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n548_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n574_), .B1(new_n577_), .B2(new_n564_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n556_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n573_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n472_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT69), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n472_), .A3(KEYINPUT69), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n547_), .A2(new_n552_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n557_), .B1(new_n585_), .B2(new_n577_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n565_), .A2(new_n572_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n544_), .A2(new_n562_), .A3(new_n563_), .A4(new_n548_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT8), .B1(new_n589_), .B2(new_n574_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n477_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n583_), .A2(KEYINPUT70), .A3(new_n584_), .A4(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT35), .ZN(new_n595_));
  XOR2_X1   g394(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n593_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT35), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n468_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n470_), .A2(KEYINPUT15), .A3(new_n465_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n579_), .B2(new_n573_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n592_), .B1(new_n604_), .B2(KEYINPUT69), .ZN(new_n605_));
  INV_X1    g404(.A(new_n584_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n600_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n581_), .A2(new_n582_), .B1(new_n477_), .B2(new_n591_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n608_), .A2(KEYINPUT70), .A3(new_n584_), .A4(new_n597_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n599_), .A2(new_n607_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G190gat), .B(G218gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(KEYINPUT36), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n613_), .B(KEYINPUT36), .Z(new_n616_));
  NAND4_X1  g415(.A1(new_n599_), .A2(new_n607_), .A3(new_n609_), .A4(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT37), .B1(new_n615_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n591_), .B2(new_n513_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT12), .ZN(new_n622_));
  INV_X1    g421(.A(new_n513_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n580_), .B2(new_n623_), .ZN(new_n624_));
  AOI211_X1 g423(.A(KEYINPUT12), .B(new_n513_), .C1(new_n573_), .C2(new_n579_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n621_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n580_), .A2(new_n623_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n573_), .A2(new_n579_), .A3(new_n513_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n620_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n626_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(G120gat), .B(G148gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n631_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n626_), .A2(new_n630_), .A3(new_n636_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n638_), .A2(KEYINPUT13), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT13), .B1(new_n638_), .B2(new_n639_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n615_), .A2(KEYINPUT37), .A3(new_n617_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n537_), .A2(new_n619_), .A3(new_n642_), .A4(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n505_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT101), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n505_), .A2(new_n648_), .A3(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n425_), .A2(G1gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OR3_X1    g452(.A1(new_n650_), .A2(new_n651_), .A3(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n615_), .A2(new_n617_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n445_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n657_));
  INV_X1    g456(.A(new_n642_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(new_n497_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n529_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n660_), .A2(new_n519_), .A3(new_n527_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(new_n532_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n642_), .A2(KEYINPUT103), .A3(new_n496_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n659_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n656_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G1gat), .B1(new_n665_), .B2(new_n425_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n651_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n654_), .A2(new_n666_), .A3(new_n667_), .ZN(G1324gat));
  NAND2_X1  g467(.A1(new_n386_), .A2(new_n400_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G8gat), .B1(new_n665_), .B2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT39), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n669_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n647_), .A2(new_n649_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n672_), .A2(KEYINPUT40), .A3(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1325gat));
  NOR2_X1   g478(.A1(new_n337_), .A2(new_n340_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G15gat), .B1(new_n665_), .B2(new_n681_), .ZN(new_n682_));
  XOR2_X1   g481(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n681_), .A2(G15gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n650_), .B2(new_n685_), .ZN(G1326gat));
  OAI21_X1  g485(.A(G22gat), .B1(new_n665_), .B2(new_n343_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n343_), .A2(G22gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n650_), .B2(new_n690_), .ZN(G1327gat));
  OAI21_X1  g490(.A(new_n535_), .B1(new_n661_), .B2(new_n532_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n530_), .A2(KEYINPUT75), .A3(new_n533_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n655_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n695_), .A2(new_n658_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n505_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n425_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n700_));
  INV_X1    g499(.A(new_n643_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(new_n618_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n700_), .B1(new_n445_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n619_), .A2(new_n643_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n503_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n659_), .A2(new_n694_), .A3(new_n663_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT44), .B1(new_n707_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n700_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n503_), .B2(new_n705_), .ZN(new_n712_));
  AOI211_X1 g511(.A(KEYINPUT43), .B(new_n702_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n713_));
  OAI211_X1 g512(.A(KEYINPUT44), .B(new_n709_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n708_), .B1(new_n703_), .B2(new_n706_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n710_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n698_), .A2(G29gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n699_), .B1(new_n719_), .B2(new_n720_), .ZN(G1328gat));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722_));
  INV_X1    g521(.A(G36gat), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n716_), .A2(new_n718_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n669_), .B1(new_n717_), .B2(KEYINPUT44), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n723_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n505_), .A2(new_n723_), .A3(new_n669_), .A4(new_n696_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n722_), .B1(new_n727_), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n728_), .B(KEYINPUT45), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n725_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n732_), .B(KEYINPUT46), .C1(new_n733_), .C2(new_n723_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(G1329gat));
  NOR2_X1   g534(.A1(new_n681_), .A2(new_n319_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI211_X1 g536(.A(new_n737_), .B(new_n710_), .C1(new_n716_), .C2(new_n718_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n697_), .A2(new_n680_), .ZN(new_n739_));
  XOR2_X1   g538(.A(KEYINPUT108), .B(G43gat), .Z(new_n740_));
  AND2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT47), .B1(new_n738_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n719_), .A2(new_n736_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n739_), .A2(new_n740_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n742_), .A2(new_n746_), .ZN(G1330gat));
  AOI21_X1  g546(.A(G50gat), .B1(new_n697_), .B2(new_n263_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n263_), .A2(G50gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n719_), .B2(new_n749_), .ZN(G1331gat));
  NOR3_X1   g549(.A1(new_n694_), .A2(new_n642_), .A3(new_n496_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n656_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(G57gat), .A3(new_n698_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT110), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n445_), .A2(new_n496_), .A3(new_n642_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n694_), .A2(new_n701_), .A3(new_n618_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(G57gat), .B1(new_n759_), .B2(new_n698_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n760_), .A2(new_n761_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n755_), .A2(new_n762_), .A3(new_n763_), .ZN(G1332gat));
  OAI21_X1  g563(.A(G64gat), .B1(new_n752_), .B2(new_n670_), .ZN(new_n765_));
  XOR2_X1   g564(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n670_), .A2(G64gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n758_), .B2(new_n768_), .ZN(G1333gat));
  OR3_X1    g568(.A1(new_n758_), .A2(G71gat), .A3(new_n681_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n753_), .A2(new_n680_), .ZN(new_n771_));
  XOR2_X1   g570(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n772_));
  AND3_X1   g571(.A1(new_n771_), .A2(G71gat), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n771_), .B2(G71gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(G1334gat));
  OAI21_X1  g574(.A(G78gat), .B1(new_n752_), .B2(new_n343_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT50), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n343_), .A2(G78gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n758_), .B2(new_n778_), .ZN(G1335gat));
  INV_X1    g578(.A(new_n695_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n756_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(G85gat), .B1(new_n782_), .B2(new_n698_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n537_), .A2(new_n642_), .A3(new_n496_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT113), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n707_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n698_), .A2(G85gat), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT114), .Z(new_n788_));
  AOI21_X1  g587(.A(new_n783_), .B1(new_n786_), .B2(new_n788_), .ZN(G1336gat));
  NOR3_X1   g588(.A1(new_n781_), .A2(G92gat), .A3(new_n670_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n786_), .A2(new_n669_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(G92gat), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(G1337gat));
  NOR4_X1   g593(.A1(new_n781_), .A2(new_n681_), .A3(new_n559_), .A4(new_n558_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n786_), .A2(new_n680_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(G99gat), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n797_), .B(new_n798_), .ZN(G1338gat));
  XNOR2_X1  g598(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n263_), .B(new_n785_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(G106gat), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n802_), .A2(new_n801_), .A3(G106gat), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n782_), .A2(new_n540_), .A3(new_n263_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n800_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n805_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n807_), .B(new_n800_), .C1(new_n809_), .C2(new_n803_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n808_), .A2(new_n811_), .ZN(G1339gat));
  NOR2_X1   g611(.A1(new_n669_), .A2(new_n425_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n499_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  XOR2_X1   g614(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n816_));
  XOR2_X1   g615(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n817_));
  INV_X1    g616(.A(new_n639_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(new_n489_), .B2(new_n495_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n628_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n620_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n626_), .A2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n621_), .B(KEYINPUT55), .C1(new_n624_), .C2(new_n625_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n637_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT56), .B1(new_n825_), .B2(new_n637_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n819_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n638_), .A2(new_n639_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830_));
  INV_X1    g629(.A(new_n475_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n493_), .A2(new_n473_), .A3(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n832_), .B(new_n449_), .C1(new_n831_), .C2(new_n486_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n495_), .A2(new_n830_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n830_), .B1(new_n495_), .B2(new_n833_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n829_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n828_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n615_), .A2(new_n617_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n817_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n840_), .B(new_n655_), .C1(new_n828_), .C2(new_n836_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n825_), .A2(new_n637_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT56), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n637_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n818_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n834_), .A2(new_n835_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(new_n848_), .A3(KEYINPUT58), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n705_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n537_), .B1(new_n842_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n757_), .A2(new_n855_), .A3(new_n497_), .A4(new_n642_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT54), .B1(new_n644_), .B2(new_n496_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n815_), .B(new_n816_), .C1(new_n854_), .C2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(G113gat), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n497_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n662_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n655_), .B1(new_n828_), .B2(new_n836_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT57), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n863_), .B2(new_n817_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n852_), .A2(new_n705_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT58), .B1(new_n847_), .B2(new_n848_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n862_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n856_), .A2(new_n857_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n814_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n859_), .B(new_n861_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n662_), .B1(new_n842_), .B2(new_n853_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n496_), .B(new_n815_), .C1(new_n874_), .C2(new_n858_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n875_), .A2(new_n876_), .A3(new_n860_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n875_), .B2(new_n860_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n873_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT121), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n881_), .B(new_n873_), .C1(new_n877_), .C2(new_n878_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1340gat));
  INV_X1    g682(.A(new_n871_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT59), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n658_), .A3(new_n859_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G120gat), .ZN(new_n887_));
  INV_X1    g686(.A(G120gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n642_), .B2(KEYINPUT60), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(KEYINPUT60), .B2(new_n888_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n887_), .B1(new_n884_), .B2(new_n890_), .ZN(G1341gat));
  AOI21_X1  g690(.A(G127gat), .B1(new_n871_), .B2(new_n537_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n885_), .A2(new_n859_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT122), .B(G127gat), .Z(new_n894_));
  NOR2_X1   g693(.A1(new_n862_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n892_), .B1(new_n893_), .B2(new_n895_), .ZN(G1342gat));
  NAND3_X1  g695(.A1(new_n885_), .A2(new_n705_), .A3(new_n859_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G134gat), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n838_), .A2(G134gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n884_), .B2(new_n899_), .ZN(G1343gat));
  NAND2_X1  g699(.A1(new_n869_), .A2(new_n870_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n813_), .A2(new_n500_), .ZN(new_n902_));
  XOR2_X1   g701(.A(new_n902_), .B(KEYINPUT123), .Z(new_n903_));
  AND2_X1   g702(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n496_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n658_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g707(.A1(new_n904_), .A2(new_n537_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT61), .B(G155gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1346gat));
  AND3_X1   g710(.A1(new_n901_), .A2(new_n655_), .A3(new_n903_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n913_));
  OR3_X1    g712(.A1(new_n912_), .A2(new_n913_), .A3(G162gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n912_), .B2(G162gat), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n705_), .A2(G162gat), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n914_), .A2(new_n915_), .B1(new_n904_), .B2(new_n916_), .ZN(G1347gat));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n854_), .A2(new_n858_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n670_), .A2(new_n698_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n345_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n919_), .A2(new_n497_), .A3(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT22), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n918_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(G169gat), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n304_), .B1(new_n924_), .B2(new_n918_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(G1348gat));
  NOR2_X1   g728(.A1(new_n919_), .A2(new_n923_), .ZN(new_n930_));
  AOI21_X1  g729(.A(G176gat), .B1(new_n930_), .B2(new_n658_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n263_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n920_), .A2(new_n680_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n933_), .A2(new_n305_), .A3(new_n642_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n931_), .B1(new_n932_), .B2(new_n934_), .ZN(G1349gat));
  NAND2_X1  g734(.A1(new_n353_), .A2(new_n354_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n930_), .A2(new_n936_), .A3(new_n662_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n933_), .A2(new_n694_), .ZN(new_n938_));
  AOI21_X1  g737(.A(KEYINPUT125), .B1(new_n932_), .B2(new_n938_), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n343_), .B(new_n938_), .C1(new_n874_), .C2(new_n858_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n295_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n937_), .B1(new_n939_), .B2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(KEYINPUT126), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n937_), .B(new_n945_), .C1(new_n939_), .C2(new_n942_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n944_), .A2(new_n946_), .ZN(G1350gat));
  NAND3_X1  g746(.A1(new_n930_), .A2(new_n272_), .A3(new_n655_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n919_), .A2(new_n702_), .A3(new_n923_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n296_), .B2(new_n949_), .ZN(G1351gat));
  NOR2_X1   g749(.A1(new_n921_), .A2(new_n341_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n901_), .A2(new_n496_), .A3(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(G197gat), .ZN(new_n953_));
  OR3_X1    g752(.A1(new_n952_), .A2(KEYINPUT127), .A3(new_n953_), .ZN(new_n954_));
  OAI21_X1  g753(.A(KEYINPUT127), .B1(new_n952_), .B2(new_n953_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n952_), .A2(new_n953_), .ZN(new_n956_));
  AND3_X1   g755(.A1(new_n954_), .A2(new_n955_), .A3(new_n956_), .ZN(G1352gat));
  AND2_X1   g756(.A1(new_n901_), .A2(new_n951_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n658_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g759(.A1(new_n958_), .A2(new_n662_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(KEYINPUT63), .B(G211gat), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n961_), .A2(new_n962_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n963_), .B1(new_n961_), .B2(new_n964_), .ZN(G1354gat));
  INV_X1    g764(.A(G218gat), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n958_), .A2(new_n966_), .A3(new_n655_), .ZN(new_n967_));
  AND2_X1   g766(.A1(new_n958_), .A2(new_n705_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n967_), .B1(new_n968_), .B2(new_n966_), .ZN(G1355gat));
endmodule


