//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n956_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_;
  INV_X1    g000(.A(KEYINPUT9), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G92gat), .ZN(new_n203_));
  INV_X1    g002(.A(G85gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n207_), .B1(new_n208_), .B2(KEYINPUT9), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n206_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G99gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT10), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT10), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G99gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(G106gat), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  AND4_X1   g019(.A1(KEYINPUT65), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n221_));
  NOR3_X1   g020(.A1(new_n215_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n210_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n208_), .A2(new_n207_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n226_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n228_));
  INV_X1    g027(.A(G106gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n211_), .B(new_n229_), .C1(new_n230_), .C2(KEYINPUT66), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(KEYINPUT66), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n224_), .B(new_n225_), .C1(new_n228_), .C2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AND3_X1   g034(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n238_), .A2(new_n227_), .A3(new_n232_), .A4(new_n231_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n224_), .B1(new_n239_), .B2(new_n225_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n223_), .B1(new_n235_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n225_), .B1(new_n228_), .B2(new_n233_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT8), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(new_n234_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(KEYINPUT67), .A3(new_n223_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT11), .ZN(new_n248_));
  XOR2_X1   g047(.A(G71gat), .B(G78gat), .Z(new_n249_));
  NAND2_X1  g048(.A1(G57gat), .A2(G64gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(G57gat), .A2(G64gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT68), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n252_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(new_n250_), .ZN(new_n256_));
  AOI211_X1 g055(.A(new_n248_), .B(new_n249_), .C1(new_n253_), .C2(new_n256_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n256_), .A2(new_n253_), .A3(new_n248_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n248_), .B1(new_n256_), .B2(new_n253_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n257_), .B1(new_n260_), .B2(new_n249_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n243_), .A2(new_n247_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n241_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT71), .B1(new_n246_), .B2(new_n223_), .ZN(new_n267_));
  OAI211_X1 g066(.A(KEYINPUT12), .B(new_n261_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G230gat), .A2(G233gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n261_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n246_), .A2(KEYINPUT67), .A3(new_n223_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT67), .B1(new_n246_), .B2(new_n223_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n264_), .A2(new_n268_), .A3(new_n269_), .A4(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n243_), .A2(new_n247_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT69), .B1(new_n276_), .B2(new_n270_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n278_));
  AOI211_X1 g077(.A(new_n278_), .B(new_n261_), .C1(new_n243_), .C2(new_n247_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT70), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n273_), .A2(new_n278_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n276_), .A2(KEYINPUT69), .A3(new_n270_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(new_n284_), .A3(new_n262_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n269_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n275_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G120gat), .B(G148gat), .Z(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(G204gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT5), .ZN(new_n290_));
  INV_X1    g089(.A(G176gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n287_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n285_), .A2(new_n286_), .ZN(new_n295_));
  AND4_X1   g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n274_), .A4(new_n292_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(new_n287_), .B2(new_n292_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n293_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT13), .ZN(new_n302_));
  OAI221_X1 g101(.A(new_n293_), .B1(KEYINPUT73), .B2(new_n302_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G113gat), .B(G141gat), .ZN(new_n305_));
  INV_X1    g104(.A(G169gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G197gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G50gat), .ZN(new_n310_));
  OR2_X1    g109(.A1(G29gat), .A2(G36gat), .ZN(new_n311_));
  INV_X1    g110(.A(G43gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G29gat), .A2(G36gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n310_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G29gat), .B(G36gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G43gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(G50gat), .A3(new_n314_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n317_), .A2(KEYINPUT15), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT15), .B1(new_n317_), .B2(new_n320_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G15gat), .B(G22gat), .ZN(new_n324_));
  INV_X1    g123(.A(G1gat), .ZN(new_n325_));
  INV_X1    g124(.A(G8gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT14), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G1gat), .B(G8gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n323_), .A2(new_n331_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n315_), .A2(new_n310_), .A3(new_n316_), .ZN(new_n333_));
  AOI21_X1  g132(.A(G50gat), .B1(new_n319_), .B2(new_n314_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT80), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n317_), .A2(new_n320_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT80), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n339_), .A3(new_n331_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n340_), .A2(KEYINPUT81), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(KEYINPUT81), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n332_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G229gat), .A2(G233gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n335_), .A2(KEYINPUT80), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n337_), .A2(new_n338_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n330_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT82), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n341_), .A2(new_n342_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n344_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n309_), .B1(new_n346_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n309_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n350_), .A2(new_n351_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n345_), .B(new_n354_), .C1(new_n355_), .C2(new_n344_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G231gat), .A2(G233gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n330_), .B(new_n359_), .Z(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(new_n270_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT79), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT16), .B(G183gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G211gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(G127gat), .B(G155gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT17), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n362_), .B(new_n368_), .Z(new_n369_));
  INV_X1    g168(.A(new_n361_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(new_n367_), .A3(new_n366_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n304_), .A2(new_n358_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n276_), .A2(new_n335_), .ZN(new_n376_));
  OAI22_X1  g175(.A1(new_n266_), .A2(new_n267_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G232gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT34), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n379_), .A2(KEYINPUT35), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT75), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n381_), .B1(new_n379_), .B2(KEYINPUT35), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n380_), .B(new_n382_), .ZN(new_n383_));
  AND4_X1   g182(.A1(KEYINPUT76), .A2(new_n376_), .A3(new_n377_), .A4(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n376_), .A2(new_n377_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT76), .B1(new_n385_), .B2(new_n380_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n376_), .A2(new_n377_), .A3(new_n383_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n384_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT74), .B(G134gat), .ZN(new_n389_));
  INV_X1    g188(.A(G162gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G190gat), .B(G218gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT36), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n393_), .A2(new_n394_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n388_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n337_), .B1(new_n243_), .B2(new_n247_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n241_), .A2(new_n265_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n246_), .A2(KEYINPUT71), .A3(new_n223_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n323_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n380_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT76), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n387_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n376_), .A2(new_n377_), .A3(KEYINPUT76), .A4(new_n383_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n395_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT77), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT77), .ZN(new_n410_));
  AOI211_X1 g209(.A(new_n410_), .B(new_n395_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n375_), .B(new_n398_), .C1(new_n409_), .C2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT37), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n410_), .B1(new_n388_), .B2(new_n395_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n407_), .A2(KEYINPUT77), .A3(new_n408_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n417_), .A2(new_n375_), .A3(KEYINPUT37), .A4(new_n398_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n414_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G228gat), .A2(G233gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT29), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n423_));
  NOR2_X1   g222(.A1(G155gat), .A2(G162gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G155gat), .A2(G162gat), .ZN(new_n426_));
  OR3_X1    g225(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G141gat), .A2(G148gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT2), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n427_), .A2(new_n430_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n425_), .A2(KEYINPUT94), .A3(new_n426_), .A4(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n423_), .A2(new_n424_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT93), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT92), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT92), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT93), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n437_), .A2(new_n439_), .A3(new_n424_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n433_), .B(new_n426_), .C1(new_n435_), .C2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT94), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n434_), .A2(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n426_), .B(KEYINPUT1), .Z(new_n445_));
  NAND2_X1  g244(.A1(new_n425_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(G141gat), .ZN(new_n447_));
  INV_X1    g246(.A(G148gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n446_), .A2(new_n428_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n422_), .B1(new_n444_), .B2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G211gat), .B(G218gat), .ZN(new_n452_));
  XOR2_X1   g251(.A(G197gat), .B(G204gat), .Z(new_n453_));
  OAI21_X1  g252(.A(new_n452_), .B1(new_n453_), .B2(KEYINPUT21), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(KEYINPUT21), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n421_), .B1(new_n451_), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G197gat), .B(G204gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT21), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n454_), .B(new_n460_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n425_), .A2(new_n445_), .B1(G141gat), .B2(G148gat), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n449_), .A2(new_n462_), .B1(new_n434_), .B2(new_n443_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n461_), .B(new_n420_), .C1(new_n463_), .C2(new_n422_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n457_), .A2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G78gat), .B(G106gat), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n457_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n466_), .B1(new_n457_), .B2(new_n464_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT96), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n444_), .A2(new_n450_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n473_), .B1(new_n474_), .B2(KEYINPUT29), .ZN(new_n475_));
  INV_X1    g274(.A(new_n473_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n463_), .A2(new_n422_), .A3(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G22gat), .B(G50gat), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n475_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n480_));
  OAI22_X1  g279(.A1(new_n471_), .A2(new_n472_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n470_), .B(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G1gat), .B(G29gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(G57gat), .B(G85gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G225gat), .A2(G233gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G113gat), .A2(G120gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G113gat), .A2(G120gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(KEYINPUT89), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT89), .ZN(new_n494_));
  INV_X1    g293(.A(new_n492_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n494_), .B1(new_n495_), .B2(new_n490_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G127gat), .B(G134gat), .Z(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n493_), .A2(new_n496_), .A3(new_n498_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(new_n444_), .A3(new_n450_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT90), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n505_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n500_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n501_), .A2(new_n504_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT91), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(new_n499_), .A3(new_n506_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n503_), .B1(new_n513_), .B2(new_n463_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT4), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n474_), .A2(new_n512_), .A3(new_n509_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT4), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n489_), .B1(new_n515_), .B2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n516_), .A2(new_n489_), .A3(new_n503_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n488_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT102), .ZN(new_n523_));
  INV_X1    g322(.A(new_n489_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n517_), .B1(new_n516_), .B2(new_n503_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n513_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT4), .B1(new_n526_), .B2(new_n474_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n524_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(new_n520_), .A3(new_n487_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n522_), .A2(new_n523_), .A3(new_n529_), .ZN(new_n530_));
  OAI211_X1 g329(.A(KEYINPUT102), .B(new_n488_), .C1(new_n519_), .C2(new_n521_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G226gat), .A2(G233gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n533_), .B(KEYINPUT97), .Z(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT19), .Z(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G183gat), .A2(G190gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT23), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT23), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n539_), .A2(G183gat), .A3(G190gat), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n540_), .A3(KEYINPUT85), .ZN(new_n541_));
  NOR2_X1   g340(.A1(G183gat), .A2(G190gat), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT85), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n544_), .A2(new_n539_), .A3(G183gat), .A4(G190gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT86), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G169gat), .A2(G176gat), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n306_), .A2(KEYINPUT22), .ZN(new_n550_));
  AOI21_X1  g349(.A(G176gat), .B1(new_n550_), .B2(KEYINPUT84), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT84), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT22), .B1(new_n552_), .B2(new_n306_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n549_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n541_), .A2(new_n555_), .A3(new_n543_), .A4(new_n545_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n547_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT25), .B(G183gat), .ZN(new_n558_));
  AND3_X1   g357(.A1(KEYINPUT83), .A2(KEYINPUT26), .A3(G190gat), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT26), .B1(KEYINPUT83), .B2(G190gat), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n306_), .A2(new_n291_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(KEYINPUT24), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n538_), .A2(new_n540_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n562_), .A2(KEYINPUT24), .A3(new_n548_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n561_), .A2(new_n564_), .A3(new_n565_), .A4(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n456_), .B1(new_n557_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n548_), .A2(KEYINPUT24), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT98), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT98), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n548_), .A2(new_n571_), .A3(KEYINPUT24), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(new_n562_), .A3(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT26), .B(G190gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n558_), .A2(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n573_), .A2(new_n545_), .A3(new_n541_), .A4(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n542_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(new_n549_), .ZN(new_n578_));
  XOR2_X1   g377(.A(KEYINPUT22), .B(G169gat), .Z(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(G176gat), .ZN(new_n580_));
  OAI22_X1  g379(.A1(new_n576_), .A2(new_n563_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT20), .B1(new_n581_), .B2(new_n461_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n536_), .B1(new_n568_), .B2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n456_), .A2(new_n567_), .A3(new_n557_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n461_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(KEYINPUT20), .A4(new_n535_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT18), .B(G64gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(G92gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G8gat), .B(G36gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n587_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT99), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT100), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n596_), .B1(new_n587_), .B2(new_n592_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n583_), .A2(KEYINPUT100), .A3(new_n591_), .A4(new_n586_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n587_), .A2(KEYINPUT99), .A3(new_n592_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n595_), .A2(new_n597_), .A3(new_n598_), .A4(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT27), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n591_), .B(KEYINPUT103), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT20), .ZN(new_n604_));
  INV_X1    g403(.A(new_n581_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n605_), .B2(new_n456_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n557_), .A2(new_n567_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n461_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n536_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  AND4_X1   g408(.A1(KEYINPUT20), .A2(new_n584_), .A3(new_n585_), .A4(new_n536_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n603_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n593_), .A2(new_n611_), .A3(KEYINPUT27), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT104), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n593_), .A2(new_n611_), .A3(KEYINPUT104), .A4(KEYINPUT27), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n602_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n482_), .B1(new_n532_), .B2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(G15gat), .B(G43gat), .Z(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT87), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G71gat), .B(G99gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G227gat), .A2(G233gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n622_), .B(new_n623_), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n607_), .B(KEYINPUT30), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT88), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT31), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n624_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n628_), .B1(new_n624_), .B2(new_n627_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n526_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n625_), .A2(new_n626_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n624_), .A2(new_n627_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT31), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n513_), .A3(new_n629_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n632_), .A2(new_n633_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n633_), .B1(new_n632_), .B2(new_n636_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n529_), .A2(KEYINPUT33), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n528_), .A2(new_n642_), .A3(new_n520_), .A4(new_n487_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n489_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n516_), .A2(new_n524_), .A3(new_n503_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n645_), .A2(new_n488_), .A3(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n600_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n644_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n468_), .A2(new_n469_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n481_), .B(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n609_), .A2(new_n610_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n592_), .A2(KEYINPUT32), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n587_), .B2(new_n653_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n530_), .A2(new_n531_), .A3(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n649_), .A2(new_n651_), .A3(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n618_), .A2(new_n640_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n659_), .B1(new_n617_), .B2(new_n482_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n532_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n651_), .A2(KEYINPUT105), .A3(new_n616_), .A4(new_n602_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n639_), .A4(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n419_), .B1(new_n658_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n374_), .A2(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n665_), .A2(G1gat), .A3(new_n661_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n407_), .A2(new_n408_), .A3(new_n396_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n658_), .B2(new_n663_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n374_), .A2(new_n669_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n672_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT107), .B1(new_n674_), .B2(new_n373_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G1gat), .B1(new_n676_), .B2(new_n661_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n668_), .A2(new_n677_), .ZN(G1324gat));
  NAND4_X1  g477(.A1(new_n374_), .A2(new_n326_), .A3(new_n617_), .A4(new_n664_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n374_), .A2(new_n617_), .A3(new_n672_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT39), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n680_), .A2(new_n681_), .A3(G8gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n680_), .B2(G8gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n679_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT108), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n686_), .B(new_n679_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n685_), .A2(KEYINPUT40), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT40), .B1(new_n685_), .B2(new_n687_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1325gat));
  INV_X1    g489(.A(G15gat), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n374_), .A2(new_n691_), .A3(new_n639_), .A4(new_n664_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n640_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(new_n691_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(KEYINPUT41), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n693_), .A2(new_n696_), .A3(new_n691_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n692_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT109), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n700_), .B(new_n692_), .C1(new_n695_), .C2(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1326gat));
  OAI21_X1  g501(.A(G22gat), .B1(new_n676_), .B2(new_n651_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT42), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n651_), .A2(G22gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n665_), .B2(new_n705_), .ZN(G1327gat));
  INV_X1    g505(.A(new_n372_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n671_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT113), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n658_), .A2(new_n663_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n304_), .A2(new_n358_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G29gat), .B1(new_n714_), .B2(new_n532_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n414_), .A2(new_n418_), .A3(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n414_), .B2(new_n418_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n716_), .B1(new_n720_), .B2(new_n710_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n710_), .A2(new_n716_), .A3(new_n419_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n713_), .B(new_n707_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT112), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n719_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n414_), .A2(new_n418_), .A3(new_n717_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n710_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT43), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n710_), .A2(new_n716_), .A3(new_n419_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n712_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(KEYINPUT44), .A4(new_n707_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n725_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n735_), .A2(new_n661_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n723_), .A2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(G29gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n715_), .B1(new_n736_), .B2(new_n739_), .ZN(G1328gat));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n741_));
  INV_X1    g540(.A(G36gat), .ZN(new_n742_));
  INV_X1    g541(.A(new_n617_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n723_), .B2(new_n737_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n734_), .B2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n714_), .A2(new_n742_), .A3(new_n617_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT45), .Z(new_n747_));
  OAI21_X1  g546(.A(new_n741_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n746_), .B(KEYINPUT45), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n738_), .A2(new_n617_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n725_), .B2(new_n733_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT46), .B(new_n749_), .C1(new_n751_), .C2(new_n742_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n748_), .A2(new_n752_), .ZN(G1329gat));
  AOI21_X1  g552(.A(new_n312_), .B1(new_n723_), .B2(new_n737_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n734_), .A2(new_n639_), .A3(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n714_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n312_), .B1(new_n756_), .B2(new_n640_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT47), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n755_), .A2(new_n760_), .A3(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1330gat));
  AOI21_X1  g561(.A(G50gat), .B1(new_n714_), .B2(new_n482_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n735_), .A2(new_n651_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n310_), .B1(new_n723_), .B2(new_n737_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(G1331gat));
  NAND3_X1  g565(.A1(new_n301_), .A2(new_n303_), .A3(new_n357_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n767_), .A2(new_n707_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n672_), .ZN(new_n769_));
  INV_X1    g568(.A(G57gat), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n661_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n768_), .A2(new_n664_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n532_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n771_), .B1(new_n770_), .B2(new_n774_), .ZN(G1332gat));
  OAI21_X1  g574(.A(G64gat), .B1(new_n769_), .B2(new_n743_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT48), .Z(new_n777_));
  NOR3_X1   g576(.A1(new_n772_), .A2(G64gat), .A3(new_n743_), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1333gat));
  OAI21_X1  g578(.A(G71gat), .B1(new_n769_), .B2(new_n640_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT49), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n640_), .A2(G71gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n772_), .B2(new_n782_), .ZN(G1334gat));
  OAI21_X1  g582(.A(G78gat), .B1(new_n769_), .B2(new_n651_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT50), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n651_), .A2(G78gat), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT114), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n785_), .B1(new_n772_), .B2(new_n787_), .ZN(G1335gat));
  INV_X1    g587(.A(new_n767_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n711_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G85gat), .B1(new_n790_), .B2(new_n532_), .ZN(new_n791_));
  AOI211_X1 g590(.A(new_n372_), .B(new_n767_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n792_), .A2(G85gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n791_), .B1(new_n793_), .B2(new_n532_), .ZN(G1336gat));
  AOI21_X1  g593(.A(G92gat), .B1(new_n790_), .B2(new_n617_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n743_), .A2(new_n203_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n792_), .B2(new_n796_), .ZN(G1337gat));
  AOI21_X1  g596(.A(new_n211_), .B1(new_n792_), .B2(new_n639_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n640_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n790_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(G1338gat));
  NAND3_X1  g601(.A1(new_n790_), .A2(new_n229_), .A3(new_n482_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n767_), .A2(new_n372_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n482_), .B(new_n807_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n808_), .A2(new_n809_), .A3(G106gat), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n808_), .B2(G106gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n806_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n808_), .A2(G106gat), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT117), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n808_), .A2(new_n809_), .A3(G106gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(KEYINPUT52), .A3(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n805_), .A2(new_n812_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT53), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n805_), .A2(new_n812_), .A3(new_n816_), .A4(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n264_), .A2(new_n269_), .A3(new_n268_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(KEYINPUT55), .A4(new_n273_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n277_), .A2(new_n279_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n264_), .A2(new_n268_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n286_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT120), .B1(new_n274_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n274_), .A2(new_n829_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n825_), .A2(new_n828_), .A3(new_n830_), .A4(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n292_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n832_), .A2(KEYINPUT56), .A3(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n295_), .A2(new_n274_), .A3(new_n292_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT72), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n287_), .A2(new_n294_), .A3(new_n292_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n357_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n344_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n343_), .A2(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n309_), .B(new_n844_), .C1(new_n355_), .C2(new_n843_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n356_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n838_), .A2(new_n842_), .B1(new_n298_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n822_), .B1(new_n848_), .B2(new_n671_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n671_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n842_), .A2(new_n838_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n840_), .A2(new_n841_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n846_), .B1(new_n852_), .B2(new_n293_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT57), .B(new_n850_), .C1(new_n851_), .C2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n832_), .A2(KEYINPUT56), .A3(new_n833_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT56), .B1(new_n832_), .B2(new_n833_), .ZN(new_n857_));
  OAI22_X1  g656(.A1(new_n856_), .A2(new_n857_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n855_), .B1(new_n858_), .B2(new_n846_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n838_), .A2(KEYINPUT58), .A3(new_n852_), .A4(new_n847_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n419_), .A3(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n849_), .A2(new_n854_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n707_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n419_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n707_), .A2(new_n358_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n304_), .A2(new_n864_), .A3(new_n866_), .A4(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT119), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n419_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n870_), .A2(new_n871_), .A3(new_n866_), .A4(new_n867_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n304_), .A2(new_n864_), .A3(new_n867_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n865_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n869_), .A2(new_n872_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n863_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n660_), .A2(new_n639_), .A3(new_n662_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n661_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(KEYINPUT59), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n876_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n876_), .A2(KEYINPUT122), .A3(new_n880_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n862_), .A2(new_n885_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n849_), .A2(new_n854_), .A3(KEYINPUT121), .A4(new_n861_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n707_), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n879_), .B1(new_n888_), .B2(new_n875_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n883_), .B(new_n884_), .C1(new_n889_), .C2(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(G113gat), .B1(new_n891_), .B2(new_n357_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n889_), .ZN(new_n893_));
  OR3_X1    g692(.A1(new_n893_), .A2(G113gat), .A3(new_n357_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1340gat));
  OAI21_X1  g694(.A(G120gat), .B1(new_n891_), .B2(new_n304_), .ZN(new_n896_));
  INV_X1    g695(.A(G120gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n304_), .B2(KEYINPUT60), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n889_), .B(new_n898_), .C1(KEYINPUT60), .C2(new_n897_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n899_), .ZN(G1341gat));
  OAI21_X1  g699(.A(G127gat), .B1(new_n891_), .B2(new_n707_), .ZN(new_n901_));
  OR3_X1    g700(.A1(new_n893_), .A2(G127gat), .A3(new_n707_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1342gat));
  OAI21_X1  g702(.A(G134gat), .B1(new_n891_), .B2(new_n864_), .ZN(new_n904_));
  OR3_X1    g703(.A1(new_n893_), .A2(G134gat), .A3(new_n850_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1343gat));
  NAND2_X1  g705(.A1(new_n888_), .A2(new_n875_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n661_), .A2(new_n639_), .A3(new_n651_), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n907_), .A2(new_n743_), .A3(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n358_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G141gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n909_), .A2(new_n447_), .A3(new_n358_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1344gat));
  INV_X1    g712(.A(new_n304_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n909_), .A2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(G148gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n909_), .A2(new_n448_), .A3(new_n914_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1345gat));
  NAND4_X1  g717(.A1(new_n907_), .A2(new_n372_), .A3(new_n743_), .A4(new_n908_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(KEYINPUT61), .B(G155gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n919_), .B(new_n920_), .ZN(G1346gat));
  NAND2_X1  g720(.A1(new_n909_), .A2(new_n671_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n718_), .A2(new_n719_), .A3(new_n390_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n922_), .A2(new_n390_), .B1(new_n909_), .B2(new_n923_), .ZN(G1347gat));
  NAND3_X1  g723(.A1(new_n661_), .A2(new_n639_), .A3(new_n617_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n358_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n876_), .A2(new_n930_), .A3(new_n651_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(G169gat), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT62), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n927_), .A2(new_n651_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n876_), .A2(new_n934_), .ZN(new_n935_));
  OR3_X1    g734(.A1(new_n935_), .A2(new_n357_), .A3(new_n579_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n933_), .A2(new_n936_), .ZN(G1348gat));
  NAND4_X1  g736(.A1(new_n907_), .A2(G176gat), .A3(new_n914_), .A4(new_n934_), .ZN(new_n938_));
  OR2_X1    g737(.A1(new_n938_), .A2(KEYINPUT125), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n291_), .B1(new_n935_), .B2(new_n304_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n938_), .A2(KEYINPUT125), .ZN(new_n941_));
  AND3_X1   g740(.A1(new_n939_), .A2(new_n940_), .A3(new_n941_), .ZN(G1349gat));
  NOR3_X1   g741(.A1(new_n935_), .A2(new_n707_), .A3(new_n558_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n907_), .A2(new_n372_), .A3(new_n934_), .ZN(new_n944_));
  INV_X1    g743(.A(G183gat), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n943_), .B1(new_n944_), .B2(new_n945_), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n935_), .B2(new_n864_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n671_), .A2(new_n574_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n935_), .B2(new_n948_), .ZN(G1351gat));
  NOR3_X1   g748(.A1(new_n639_), .A2(new_n532_), .A3(new_n651_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(KEYINPUT126), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(new_n617_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n952_), .B1(new_n888_), .B2(new_n875_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(new_n358_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g754(.A1(new_n953_), .A2(new_n914_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g756(.A1(new_n953_), .A2(new_n372_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  AND2_X1   g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n958_), .B1(new_n959_), .B2(new_n960_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n961_), .B1(new_n958_), .B2(new_n959_), .ZN(G1354gat));
  INV_X1    g761(.A(G218gat), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n963_), .B1(new_n953_), .B2(new_n419_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n671_), .A2(new_n963_), .ZN(new_n965_));
  AOI211_X1 g764(.A(new_n952_), .B(new_n965_), .C1(new_n888_), .C2(new_n875_), .ZN(new_n966_));
  OAI21_X1  g765(.A(KEYINPUT127), .B1(new_n964_), .B2(new_n966_), .ZN(new_n967_));
  INV_X1    g766(.A(new_n965_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n953_), .A2(new_n968_), .ZN(new_n969_));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970_));
  AOI211_X1 g769(.A(new_n864_), .B(new_n952_), .C1(new_n888_), .C2(new_n875_), .ZN(new_n971_));
  OAI211_X1 g770(.A(new_n969_), .B(new_n970_), .C1(new_n971_), .C2(new_n963_), .ZN(new_n972_));
  AND2_X1   g771(.A1(new_n967_), .A2(new_n972_), .ZN(G1355gat));
endmodule


