//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_;
  AOI21_X1  g000(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND3_X1  g002(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n204_), .A3(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n209_));
  OR3_X1    g008(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT24), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n212_), .B1(G169gat), .B2(G176gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT78), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT24), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n218_), .A2(new_n219_), .A3(new_n214_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n222_));
  AND3_X1   g021(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n202_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n205_), .A2(KEYINPUT25), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT25), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(G183gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n206_), .A2(KEYINPUT26), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G190gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .A4(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n211_), .B1(new_n221_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT79), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n231_), .B(new_n224_), .C1(new_n216_), .C2(new_n220_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT79), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n211_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G71gat), .B(G99gat), .ZN(new_n239_));
  INV_X1    g038(.A(G43gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n238_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT80), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G113gat), .B(G120gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n242_), .B(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G227gat), .A2(G233gat), .ZN(new_n248_));
  INV_X1    g047(.A(G15gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT30), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT31), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n247_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n247_), .A2(new_n253_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G22gat), .B(G50gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G141gat), .A2(G148gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT81), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G141gat), .ZN(new_n263_));
  INV_X1    g062(.A(G148gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT82), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(KEYINPUT1), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n269_), .B1(KEYINPUT1), .B2(new_n267_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n262_), .A2(new_n266_), .A3(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G155gat), .B(G162gat), .Z(new_n272_));
  NOR2_X1   g071(.A1(new_n261_), .A2(KEYINPUT2), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n265_), .A2(KEYINPUT3), .ZN(new_n274_));
  INV_X1    g073(.A(new_n259_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT2), .ZN(new_n276_));
  OR3_X1    g075(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  OAI211_X1 g077(.A(KEYINPUT83), .B(new_n272_), .C1(new_n273_), .C2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n275_), .A2(KEYINPUT2), .B1(new_n265_), .B2(KEYINPUT3), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n281_), .B(new_n277_), .C1(new_n261_), .C2(KEYINPUT2), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT83), .B1(new_n282_), .B2(new_n272_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n271_), .B1(new_n280_), .B2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n284_), .A2(KEYINPUT29), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT28), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n285_), .A2(new_n286_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n258_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n289_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(new_n287_), .A3(new_n257_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT90), .ZN(new_n294_));
  INV_X1    g093(.A(G218gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G211gat), .ZN(new_n296_));
  INV_X1    g095(.A(G211gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G218gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT89), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n296_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n299_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n294_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n296_), .A2(new_n298_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT89), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(KEYINPUT90), .A3(new_n300_), .ZN(new_n306_));
  INV_X1    g105(.A(G204gat), .ZN(new_n307_));
  INV_X1    g106(.A(G197gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT86), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT86), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(G197gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n307_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT21), .ZN(new_n313_));
  NOR2_X1   g112(.A1(G197gat), .A2(G204gat), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n312_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n303_), .A2(new_n306_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT88), .ZN(new_n317_));
  AOI21_X1  g116(.A(G204gat), .B1(new_n309_), .B2(new_n311_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT87), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n313_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n319_), .B1(new_n308_), .B2(G204gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT86), .B(G197gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n321_), .B1(new_n322_), .B2(G204gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n317_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n313_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n305_), .A2(new_n300_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n320_), .A2(new_n317_), .A3(new_n323_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n316_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(KEYINPUT85), .ZN(new_n331_));
  INV_X1    g130(.A(G233gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(KEYINPUT84), .A2(G228gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(KEYINPUT84), .A2(G228gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n284_), .A2(KEYINPUT29), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n331_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n337_), .B1(new_n331_), .B2(new_n338_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G78gat), .B(G106gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n293_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT93), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n331_), .A2(new_n338_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n336_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n339_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n344_), .B1(new_n349_), .B2(KEYINPUT92), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT92), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n348_), .A2(new_n351_), .A3(new_n339_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n346_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT92), .B1(new_n340_), .B2(new_n341_), .ZN(new_n354_));
  AND4_X1   g153(.A1(new_n346_), .A2(new_n354_), .A3(new_n343_), .A4(new_n352_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n345_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT91), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n349_), .B2(new_n343_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n349_), .A2(new_n357_), .A3(new_n343_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n293_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n246_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n284_), .A2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n246_), .B(new_n271_), .C1(new_n283_), .C2(new_n280_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(KEYINPUT4), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n284_), .A2(new_n368_), .A3(new_n364_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n363_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G1gat), .B(G29gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(G85gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT0), .B(G57gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n363_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n376_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n377_));
  OR3_X1    g176(.A1(new_n370_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n375_), .B1(new_n370_), .B2(new_n377_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n309_), .A2(new_n311_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(new_n319_), .A3(new_n307_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT21), .ZN(new_n383_));
  INV_X1    g182(.A(new_n321_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n318_), .A2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT88), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n314_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n322_), .B2(new_n307_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n388_), .A2(new_n313_), .B1(new_n305_), .B2(new_n300_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n329_), .A3(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n303_), .A2(new_n306_), .A3(new_n315_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT22), .B(G169gat), .ZN(new_n393_));
  INV_X1    g192(.A(G176gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n217_), .A2(KEYINPUT97), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n217_), .A2(KEYINPUT97), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n395_), .A2(new_n208_), .A3(new_n396_), .A4(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n224_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT95), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n217_), .A2(KEYINPUT94), .A3(KEYINPUT24), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT94), .B1(new_n217_), .B2(KEYINPUT24), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n401_), .A2(new_n402_), .A3(new_n214_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n231_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n400_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT94), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n218_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n217_), .A2(KEYINPUT94), .A3(KEYINPUT24), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n215_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(KEYINPUT95), .A3(new_n231_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n399_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT96), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n398_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n409_), .A2(KEYINPUT95), .A3(new_n231_), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT95), .B1(new_n409_), .B2(new_n231_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n224_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n416_), .A2(KEYINPUT96), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n392_), .B1(new_n413_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT20), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n235_), .A2(new_n236_), .A3(new_n211_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n236_), .B1(new_n235_), .B2(new_n211_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n419_), .B1(new_n330_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G226gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT19), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n418_), .A2(new_n423_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n419_), .B1(new_n392_), .B2(new_n238_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n390_), .A2(new_n416_), .A3(new_n391_), .A4(new_n398_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n426_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT102), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n427_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n418_), .A2(new_n423_), .A3(KEYINPUT102), .A4(new_n426_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G8gat), .B(G36gat), .Z(new_n435_));
  XNOR2_X1  g234(.A(G64gat), .B(G92gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n440_), .A2(KEYINPUT32), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n434_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n398_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n443_), .B1(new_n416_), .B2(KEYINPUT96), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n411_), .A2(new_n412_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n330_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT99), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT99), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n444_), .A2(new_n330_), .A3(new_n448_), .A4(new_n445_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n428_), .A2(new_n426_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n418_), .A2(new_n423_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT98), .B1(new_n453_), .B2(new_n425_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT98), .ZN(new_n455_));
  AOI211_X1 g254(.A(new_n455_), .B(new_n426_), .C1(new_n418_), .C2(new_n423_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n452_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n441_), .B(KEYINPUT101), .Z(new_n458_));
  OAI211_X1 g257(.A(new_n380_), .B(new_n442_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n439_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n365_), .A2(new_n366_), .A3(new_n376_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n461_), .A2(new_n374_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n367_), .A2(new_n363_), .A3(new_n369_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT33), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n379_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n452_), .B(new_n440_), .C1(new_n454_), .C2(new_n456_), .ZN(new_n467_));
  OAI211_X1 g266(.A(KEYINPUT33), .B(new_n375_), .C1(new_n370_), .C2(new_n377_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n460_), .A2(new_n466_), .A3(new_n467_), .A4(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n459_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n362_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n356_), .A2(new_n361_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n380_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT27), .ZN(new_n474_));
  INV_X1    g273(.A(new_n467_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n444_), .A2(new_n445_), .B1(new_n391_), .B2(new_n390_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT20), .B1(new_n392_), .B2(new_n238_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n425_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n455_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n453_), .A2(KEYINPUT98), .A3(new_n425_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n440_), .B1(new_n481_), .B2(new_n452_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n474_), .B1(new_n475_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT103), .ZN(new_n484_));
  AND4_X1   g283(.A1(KEYINPUT102), .A2(new_n418_), .A3(new_n423_), .A4(new_n426_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n429_), .B(KEYINPUT20), .C1(new_n330_), .C2(new_n422_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n425_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT102), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n485_), .B1(new_n488_), .B2(new_n427_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n484_), .B1(new_n489_), .B2(new_n440_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n434_), .A2(KEYINPUT103), .A3(new_n439_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n490_), .A2(KEYINPUT27), .A3(new_n467_), .A4(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n472_), .A2(new_n473_), .A3(new_n483_), .A4(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n256_), .B1(new_n471_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n256_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(new_n380_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n492_), .A2(new_n483_), .A3(KEYINPUT104), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT104), .B1(new_n492_), .B2(new_n483_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n362_), .B(new_n497_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(KEYINPUT105), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT105), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT104), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n467_), .A2(KEYINPUT27), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT103), .B1(new_n434_), .B2(new_n439_), .ZN(new_n505_));
  AOI211_X1 g304(.A(new_n484_), .B(new_n440_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT27), .B1(new_n460_), .B2(new_n467_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n503_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n492_), .A2(new_n483_), .A3(KEYINPUT104), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n472_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n502_), .B1(new_n511_), .B2(new_n497_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n495_), .B1(new_n501_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514_));
  INV_X1    g313(.A(G1gat), .ZN(new_n515_));
  INV_X1    g314(.A(G8gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT14), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G1gat), .B(G8gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G29gat), .B(G36gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G43gat), .B(G50gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n520_), .B(new_n523_), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT76), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(G229gat), .A3(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n523_), .B(KEYINPUT15), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n520_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529_));
  INV_X1    g328(.A(new_n520_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n523_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n528_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n526_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G113gat), .B(G141gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT77), .ZN(new_n535_));
  XOR2_X1   g334(.A(G169gat), .B(G197gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n533_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n513_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n541_), .B(KEYINPUT6), .Z(new_n542_));
  OR3_X1    g341(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(G85gat), .ZN(new_n546_));
  INV_X1    g345(.A(G92gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G85gat), .A2(G92gat), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n548_), .A2(KEYINPUT66), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT66), .B1(new_n548_), .B2(new_n549_), .ZN(new_n551_));
  OAI22_X1  g350(.A1(new_n542_), .A2(new_n545_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT8), .ZN(new_n553_));
  INV_X1    g352(.A(G106gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT10), .B(G99gat), .Z(new_n555_));
  AOI21_X1  g354(.A(new_n542_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n557_));
  INV_X1    g356(.A(new_n549_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT65), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT9), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n548_), .B1(new_n561_), .B2(new_n549_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n556_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n553_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT35), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT71), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n565_), .A2(new_n523_), .B1(new_n566_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n564_), .A2(KEYINPUT69), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT69), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n553_), .A2(new_n574_), .A3(new_n563_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n527_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n572_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n571_), .A2(new_n566_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G190gat), .B(G218gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(KEYINPUT36), .ZN(new_n584_));
  INV_X1    g383(.A(new_n579_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n572_), .B(new_n585_), .C1(new_n576_), .C2(new_n577_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n580_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT72), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT72), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n580_), .A2(new_n589_), .A3(new_n584_), .A4(new_n586_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n580_), .A2(new_n586_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n583_), .B(KEYINPUT36), .Z(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(KEYINPUT73), .A3(KEYINPUT37), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT67), .B(G71gat), .ZN(new_n598_));
  INV_X1    g397(.A(G78gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G57gat), .B(G64gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT11), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n601_), .B(KEYINPUT11), .Z(new_n604_));
  OAI21_X1  g403(.A(new_n603_), .B1(new_n604_), .B2(new_n600_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n564_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT68), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n597_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n564_), .A2(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT68), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n608_), .B1(new_n606_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT12), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n609_), .B1(new_n606_), .B2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n573_), .A2(KEYINPUT12), .A3(new_n605_), .A4(new_n575_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(new_n597_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT5), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G176gat), .B(G204gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n618_), .B(new_n619_), .Z(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n620_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n611_), .A2(new_n615_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT13), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n621_), .A2(KEYINPUT13), .A3(new_n623_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT37), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n591_), .A2(new_n594_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT73), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n629_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n520_), .B(KEYINPUT74), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n633_), .B(new_n634_), .Z(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(new_n605_), .Z(new_n636_));
  XOR2_X1   g435(.A(G127gat), .B(G155gat), .Z(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G183gat), .B(G211gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(KEYINPUT17), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n636_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n641_), .A2(KEYINPUT17), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n636_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n596_), .A2(new_n628_), .A3(new_n632_), .A4(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n540_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n515_), .A3(new_n380_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT38), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n500_), .A2(KEYINPUT105), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n509_), .A2(new_n510_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n653_), .A2(new_n502_), .A3(new_n362_), .A4(new_n497_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n494_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n595_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n628_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n646_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n657_), .A2(new_n538_), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n656_), .A2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G1gat), .B1(new_n660_), .B2(new_n473_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n649_), .A2(new_n650_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n651_), .A2(new_n661_), .A3(new_n662_), .ZN(G1324gat));
  NOR4_X1   g462(.A1(new_n540_), .A2(G8gat), .A3(new_n653_), .A4(new_n647_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G8gat), .B1(new_n660_), .B2(new_n653_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT39), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n667_), .B(G8gat), .C1(new_n660_), .C2(new_n653_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n664_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n669_), .B(new_n670_), .Z(G1325gat));
  NAND3_X1  g470(.A1(new_n648_), .A2(new_n249_), .A3(new_n256_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT107), .Z(new_n673_));
  OAI21_X1  g472(.A(G15gat), .B1(new_n660_), .B2(new_n496_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT41), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(KEYINPUT41), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n673_), .A2(new_n675_), .A3(new_n676_), .ZN(G1326gat));
  OAI21_X1  g476(.A(G22gat), .B1(new_n660_), .B2(new_n362_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT42), .ZN(new_n679_));
  INV_X1    g478(.A(G22gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n648_), .A2(new_n680_), .A3(new_n472_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1327gat));
  NAND2_X1  g481(.A1(new_n595_), .A2(new_n658_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n540_), .A2(new_n657_), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n380_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n657_), .A2(new_n538_), .A3(new_n646_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT37), .B1(new_n595_), .B2(KEYINPUT73), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n630_), .A2(new_n631_), .A3(new_n629_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n687_), .B1(new_n513_), .B2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n655_), .A2(KEYINPUT43), .A3(new_n690_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n686_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n513_), .A2(new_n687_), .A3(new_n691_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT43), .B1(new_n655_), .B2(new_n690_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(KEYINPUT44), .A3(new_n686_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n696_), .A2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n380_), .A2(G29gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n685_), .B1(new_n701_), .B2(new_n702_), .ZN(G1328gat));
  XNOR2_X1  g502(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n704_));
  INV_X1    g503(.A(new_n653_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n696_), .A2(new_n705_), .A3(new_n700_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G36gat), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n683_), .A2(new_n657_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n653_), .A2(G36gat), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n513_), .A2(new_n539_), .A3(new_n708_), .A4(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n704_), .B1(new_n707_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n704_), .ZN(new_n715_));
  AOI211_X1 g514(.A(new_n712_), .B(new_n715_), .C1(new_n706_), .C2(G36gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1329gat));
  NAND4_X1  g516(.A1(new_n696_), .A2(G43gat), .A3(new_n256_), .A4(new_n700_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n684_), .A2(new_n256_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n240_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT47), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n718_), .A2(new_n723_), .A3(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1330gat));
  AOI21_X1  g524(.A(G50gat), .B1(new_n684_), .B2(new_n472_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n472_), .A2(G50gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n701_), .B2(new_n727_), .ZN(G1331gat));
  NOR2_X1   g527(.A1(new_n655_), .A2(new_n539_), .ZN(new_n729_));
  AND4_X1   g528(.A1(new_n657_), .A2(new_n729_), .A3(new_n646_), .A4(new_n690_), .ZN(new_n730_));
  INV_X1    g529(.A(G57gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n380_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n657_), .A2(new_n538_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n658_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n656_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n737_), .A2(new_n380_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n732_), .B1(new_n738_), .B2(new_n731_), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n730_), .A2(new_n740_), .A3(new_n705_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n737_), .A2(new_n705_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(G64gat), .ZN(new_n744_));
  AOI211_X1 g543(.A(KEYINPUT48), .B(new_n740_), .C1(new_n737_), .C2(new_n705_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1333gat));
  NOR2_X1   g545(.A1(new_n496_), .A2(G71gat), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT111), .Z(new_n748_));
  NAND2_X1  g547(.A1(new_n730_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n737_), .A2(new_n256_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n750_), .A2(G71gat), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n750_), .B2(G71gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(G1334gat));
  NAND3_X1  g553(.A1(new_n730_), .A2(new_n599_), .A3(new_n472_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n737_), .A2(new_n472_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(G78gat), .ZN(new_n758_));
  AOI211_X1 g557(.A(KEYINPUT50), .B(new_n599_), .C1(new_n737_), .C2(new_n472_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n683_), .A2(new_n628_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n729_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(new_n546_), .A3(new_n380_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n692_), .A2(new_n693_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n733_), .A2(new_n646_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n765_), .A2(new_n473_), .A3(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n768_), .B2(new_n546_), .ZN(G1336gat));
  OAI21_X1  g568(.A(new_n547_), .B1(new_n762_), .B2(new_n653_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT112), .Z(new_n771_));
  NOR2_X1   g570(.A1(new_n765_), .A2(new_n767_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n653_), .A2(new_n547_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n771_), .B1(new_n772_), .B2(new_n773_), .ZN(G1337gat));
  INV_X1    g573(.A(G99gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n772_), .B2(new_n256_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n763_), .A2(new_n256_), .A3(new_n555_), .ZN(new_n777_));
  OR3_X1    g576(.A1(new_n776_), .A2(KEYINPUT51), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT51), .B1(new_n776_), .B2(new_n777_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1338gat));
  NAND3_X1  g579(.A1(new_n763_), .A2(new_n554_), .A3(new_n472_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n699_), .A2(new_n472_), .A3(new_n766_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n554_), .B1(KEYINPUT113), .B2(KEYINPUT52), .ZN(new_n783_));
  NOR2_X1   g582(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n781_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n781_), .B(new_n788_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1339gat));
  AOI21_X1  g591(.A(new_n597_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n615_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n613_), .A2(new_n614_), .A3(KEYINPUT55), .A4(new_n597_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n620_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n797_), .A2(KEYINPUT56), .A3(new_n620_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n526_), .A2(new_n532_), .A3(new_n537_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n525_), .A2(new_n529_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n529_), .B1(new_n530_), .B2(new_n523_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n537_), .B1(new_n528_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n803_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n809_), .A2(new_n623_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n802_), .A2(KEYINPUT58), .A3(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT58), .B1(new_n802_), .B2(new_n810_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n801_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT56), .B1(new_n797_), .B2(new_n620_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n539_), .B(new_n623_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n624_), .A2(new_n809_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n595_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  OAI22_X1  g617(.A1(new_n812_), .A2(new_n813_), .B1(new_n818_), .B2(KEYINPUT57), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n818_), .A2(KEYINPUT57), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n658_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OR3_X1    g620(.A1(new_n647_), .A2(KEYINPUT54), .A3(new_n539_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT54), .B1(new_n647_), .B2(new_n539_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n821_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n511_), .A2(new_n380_), .A3(new_n256_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n827_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n825_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n821_), .A2(new_n824_), .B1(new_n827_), .B2(new_n826_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT59), .B1(new_n833_), .B2(new_n828_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(G113gat), .B1(new_n835_), .B2(new_n538_), .ZN(new_n836_));
  OR3_X1    g635(.A1(new_n830_), .A2(G113gat), .A3(new_n538_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1340gat));
  OAI21_X1  g637(.A(G120gat), .B1(new_n835_), .B2(new_n628_), .ZN(new_n839_));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n628_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(KEYINPUT60), .B2(new_n840_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n839_), .B1(new_n830_), .B2(new_n842_), .ZN(G1341gat));
  OAI21_X1  g642(.A(G127gat), .B1(new_n835_), .B2(new_n658_), .ZN(new_n844_));
  OR3_X1    g643(.A1(new_n830_), .A2(G127gat), .A3(new_n658_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1342gat));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n825_), .A2(new_n595_), .A3(new_n828_), .A4(new_n829_), .ZN(new_n848_));
  INV_X1    g647(.A(G134gat), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n848_), .A2(KEYINPUT116), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT116), .B1(new_n848_), .B2(new_n849_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT117), .B(G134gat), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n691_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n830_), .A2(new_n831_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n833_), .A2(KEYINPUT59), .A3(new_n828_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n847_), .B1(new_n852_), .B2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n691_), .B(new_n854_), .C1(new_n832_), .C2(new_n834_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n860_), .B(KEYINPUT118), .C1(new_n851_), .C2(new_n850_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1343gat));
  AOI21_X1  g661(.A(new_n256_), .B1(new_n821_), .B2(new_n824_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n863_), .A2(new_n380_), .A3(new_n472_), .A4(new_n653_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n538_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(new_n263_), .ZN(G1344gat));
  NOR2_X1   g665(.A1(new_n864_), .A2(new_n628_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(new_n264_), .ZN(G1345gat));
  NOR2_X1   g667(.A1(new_n864_), .A2(new_n658_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT61), .B(G155gat), .Z(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1346gat));
  OAI21_X1  g670(.A(G162gat), .B1(new_n864_), .B2(new_n690_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n630_), .A2(G162gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n864_), .B2(new_n873_), .ZN(G1347gat));
  NAND2_X1  g673(.A1(new_n825_), .A2(new_n362_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n705_), .A2(new_n497_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n393_), .A3(new_n539_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n876_), .A2(new_n538_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT119), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n825_), .A2(new_n880_), .A3(new_n362_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n881_), .A2(new_n882_), .A3(G169gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n881_), .B2(G169gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n878_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT120), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n878_), .B(new_n887_), .C1(new_n884_), .C2(new_n883_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1348gat));
  AOI21_X1  g688(.A(G176gat), .B1(new_n877_), .B2(new_n657_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n875_), .B(KEYINPUT121), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n876_), .A2(new_n394_), .A3(new_n628_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n891_), .B2(new_n892_), .ZN(G1349gat));
  NAND2_X1  g692(.A1(new_n225_), .A2(new_n227_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n877_), .A2(new_n894_), .A3(new_n646_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n891_), .A2(new_n705_), .A3(new_n497_), .A4(new_n646_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n205_), .ZN(G1350gat));
  INV_X1    g696(.A(new_n877_), .ZN(new_n898_));
  OAI21_X1  g697(.A(G190gat), .B1(new_n898_), .B2(new_n690_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n595_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(new_n900_), .ZN(G1351gat));
  NOR2_X1   g700(.A1(new_n362_), .A2(new_n380_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n863_), .A2(new_n902_), .A3(new_n705_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n904_), .B(new_n539_), .C1(KEYINPUT122), .C2(G197gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT122), .B(G197gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(new_n903_), .B2(new_n538_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1352gat));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n904_), .B(new_n657_), .C1(new_n909_), .C2(new_n307_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n307_), .B2(KEYINPUT123), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1353gat));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n658_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n904_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n904_), .B2(new_n914_), .ZN(new_n916_));
  OAI22_X1  g715(.A1(new_n915_), .A2(new_n916_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n904_), .A2(new_n914_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT125), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n904_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n919_), .A2(new_n920_), .A3(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n917_), .A2(new_n922_), .ZN(G1354gat));
  XOR2_X1   g722(.A(KEYINPUT126), .B(G218gat), .Z(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n903_), .B2(new_n630_), .ZN(new_n925_));
  OR2_X1    g724(.A1(new_n690_), .A2(new_n924_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n903_), .B2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT127), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n925_), .B(new_n929_), .C1(new_n903_), .C2(new_n926_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1355gat));
endmodule


