//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n955_, new_n956_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT72), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n202_), .A2(KEYINPUT72), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n202_), .A2(KEYINPUT72), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(new_n208_), .A3(new_n204_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G85gat), .ZN(new_n216_));
  INV_X1    g015(.A(G92gat), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n216_), .A2(new_n217_), .A3(KEYINPUT9), .ZN(new_n218_));
  XOR2_X1   g017(.A(G85gat), .B(G92gat), .Z(new_n219_));
  AOI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(KEYINPUT9), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT10), .B(G99gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n215_), .B(new_n220_), .C1(G106gat), .C2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT6), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT65), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT6), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n226_), .A2(new_n228_), .A3(new_n214_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n214_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n224_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n226_), .A2(new_n228_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n214_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n226_), .A2(new_n228_), .A3(new_n214_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(KEYINPUT66), .A3(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G99gat), .A2(G106gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT7), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n231_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n223_), .B1(new_n239_), .B2(new_n219_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n219_), .A2(new_n223_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n241_), .B1(new_n215_), .B2(new_n238_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n222_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n212_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n210_), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n245_), .B(new_n222_), .C1(new_n240_), .C2(new_n242_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G232gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT34), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT35), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n244_), .A2(new_n246_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(KEYINPUT35), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n253_), .B(KEYINPUT71), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n212_), .A2(new_n243_), .B1(new_n250_), .B2(new_n249_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n254_), .B1(new_n257_), .B2(new_n246_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G190gat), .B(G218gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(G134gat), .B(G162gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n263_), .A2(KEYINPUT36), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(KEYINPUT36), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n259_), .B(KEYINPUT74), .C1(new_n264_), .C2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n252_), .A2(new_n255_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n257_), .A2(new_n254_), .A3(new_n246_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(KEYINPUT74), .A3(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n266_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n270_), .B(new_n271_), .C1(KEYINPUT36), .C2(new_n263_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n267_), .A2(new_n272_), .A3(KEYINPUT37), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT37), .B1(new_n267_), .B2(new_n272_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G57gat), .B(G64gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n276_), .A2(new_n277_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT11), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n276_), .A2(new_n277_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT11), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(new_n278_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT67), .B(G71gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(G78gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n281_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G78gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n285_), .B(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n289_), .B(KEYINPUT11), .C1(new_n279_), .C2(new_n280_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n243_), .A2(new_n292_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n291_), .B(new_n222_), .C1(new_n240_), .C2(new_n242_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(KEYINPUT69), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G230gat), .A2(G233gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n295_), .B(new_n297_), .C1(KEYINPUT69), .C2(new_n293_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(KEYINPUT70), .A2(KEYINPUT12), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(KEYINPUT70), .A2(KEYINPUT12), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n243_), .A2(new_n292_), .A3(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n301_), .B1(new_n243_), .B2(new_n292_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n300_), .B(new_n296_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n298_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G120gat), .B(G148gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT5), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G176gat), .B(G204gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n309_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n298_), .A2(new_n304_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT13), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(KEYINPUT13), .A3(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G15gat), .B(G22gat), .ZN(new_n318_));
  INV_X1    g117(.A(G1gat), .ZN(new_n319_));
  INV_X1    g118(.A(G8gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT14), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G1gat), .B(G8gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G231gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n292_), .B(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G127gat), .B(G155gat), .Z(new_n328_));
  XNOR2_X1  g127(.A(G183gat), .B(G211gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n327_), .A2(KEYINPUT17), .A3(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n332_), .B(KEYINPUT17), .Z(new_n335_));
  OAI21_X1  g134(.A(new_n334_), .B1(new_n327_), .B2(new_n335_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n275_), .A2(new_n317_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT100), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n341_), .B(new_n342_), .C1(G183gat), .C2(G190gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT22), .ZN(new_n345_));
  INV_X1    g144(.A(G169gat), .ZN(new_n346_));
  INV_X1    g145(.A(G176gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n343_), .A2(new_n344_), .A3(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT26), .B(G190gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G183gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT25), .B(G183gat), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n350_), .B(new_n354_), .C1(new_n355_), .C2(new_n353_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT24), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n357_), .B1(G169gat), .B2(G176gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n361_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n357_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n341_), .A2(new_n342_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n349_), .B1(new_n363_), .B2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G71gat), .B(G99gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(G43gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n370_), .B(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G227gat), .A2(G233gat), .ZN(new_n374_));
  INV_X1    g173(.A(G15gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT30), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT31), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n373_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(new_n378_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n381_), .A2(KEYINPUT79), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(KEYINPUT79), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(G134gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G127gat), .ZN(new_n386_));
  INV_X1    g185(.A(G127gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G134gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G120gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G113gat), .ZN(new_n391_));
  INV_X1    g190(.A(G113gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G120gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n386_), .A2(new_n388_), .A3(new_n391_), .A4(new_n393_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n384_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n397_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n382_), .A2(new_n399_), .A3(new_n383_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n402_));
  INV_X1    g201(.A(G141gat), .ZN(new_n403_));
  INV_X1    g202(.A(G148gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G141gat), .A2(G148gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT2), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n405_), .A2(new_n408_), .A3(new_n409_), .A4(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G155gat), .A2(G162gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n412_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  OR2_X1    g215(.A1(G155gat), .A2(G162gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(KEYINPUT80), .A3(new_n413_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n411_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n403_), .A2(new_n404_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n413_), .A2(KEYINPUT1), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n417_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n413_), .A2(KEYINPUT1), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n406_), .B(new_n420_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT29), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n419_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT28), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT28), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n419_), .A2(new_n424_), .A3(new_n428_), .A4(new_n425_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G22gat), .B(G50gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n427_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(KEYINPUT84), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G218gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G211gat), .ZN(new_n437_));
  INV_X1    g236(.A(G211gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(G218gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(G197gat), .A2(G204gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(G197gat), .A2(G204gat), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n442_), .A2(new_n443_), .A3(KEYINPUT21), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT21), .ZN(new_n445_));
  OR2_X1    g244(.A1(G197gat), .A2(G204gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G197gat), .A2(G204gat), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n441_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT82), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n446_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT21), .B1(new_n442_), .B2(new_n443_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n440_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT82), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n446_), .A2(new_n456_), .A3(new_n447_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT83), .B1(new_n442_), .B2(new_n443_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(KEYINPUT21), .A4(new_n440_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n451_), .A2(new_n455_), .A3(new_n459_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n460_), .A2(KEYINPUT81), .B1(G228gat), .B2(G233gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n419_), .A2(new_n424_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT29), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n463_), .A3(new_n460_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G228gat), .A2(G233gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n459_), .B1(new_n454_), .B2(KEYINPUT82), .ZN(new_n466_));
  AOI211_X1 g265(.A(new_n450_), .B(new_n440_), .C1(new_n453_), .C2(new_n452_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT81), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n465_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n460_), .A2(new_n463_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n435_), .A2(new_n464_), .A3(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G78gat), .B(G106gat), .Z(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n433_), .A2(new_n434_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT84), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n427_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n431_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n477_), .B(new_n475_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n473_), .B1(new_n478_), .B2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n477_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n474_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n461_), .B(new_n471_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n435_), .A4(new_n481_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G226gat), .A2(G233gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT19), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n370_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n491_), .B1(new_n492_), .B2(new_n468_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n358_), .A2(KEYINPUT86), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G169gat), .A2(G176gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(KEYINPUT86), .A3(KEYINPUT24), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n366_), .B(new_n368_), .C1(new_n494_), .C2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G183gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT25), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT85), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n352_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n352_), .B2(new_n500_), .ZN(new_n503_));
  XOR2_X1   g302(.A(KEYINPUT26), .B(G190gat), .Z(new_n504_));
  NOR3_X1   g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT22), .B(G169gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n345_), .A2(G169gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n346_), .A2(KEYINPUT22), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT87), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(G176gat), .B1(new_n508_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n343_), .A2(new_n495_), .ZN(new_n513_));
  OAI22_X1  g312(.A1(new_n498_), .A2(new_n505_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT20), .B1(new_n460_), .B2(new_n514_), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n493_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT20), .B1(new_n460_), .B2(new_n370_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n460_), .A2(new_n514_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT88), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT88), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n460_), .A2(new_n514_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n517_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n516_), .B1(new_n522_), .B2(new_n491_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G8gat), .B(G36gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT18), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G64gat), .B(G92gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT32), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n462_), .A2(new_n399_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n419_), .A2(new_n397_), .A3(new_n424_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G225gat), .A2(G233gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT92), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT92), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n530_), .A2(new_n535_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G57gat), .B(G85gat), .Z(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT91), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G85gat), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT91), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n539_), .A2(new_n319_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n319_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(G29gat), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n544_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(G29gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n546_), .B(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n539_), .A2(new_n542_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(G1gat), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n552_), .B2(new_n543_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n548_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n530_), .A2(KEYINPUT4), .A3(new_n531_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n397_), .B1(new_n419_), .B2(new_n424_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT4), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n532_), .B(KEYINPUT89), .Z(new_n559_));
  NAND3_X1  g358(.A1(new_n555_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n537_), .A2(new_n554_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n554_), .B1(new_n537_), .B2(new_n560_), .ZN(new_n562_));
  OAI22_X1  g361(.A1(new_n523_), .A2(new_n529_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  AOI22_X1  g362(.A1(new_n515_), .A2(KEYINPUT95), .B1(new_n460_), .B2(new_n370_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT95), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n565_), .B(KEYINPUT20), .C1(new_n460_), .C2(new_n514_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n491_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT20), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n492_), .B2(new_n468_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n460_), .A2(new_n514_), .A3(new_n520_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n520_), .B1(new_n460_), .B2(new_n514_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n491_), .B(new_n569_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n529_), .B1(new_n567_), .B2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n563_), .B1(KEYINPUT96), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT96), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n576_), .B(new_n529_), .C1(new_n567_), .C2(new_n573_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n548_), .A2(new_n553_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n419_), .A2(new_n397_), .A3(new_n424_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(new_n556_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n559_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n555_), .A2(new_n558_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n582_), .B1(new_n583_), .B2(new_n532_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n535_), .B1(new_n580_), .B2(new_n532_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n536_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n554_), .B(new_n560_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT93), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n584_), .B1(new_n588_), .B2(KEYINPUT33), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n493_), .A2(new_n515_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n569_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n591_), .B2(new_n490_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n527_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n527_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n523_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT33), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n587_), .A2(KEYINPUT93), .A3(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n589_), .A2(new_n593_), .A3(new_n595_), .A4(new_n597_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n575_), .A2(new_n577_), .B1(new_n598_), .B2(KEYINPUT94), .ZN(new_n599_));
  AOI211_X1 g398(.A(new_n594_), .B(new_n590_), .C1(new_n490_), .C2(new_n591_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n591_), .A2(new_n490_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n527_), .B1(new_n601_), .B2(new_n516_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT94), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n597_), .A4(new_n589_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n488_), .B1(new_n599_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n595_), .A2(new_n593_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT27), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n527_), .B(KEYINPUT98), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n609_), .B1(new_n567_), .B2(new_n573_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n608_), .B1(new_n592_), .B2(new_n527_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n607_), .A2(new_n608_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n613_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n537_), .A2(new_n560_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n578_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(KEYINPUT97), .A3(new_n587_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n612_), .A2(KEYINPUT99), .A3(new_n488_), .A4(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT99), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n608_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n611_), .A2(new_n610_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n488_), .A2(new_n617_), .A3(new_n614_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n621_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n620_), .A2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n401_), .B1(new_n606_), .B2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n483_), .A2(new_n487_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n612_), .A2(new_n629_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n401_), .A2(new_n630_), .A3(new_n618_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n628_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n210_), .B(new_n324_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(G229gat), .A3(G233gat), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n212_), .A2(new_n324_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(G229gat), .A2(G233gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT76), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n638_), .B1(new_n210_), .B2(new_n324_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n636_), .B2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G113gat), .B(G141gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G169gat), .B(G197gat), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n641_), .B(new_n642_), .Z(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n640_), .B(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n338_), .B1(new_n633_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n645_), .ZN(new_n647_));
  AOI211_X1 g446(.A(KEYINPUT100), .B(new_n647_), .C1(new_n628_), .C2(new_n632_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n337_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n598_), .A2(KEYINPUT94), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n574_), .A2(KEYINPUT96), .ZN(new_n653_));
  AOI22_X1  g452(.A1(new_n587_), .A2(new_n616_), .B1(new_n592_), .B2(new_n528_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n577_), .A3(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n652_), .A2(new_n605_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n629_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n626_), .A3(new_n620_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n631_), .B1(new_n658_), .B2(new_n401_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT100), .B1(new_n659_), .B2(new_n647_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n633_), .A2(new_n338_), .A3(new_n645_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(KEYINPUT101), .A3(new_n337_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n619_), .A2(G1gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n651_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT38), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n317_), .A2(new_n647_), .A3(new_n336_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT102), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n267_), .A2(new_n272_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n659_), .A2(new_n672_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n669_), .A2(new_n673_), .A3(KEYINPUT104), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT104), .B1(new_n669_), .B2(new_n673_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G1gat), .B1(new_n676_), .B2(new_n619_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n651_), .A2(KEYINPUT38), .A3(new_n663_), .A4(new_n664_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n667_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT105), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n667_), .A2(new_n677_), .A3(new_n681_), .A4(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(G1324gat));
  NAND3_X1  g482(.A1(new_n669_), .A2(new_n673_), .A3(new_n624_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT39), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT106), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n684_), .A2(G8gat), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n684_), .B2(G8gat), .ZN(new_n688_));
  OAI22_X1  g487(.A1(new_n687_), .A2(new_n688_), .B1(KEYINPUT106), .B2(new_n685_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n651_), .A2(new_n320_), .A3(new_n663_), .A4(new_n624_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(G1325gat));
  OAI21_X1  g492(.A(G15gat), .B1(new_n676_), .B2(new_n401_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n694_), .A2(KEYINPUT41), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(KEYINPUT41), .ZN(new_n696_));
  INV_X1    g495(.A(new_n401_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n662_), .A2(new_n375_), .A3(new_n697_), .A4(new_n337_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n698_), .A2(KEYINPUT108), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(KEYINPUT108), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n695_), .A2(new_n696_), .A3(new_n699_), .A4(new_n700_), .ZN(G1326gat));
  OR3_X1    g500(.A1(new_n649_), .A2(G22gat), .A3(new_n629_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G22gat), .B1(new_n676_), .B2(new_n629_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(KEYINPUT42), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(KEYINPUT42), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n702_), .B1(new_n704_), .B2(new_n705_), .ZN(G1327gat));
  NAND2_X1  g505(.A1(new_n670_), .A2(new_n336_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n709_), .A2(new_n317_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G29gat), .B1(new_n711_), .B2(new_n618_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n315_), .A2(new_n316_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n645_), .A3(new_n336_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT37), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n670_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n267_), .A2(new_n272_), .A3(KEYINPUT37), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n275_), .B2(new_n721_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n659_), .A2(new_n719_), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n719_), .B2(KEYINPUT109), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n633_), .B2(new_n275_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n715_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT110), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n722_), .B1(new_n659_), .B2(new_n719_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n633_), .A2(new_n275_), .A3(new_n724_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n714_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n727_), .A2(new_n728_), .A3(new_n733_), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n549_), .B(new_n619_), .C1(new_n731_), .C2(KEYINPUT44), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n712_), .B1(new_n734_), .B2(new_n735_), .ZN(G1328gat));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739_));
  INV_X1    g538(.A(new_n710_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n612_), .A2(G36gat), .ZN(new_n741_));
  AND4_X1   g540(.A1(new_n739_), .A2(new_n662_), .A3(new_n740_), .A4(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n739_), .B1(new_n711_), .B2(new_n741_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n738_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n662_), .A2(new_n740_), .A3(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT112), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n711_), .A2(new_n739_), .A3(new_n741_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(KEYINPUT45), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n744_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(G36gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n612_), .B1(new_n731_), .B2(KEYINPUT44), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n734_), .B2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n737_), .B1(new_n749_), .B2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n754_));
  AOI211_X1 g553(.A(KEYINPUT110), .B(new_n714_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(G36gat), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n757_), .A2(KEYINPUT46), .A3(new_n748_), .A4(new_n744_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n753_), .A2(new_n758_), .ZN(G1329gat));
  NAND2_X1  g558(.A1(new_n731_), .A2(KEYINPUT44), .ZN(new_n760_));
  INV_X1    g559(.A(G43gat), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n401_), .A2(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n760_), .B(new_n762_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n711_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n764_), .B2(new_n401_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n763_), .A2(KEYINPUT47), .A3(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT47), .B1(new_n763_), .B2(new_n765_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1330gat));
  AND3_X1   g567(.A1(new_n734_), .A2(new_n760_), .A3(new_n488_), .ZN(new_n769_));
  INV_X1    g568(.A(G50gat), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n488_), .A2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT113), .ZN(new_n772_));
  OAI22_X1  g571(.A1(new_n769_), .A2(new_n770_), .B1(new_n764_), .B2(new_n772_), .ZN(G1331gat));
  NAND2_X1  g572(.A1(new_n317_), .A2(new_n647_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n774_), .A2(new_n336_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n673_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(G57gat), .A3(new_n618_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT115), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n659_), .A2(KEYINPUT114), .A3(new_n645_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n633_), .B2(new_n647_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n336_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n719_), .A2(new_n317_), .A3(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G57gat), .B1(new_n786_), .B2(new_n618_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n779_), .A2(new_n787_), .ZN(G1332gat));
  INV_X1    g587(.A(G64gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n789_), .A3(new_n624_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT48), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n777_), .A2(new_n624_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(G64gat), .ZN(new_n793_));
  AOI211_X1 g592(.A(KEYINPUT48), .B(new_n789_), .C1(new_n777_), .C2(new_n624_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT116), .ZN(G1333gat));
  OAI21_X1  g595(.A(G71gat), .B1(new_n776_), .B2(new_n401_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT49), .ZN(new_n798_));
  INV_X1    g597(.A(G71gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n786_), .A2(new_n799_), .A3(new_n697_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1334gat));
  NAND2_X1  g600(.A1(new_n777_), .A2(new_n488_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(G78gat), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT117), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(new_n805_), .A3(G78gat), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n786_), .A2(new_n288_), .A3(new_n488_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n804_), .A2(KEYINPUT50), .A3(new_n806_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(G1335gat));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n774_), .A2(new_n784_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n729_), .A2(KEYINPUT118), .A3(new_n730_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n814_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(G85gat), .B1(new_n817_), .B2(new_n619_), .ZN(new_n818_));
  OR3_X1    g617(.A1(new_n783_), .A2(new_n713_), .A3(new_n709_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n618_), .A2(new_n216_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n818_), .B1(new_n819_), .B2(new_n820_), .ZN(G1336gat));
  OAI21_X1  g620(.A(G92gat), .B1(new_n817_), .B2(new_n612_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n624_), .A2(new_n217_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n819_), .B2(new_n823_), .ZN(G1337gat));
  NAND4_X1  g623(.A1(new_n814_), .A2(new_n697_), .A3(new_n815_), .A4(new_n816_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G99gat), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n401_), .A2(new_n221_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n819_), .B2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g628(.A(new_n488_), .B(new_n815_), .C1(new_n723_), .C2(new_n725_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n830_), .A2(new_n831_), .A3(G106gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n830_), .B2(G106gat), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n629_), .A2(G106gat), .ZN(new_n834_));
  OAI22_X1  g633(.A1(new_n832_), .A2(new_n833_), .B1(new_n819_), .B2(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g635(.A1(new_n401_), .A2(new_n630_), .A3(new_n619_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n645_), .A2(new_n312_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n294_), .A2(new_n299_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n301_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n293_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n243_), .A2(new_n292_), .A3(new_n301_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n841_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT55), .B1(new_n845_), .B2(new_n296_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n304_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(KEYINPUT55), .A3(new_n296_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT56), .B1(new_n849_), .B2(new_n309_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n851_), .B(new_n311_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n840_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n640_), .A2(new_n644_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n210_), .A2(new_n324_), .ZN(new_n855_));
  OR3_X1    g654(.A1(new_n636_), .A2(new_n855_), .A3(new_n638_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n643_), .B1(new_n634_), .B2(new_n638_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n854_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n313_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n670_), .B1(new_n853_), .B2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n858_), .A2(new_n312_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n862_), .B(new_n863_), .C1(new_n850_), .C2(new_n852_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n275_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n300_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n297_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n304_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n848_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n309_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n851_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n849_), .A2(KEYINPUT56), .A3(new_n309_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n862_), .B1(new_n875_), .B2(new_n863_), .ZN(new_n876_));
  OAI22_X1  g675(.A1(new_n860_), .A2(KEYINPUT57), .B1(new_n865_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n670_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n839_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n859_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n336_), .B1(new_n877_), .B2(new_n883_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n719_), .A2(new_n647_), .A3(new_n713_), .A4(new_n784_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT54), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n838_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(G113gat), .B1(new_n887_), .B2(new_n645_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n885_), .B(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n860_), .A2(KEYINPUT57), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n881_), .A2(new_n882_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n891_), .B(new_n892_), .C1(new_n876_), .C2(new_n865_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n890_), .B1(new_n893_), .B2(new_n336_), .ZN(new_n894_));
  AOI21_X1  g693(.A(KEYINPUT59), .B1(new_n837_), .B2(KEYINPUT121), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(KEYINPUT121), .B2(new_n837_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT120), .B1(new_n887_), .B2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n900_), .B(KEYINPUT59), .C1(new_n894_), .C2(new_n838_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n897_), .B1(new_n899_), .B2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n647_), .A2(new_n392_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n888_), .B1(new_n902_), .B2(new_n903_), .ZN(G1340gat));
  OAI21_X1  g703(.A(new_n390_), .B1(new_n713_), .B2(KEYINPUT60), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n887_), .B(new_n905_), .C1(KEYINPUT60), .C2(new_n390_), .ZN(new_n906_));
  AOI211_X1 g705(.A(new_n713_), .B(new_n897_), .C1(new_n899_), .C2(new_n901_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n390_), .ZN(G1341gat));
  INV_X1    g707(.A(new_n887_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n387_), .B1(new_n909_), .B2(new_n336_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT122), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n912_), .B(new_n387_), .C1(new_n909_), .C2(new_n336_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n336_), .A2(new_n387_), .ZN(new_n914_));
  AOI22_X1  g713(.A1(new_n911_), .A2(new_n913_), .B1(new_n902_), .B2(new_n914_), .ZN(G1342gat));
  AOI21_X1  g714(.A(G134gat), .B1(new_n887_), .B2(new_n672_), .ZN(new_n916_));
  XOR2_X1   g715(.A(KEYINPUT123), .B(G134gat), .Z(new_n917_));
  NOR2_X1   g716(.A1(new_n719_), .A2(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n902_), .B2(new_n918_), .ZN(G1343gat));
  NAND2_X1  g718(.A1(new_n884_), .A2(new_n886_), .ZN(new_n920_));
  NOR4_X1   g719(.A1(new_n697_), .A2(new_n629_), .A3(new_n624_), .A4(new_n619_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n647_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(new_n403_), .ZN(G1344gat));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n713_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n404_), .ZN(G1345gat));
  AND2_X1   g725(.A1(new_n920_), .A2(new_n921_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n927_), .A2(new_n928_), .A3(new_n784_), .ZN(new_n929_));
  OAI21_X1  g728(.A(KEYINPUT124), .B1(new_n922_), .B2(new_n336_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT61), .B(G155gat), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n933_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n929_), .A2(new_n930_), .A3(new_n932_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1346gat));
  AOI21_X1  g735(.A(G162gat), .B1(new_n927_), .B2(new_n672_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n275_), .A2(G162gat), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(KEYINPUT125), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n927_), .B2(new_n939_), .ZN(G1347gat));
  XOR2_X1   g739(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n941_));
  NOR3_X1   g740(.A1(new_n401_), .A2(new_n612_), .A3(new_n618_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(KEYINPUT126), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n943_), .A2(new_n488_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n920_), .A2(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n647_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n941_), .B1(new_n946_), .B2(new_n346_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n508_), .A2(new_n511_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n948_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n941_), .ZN(new_n950_));
  OAI211_X1 g749(.A(G169gat), .B(new_n950_), .C1(new_n945_), .C2(new_n647_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n947_), .A2(new_n949_), .A3(new_n951_), .ZN(G1348gat));
  NOR2_X1   g751(.A1(new_n945_), .A2(new_n713_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(new_n347_), .ZN(G1349gat));
  NOR2_X1   g753(.A1(new_n502_), .A2(new_n503_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n945_), .A2(new_n336_), .ZN(new_n956_));
  MUX2_X1   g755(.A(G183gat), .B(new_n955_), .S(new_n956_), .Z(G1350gat));
  OAI21_X1  g756(.A(G190gat), .B1(new_n945_), .B2(new_n719_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n672_), .A2(new_n350_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n945_), .B2(new_n959_), .ZN(G1351gat));
  NOR3_X1   g759(.A1(new_n697_), .A2(new_n612_), .A3(new_n625_), .ZN(new_n961_));
  AND2_X1   g760(.A1(new_n920_), .A2(new_n961_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(new_n645_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g763(.A1(new_n962_), .A2(new_n317_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g765(.A1(new_n962_), .A2(new_n784_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(KEYINPUT63), .B(G211gat), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n967_), .A2(new_n968_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n969_), .B1(new_n967_), .B2(new_n970_), .ZN(G1354gat));
  NAND3_X1  g770(.A1(new_n962_), .A2(new_n436_), .A3(new_n672_), .ZN(new_n972_));
  AND2_X1   g771(.A1(new_n962_), .A2(new_n275_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n972_), .B1(new_n973_), .B2(new_n436_), .ZN(G1355gat));
endmodule


