//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n597_, new_n598_, new_n599_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT74), .B(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT75), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT75), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n209_), .A3(new_n206_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G1gat), .B(G8gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n208_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G29gat), .B(G36gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n214_), .A2(new_n215_), .A3(new_n219_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT77), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n221_), .A2(KEYINPUT77), .A3(new_n222_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n202_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n228_));
  XNOR2_X1  g027(.A(new_n219_), .B(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n216_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(new_n222_), .A3(new_n202_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G113gat), .B(G141gat), .Z(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT78), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G169gat), .B(G197gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n234_), .B(new_n235_), .Z(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n227_), .A2(new_n232_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n237_), .B1(new_n227_), .B2(new_n232_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(KEYINPUT79), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT79), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n242_), .B(new_n237_), .C1(new_n227_), .C2(new_n232_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G225gat), .A2(G233gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G141gat), .A2(G148gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT86), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT2), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(G141gat), .A2(G148gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT3), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n250_), .B(new_n252_), .C1(new_n249_), .C2(new_n247_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G155gat), .B(G162gat), .Z(new_n254_));
  AND2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n248_), .B(new_n256_), .C1(G141gat), .C2(G148gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(new_n254_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G127gat), .B(G134gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT85), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G113gat), .B(G120gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n246_), .B1(new_n267_), .B2(KEYINPUT4), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT92), .B1(new_n260_), .B2(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n261_), .A2(KEYINPUT92), .A3(new_n266_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n268_), .B1(new_n272_), .B2(KEYINPUT4), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT93), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n276_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT93), .B1(new_n277_), .B2(new_n268_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n272_), .A2(new_n245_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G1gat), .B(G29gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(G85gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT0), .B(G57gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n282_), .B(new_n283_), .Z(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n285_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n275_), .A2(new_n284_), .A3(new_n278_), .A4(new_n279_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G183gat), .ZN(new_n289_));
  INV_X1    g088(.A(G190gat), .ZN(new_n290_));
  OR3_X1    g089(.A1(new_n289_), .A2(new_n290_), .A3(KEYINPUT23), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT23), .B1(new_n289_), .B2(new_n290_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT80), .B(G183gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(G190gat), .B2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(KEYINPUT84), .B(G176gat), .Z(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT22), .B(G169gat), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n297_), .A2(new_n298_), .B1(G169gat), .B2(G176gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(KEYINPUT26), .B(G190gat), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n294_), .A2(KEYINPUT25), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT81), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT25), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(KEYINPUT82), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n289_), .B1(KEYINPUT82), .B2(new_n304_), .ZN(new_n306_));
  AOI211_X1 g105(.A(new_n301_), .B(new_n303_), .C1(new_n305_), .C2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n292_), .B(KEYINPUT83), .Z(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n291_), .ZN(new_n309_));
  INV_X1    g108(.A(G169gat), .ZN(new_n310_));
  INV_X1    g109(.A(G176gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT24), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313_));
  MUX2_X1   g112(.A(new_n312_), .B(KEYINPUT24), .S(new_n313_), .Z(new_n314_));
  NAND2_X1  g113(.A1(new_n309_), .A2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n300_), .B1(new_n307_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT21), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G197gat), .B(G204gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT89), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G211gat), .B(G218gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n320_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n318_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n317_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT21), .B1(new_n319_), .B2(new_n320_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n316_), .A2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n309_), .B1(G183gat), .B2(G190gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n299_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT25), .B(G183gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n314_), .B(new_n293_), .C1(new_n301_), .C2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n333_), .A2(new_n326_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n327_), .A2(new_n334_), .A3(KEYINPUT20), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT19), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n316_), .A2(new_n326_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT20), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n333_), .B2(new_n326_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n337_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G8gat), .B(G36gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT18), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT32), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n338_), .A2(new_n343_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n335_), .A2(new_n337_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n350_), .B1(new_n337_), .B2(new_n342_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n348_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n349_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n288_), .A2(new_n353_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n338_), .A2(new_n343_), .A3(new_n347_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n347_), .B1(new_n338_), .B2(new_n343_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT33), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n287_), .A2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n284_), .B1(new_n272_), .B2(new_n246_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n245_), .B1(new_n267_), .B2(KEYINPUT4), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n360_), .B1(new_n277_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT94), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT94), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n360_), .B(new_n364_), .C1(new_n277_), .C2(new_n361_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n273_), .A2(new_n274_), .B1(new_n272_), .B2(new_n245_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n367_), .A2(KEYINPUT33), .A3(new_n284_), .A4(new_n278_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n357_), .A2(new_n359_), .A3(new_n366_), .A4(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n354_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT91), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n260_), .A2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n375_), .B(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G22gat), .B(G50gat), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n375_), .B(new_n376_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(new_n379_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n373_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n379_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n378_), .A2(new_n380_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n371_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n326_), .B1(new_n260_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT88), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(G228gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(G228gat), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n392_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n391_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n397_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n399_), .B(new_n326_), .C1(new_n260_), .C2(new_n374_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n389_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n384_), .A2(new_n401_), .A3(new_n388_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G71gat), .B(G99gat), .ZN(new_n406_));
  INV_X1    g205(.A(G43gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n316_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n408_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n410_), .B(new_n300_), .C1(new_n307_), .C2(new_n315_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n266_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414_));
  INV_X1    g213(.A(G15gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT30), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT31), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n266_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n420_));
  OR3_X1    g219(.A1(new_n413_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n413_), .B2(new_n420_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n405_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n370_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n338_), .A2(new_n343_), .A3(new_n347_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT27), .ZN(new_n427_));
  INV_X1    g226(.A(new_n347_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n428_), .B2(new_n351_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n356_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT27), .B1(new_n430_), .B2(new_n426_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n423_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n384_), .A2(new_n401_), .A3(new_n388_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n401_), .B1(new_n384_), .B2(new_n388_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n403_), .A2(new_n404_), .A3(new_n423_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n288_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n432_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n244_), .B1(new_n425_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G230gat), .A2(G233gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT10), .B(G99gat), .Z(new_n444_));
  INV_X1    g243(.A(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(G85gat), .ZN(new_n447_));
  INV_X1    g246(.A(G92gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G85gat), .A2(G92gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(KEYINPUT9), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n446_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n450_), .A2(KEYINPUT9), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n452_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT7), .ZN(new_n458_));
  INV_X1    g257(.A(G99gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n445_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n456_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n450_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT64), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT64), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n449_), .A2(new_n467_), .A3(new_n450_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n463_), .A2(KEYINPUT8), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n455_), .A2(KEYINPUT65), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT65), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT6), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n471_), .A2(new_n473_), .A3(new_n454_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n454_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n462_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT8), .B1(new_n476_), .B2(new_n469_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n470_), .B1(new_n477_), .B2(KEYINPUT66), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT8), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n460_), .A2(new_n461_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n454_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n472_), .A2(KEYINPUT6), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n455_), .A2(KEYINPUT65), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n471_), .A2(new_n473_), .A3(new_n454_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n480_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n466_), .A2(new_n468_), .ZN(new_n487_));
  AOI211_X1 g286(.A(KEYINPUT66), .B(new_n479_), .C1(new_n486_), .C2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n457_), .B1(new_n478_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G57gat), .B(G64gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT11), .ZN(new_n492_));
  XOR2_X1   g291(.A(G71gat), .B(G78gat), .Z(new_n493_));
  OR2_X1    g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n491_), .A2(KEYINPUT11), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n493_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n490_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n490_), .A2(new_n497_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n443_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n457_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n487_), .B(new_n479_), .C1(new_n456_), .C2(new_n462_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n479_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT66), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n502_), .B1(new_n506_), .B2(new_n488_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT67), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(KEYINPUT67), .B(new_n502_), .C1(new_n506_), .C2(new_n488_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT12), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n497_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(new_n510_), .A3(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n511_), .B1(new_n490_), .B2(new_n497_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n443_), .B1(new_n490_), .B2(new_n497_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n501_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G120gat), .B(G148gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G176gat), .B(G204gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT69), .B1(new_n518_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT69), .ZN(new_n525_));
  INV_X1    g324(.A(new_n523_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n501_), .A2(new_n517_), .A3(new_n525_), .A4(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n518_), .A2(new_n523_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT13), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n528_), .A2(KEYINPUT13), .A3(new_n529_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT37), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G232gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT35), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n540_), .A2(KEYINPUT72), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n509_), .A2(new_n229_), .A3(new_n510_), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n490_), .A2(new_n219_), .B1(new_n539_), .B2(new_n538_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(KEYINPUT72), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT73), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n542_), .A2(KEYINPUT72), .A3(new_n543_), .A4(new_n540_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G190gat), .B(G218gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT36), .Z(new_n552_));
  NAND4_X1  g351(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .A4(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n546_), .A2(new_n548_), .A3(new_n552_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT73), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n551_), .A2(KEYINPUT36), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n535_), .B(new_n553_), .C1(new_n555_), .C2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n497_), .B(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(new_n216_), .Z(new_n562_));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G127gat), .B(G155gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT16), .ZN(new_n565_));
  XOR2_X1   g364(.A(G183gat), .B(G211gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n562_), .B1(new_n563_), .B2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(KEYINPUT17), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n568_), .B1(new_n562_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT76), .ZN(new_n571_));
  INV_X1    g370(.A(new_n558_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(KEYINPUT37), .A3(new_n554_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n559_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n534_), .A2(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n441_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(new_n203_), .A3(new_n288_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT38), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n553_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n580_), .B1(new_n425_), .B2(new_n440_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n534_), .A2(new_n244_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n581_), .A2(new_n571_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(G1gat), .B1(new_n584_), .B2(new_n439_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n577_), .A2(new_n578_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(new_n585_), .A3(new_n586_), .ZN(G1324gat));
  INV_X1    g386(.A(new_n432_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n576_), .A2(new_n204_), .A3(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(G8gat), .B1(new_n584_), .B2(new_n432_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n590_), .A2(KEYINPUT39), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(KEYINPUT39), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n589_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT95), .B(KEYINPUT40), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n593_), .B(new_n595_), .ZN(G1325gat));
  AOI21_X1  g395(.A(new_n415_), .B1(new_n583_), .B2(new_n423_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT41), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n576_), .A2(new_n415_), .A3(new_n423_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(G1326gat));
  INV_X1    g399(.A(G22gat), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n576_), .A2(new_n601_), .A3(new_n405_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n405_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G22gat), .B1(new_n584_), .B2(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n604_), .A2(KEYINPUT42), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(KEYINPUT42), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n602_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT96), .ZN(G1327gat));
  INV_X1    g407(.A(new_n534_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n580_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n571_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n441_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n612_));
  OR3_X1    g411(.A1(new_n612_), .A2(G29gat), .A3(new_n439_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n534_), .A2(new_n244_), .A3(new_n571_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT43), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n425_), .A2(new_n440_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n559_), .A2(new_n573_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n615_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n617_), .ZN(new_n619_));
  AOI211_X1 g418(.A(KEYINPUT43), .B(new_n619_), .C1(new_n425_), .C2(new_n440_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n614_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT44), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(KEYINPUT44), .B(new_n614_), .C1(new_n618_), .C2(new_n620_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(new_n288_), .A3(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(KEYINPUT97), .ZN(new_n626_));
  OAI21_X1  g425(.A(G29gat), .B1(new_n625_), .B2(KEYINPUT97), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n613_), .B1(new_n626_), .B2(new_n627_), .ZN(G1328gat));
  NOR2_X1   g427(.A1(new_n432_), .A2(G36gat), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n441_), .A2(new_n609_), .A3(new_n611_), .A4(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT45), .Z(new_n631_));
  NAND3_X1  g430(.A1(new_n623_), .A2(new_n588_), .A3(new_n624_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n632_), .B2(G36gat), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT46), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n633_), .A2(KEYINPUT98), .A3(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n634_), .A2(KEYINPUT98), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n634_), .A2(KEYINPUT98), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n633_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n635_), .A2(new_n638_), .ZN(G1329gat));
  NOR3_X1   g438(.A1(new_n612_), .A2(G43gat), .A3(new_n433_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n623_), .A2(new_n423_), .A3(new_n624_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n641_), .B2(G43gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g442(.A1(new_n623_), .A2(G50gat), .A3(new_n405_), .A4(new_n624_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n612_), .A2(new_n603_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(G50gat), .B2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT99), .Z(G1331gat));
  INV_X1    g446(.A(new_n244_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n609_), .A2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n616_), .A2(new_n649_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n650_), .A2(new_n571_), .A3(new_n619_), .ZN(new_n651_));
  INV_X1    g450(.A(G57gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(new_n652_), .A3(new_n288_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n581_), .A2(new_n571_), .A3(new_n649_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(new_n288_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n653_), .B1(new_n655_), .B2(new_n652_), .ZN(G1332gat));
  INV_X1    g455(.A(G64gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n654_), .B2(new_n588_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT48), .Z(new_n659_));
  NAND3_X1  g458(.A1(new_n651_), .A2(new_n657_), .A3(new_n588_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1333gat));
  INV_X1    g460(.A(G71gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n651_), .A2(new_n662_), .A3(new_n423_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n654_), .A2(new_n423_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G71gat), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n665_), .A2(KEYINPUT101), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(KEYINPUT101), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT100), .B(KEYINPUT49), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n663_), .B1(new_n669_), .B2(new_n670_), .ZN(G1334gat));
  INV_X1    g470(.A(G78gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n654_), .B2(new_n405_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT50), .Z(new_n674_));
  NAND3_X1  g473(.A1(new_n651_), .A2(new_n672_), .A3(new_n405_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1335gat));
  NOR2_X1   g475(.A1(new_n618_), .A2(new_n620_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n571_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n649_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n288_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n650_), .A2(new_n611_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n439_), .A2(G85gat), .ZN(new_n683_));
  AOI22_X1  g482(.A1(new_n681_), .A2(G85gat), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT102), .Z(G1336gat));
  NAND3_X1  g484(.A1(new_n682_), .A2(new_n448_), .A3(new_n588_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n680_), .A2(new_n588_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n688_), .B2(new_n448_), .ZN(G1337gat));
  AOI21_X1  g488(.A(new_n459_), .B1(new_n680_), .B2(new_n423_), .ZN(new_n690_));
  AND2_X1   g489(.A1(KEYINPUT103), .A2(KEYINPUT51), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n682_), .A2(new_n423_), .A3(new_n444_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n690_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(KEYINPUT103), .A2(KEYINPUT51), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT104), .Z(new_n695_));
  XNOR2_X1  g494(.A(new_n693_), .B(new_n695_), .ZN(G1338gat));
  NAND3_X1  g495(.A1(new_n682_), .A2(new_n445_), .A3(new_n405_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n679_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n405_), .B(new_n698_), .C1(new_n618_), .C2(new_n620_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT106), .B1(new_n699_), .B2(G106gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(KEYINPUT106), .A3(G106gat), .ZN(new_n701_));
  XOR2_X1   g500(.A(KEYINPUT105), .B(KEYINPUT52), .Z(new_n702_));
  AND3_X1   g501(.A1(new_n700_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n700_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n697_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT53), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT53), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n707_), .B(new_n697_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1339gat));
  INV_X1    g508(.A(KEYINPUT54), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n575_), .B2(new_n244_), .ZN(new_n711_));
  NOR4_X1   g510(.A1(new_n534_), .A2(new_n574_), .A3(new_n648_), .A4(KEYINPUT54), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT58), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT55), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n514_), .A2(new_n498_), .A3(new_n515_), .ZN(new_n716_));
  AOI22_X1  g515(.A1(new_n715_), .A2(new_n517_), .B1(new_n716_), .B2(new_n443_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n514_), .A2(KEYINPUT55), .A3(new_n515_), .A4(new_n516_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n718_), .A2(new_n719_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT56), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n526_), .A2(new_n723_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n722_), .A2(KEYINPUT111), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT56), .B1(new_n722_), .B2(new_n523_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT111), .B1(new_n722_), .B2(new_n724_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n230_), .A2(G229gat), .A3(G233gat), .A4(new_n222_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n237_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n225_), .A2(new_n226_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(new_n202_), .ZN(new_n732_));
  OR3_X1    g531(.A1(new_n238_), .A2(KEYINPUT109), .A3(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT109), .B1(new_n238_), .B2(new_n732_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n528_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n714_), .B1(new_n728_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n528_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n724_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n718_), .B(new_n719_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(new_n717_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n526_), .B1(new_n741_), .B2(new_n717_), .ZN(new_n743_));
  OAI22_X1  g542(.A1(KEYINPUT111), .A2(new_n742_), .B1(new_n743_), .B2(KEYINPUT56), .ZN(new_n744_));
  OAI211_X1 g543(.A(KEYINPUT58), .B(new_n739_), .C1(new_n744_), .C2(new_n725_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n737_), .A2(new_n617_), .A3(new_n745_), .ZN(new_n746_));
  XOR2_X1   g545(.A(KEYINPUT110), .B(KEYINPUT57), .Z(new_n747_));
  AOI22_X1  g546(.A1(new_n733_), .A2(new_n734_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n722_), .A2(new_n523_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n723_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n718_), .B(KEYINPUT107), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n517_), .A2(new_n715_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n716_), .A2(new_n443_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n724_), .B1(new_n751_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n722_), .A2(KEYINPUT108), .A3(new_n724_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n750_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n241_), .A2(new_n528_), .A3(new_n243_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n748_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n747_), .B1(new_n762_), .B2(new_n580_), .ZN(new_n763_));
  AOI22_X1  g562(.A1(new_n723_), .A2(new_n749_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n760_), .B1(new_n764_), .B2(new_n758_), .ZN(new_n765_));
  OAI211_X1 g564(.A(KEYINPUT57), .B(new_n610_), .C1(new_n765_), .C2(new_n748_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n746_), .A2(new_n763_), .A3(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n713_), .B1(new_n767_), .B2(new_n678_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n588_), .A2(new_n439_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n437_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  OR3_X1    g570(.A1(new_n768_), .A2(KEYINPUT112), .A3(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT112), .B1(new_n768_), .B2(new_n771_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n648_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(G113gat), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n774_), .A2(KEYINPUT113), .A3(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n767_), .A2(new_n678_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n713_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n782_), .A2(KEYINPUT114), .A3(new_n770_), .A4(new_n769_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT59), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n784_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n244_), .A2(new_n775_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n778_), .A2(new_n779_), .B1(new_n787_), .B2(new_n788_), .ZN(G1340gat));
  AND2_X1   g588(.A1(new_n772_), .A2(new_n773_), .ZN(new_n790_));
  INV_X1    g589(.A(G120gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n609_), .B2(KEYINPUT60), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT115), .B1(new_n791_), .B2(KEYINPUT60), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n790_), .B(new_n794_), .C1(new_n795_), .C2(new_n792_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n609_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n791_), .ZN(G1341gat));
  INV_X1    g597(.A(G127gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n790_), .A2(new_n799_), .A3(new_n571_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n678_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(new_n799_), .ZN(G1342gat));
  INV_X1    g601(.A(G134gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n790_), .A2(new_n803_), .A3(new_n580_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n619_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n803_), .ZN(G1343gat));
  INV_X1    g605(.A(new_n436_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n769_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n782_), .A2(KEYINPUT116), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n768_), .B2(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n648_), .ZN(new_n814_));
  XOR2_X1   g613(.A(KEYINPUT117), .B(G141gat), .Z(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(G1344gat));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n534_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(G148gat), .ZN(G1345gat));
  AOI21_X1  g617(.A(KEYINPUT118), .B1(new_n813_), .B2(new_n571_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n820_), .B(new_n678_), .C1(new_n810_), .C2(new_n812_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT61), .B(G155gat), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n819_), .A2(new_n821_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT116), .B1(new_n782_), .B2(new_n809_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n768_), .A2(new_n811_), .A3(new_n808_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n571_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n820_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n813_), .A2(KEYINPUT118), .A3(new_n571_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n822_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n824_), .A2(new_n830_), .ZN(G1346gat));
  INV_X1    g630(.A(G162gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n813_), .A2(new_n832_), .A3(new_n580_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n619_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT119), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n833_), .B(new_n837_), .C1(new_n832_), .C2(new_n834_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1347gat));
  NOR2_X1   g638(.A1(new_n432_), .A2(new_n288_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n648_), .A3(new_n423_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT120), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n405_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n310_), .B1(new_n843_), .B2(new_n782_), .ZN(new_n844_));
  XOR2_X1   g643(.A(new_n844_), .B(KEYINPUT62), .Z(new_n845_));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n840_), .A2(new_n603_), .A3(new_n423_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n782_), .A2(new_n846_), .A3(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT121), .B1(new_n768_), .B2(new_n847_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(new_n648_), .A3(new_n298_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n845_), .A2(new_n852_), .ZN(G1348gat));
  NOR2_X1   g652(.A1(new_n768_), .A2(new_n847_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(G176gat), .A3(new_n534_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n609_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n297_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1349gat));
  AOI21_X1  g659(.A(new_n295_), .B1(new_n854_), .B2(new_n571_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n678_), .A2(new_n330_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n851_), .B2(new_n862_), .ZN(G1350gat));
  NOR2_X1   g662(.A1(new_n610_), .A2(new_n301_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT124), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n851_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n851_), .A2(new_n617_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(G190gat), .ZN(new_n869_));
  AOI211_X1 g668(.A(KEYINPUT123), .B(new_n290_), .C1(new_n851_), .C2(new_n617_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n866_), .B1(new_n869_), .B2(new_n870_), .ZN(G1351gat));
  NAND4_X1  g670(.A1(new_n782_), .A2(KEYINPUT125), .A3(new_n807_), .A4(new_n840_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n840_), .A2(new_n807_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n768_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n648_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT126), .B(G197gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1352gat));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n534_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n876_), .A2(new_n571_), .A3(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n883_), .B(new_n884_), .Z(G1354gat));
  NOR2_X1   g684(.A1(new_n610_), .A2(G218gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n876_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(G218gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n619_), .B1(new_n872_), .B2(new_n875_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT127), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT127), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n887_), .B(new_n892_), .C1(new_n888_), .C2(new_n889_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1355gat));
endmodule


