//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G113gat), .B(G120gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(new_n202_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(G71gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G227gat), .A2(G233gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT82), .B(G99gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G15gat), .B(G43gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT31), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT83), .B(KEYINPUT30), .Z(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT80), .ZN(new_n218_));
  INV_X1    g017(.A(G169gat), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n223_), .A2(KEYINPUT81), .A3(KEYINPUT24), .A4(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n221_), .A2(new_n222_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT24), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT26), .B(G190gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT25), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G183gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n235_), .A2(KEYINPUT79), .A3(G183gat), .ZN(new_n239_));
  INV_X1    g038(.A(G183gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT25), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n234_), .A2(new_n238_), .A3(new_n239_), .A4(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n221_), .A2(KEYINPUT24), .A3(new_n224_), .A4(new_n222_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT81), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n225_), .A2(new_n233_), .A3(new_n242_), .A4(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT22), .B(G169gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n220_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n248_), .B(new_n224_), .C1(new_n230_), .C2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n217_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n213_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n213_), .A2(new_n253_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT93), .B(KEYINPUT0), .Z(new_n257_));
  XNOR2_X1  g056(.A(G1gat), .B(G29gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G57gat), .B(G85gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G225gat), .A2(G233gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n208_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT87), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NOR3_X1   g068(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT86), .ZN(new_n272_));
  OR2_X1    g071(.A1(G141gat), .A2(G148gat), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT3), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT85), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT3), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n273_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n278_));
  OAI22_X1  g077(.A1(new_n276_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT2), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n272_), .B1(new_n278_), .B2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G141gat), .A2(G148gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n276_), .A2(KEYINPUT3), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n274_), .A2(KEYINPUT85), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n286_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n289_), .A2(KEYINPUT86), .A3(new_n292_), .A4(new_n279_), .ZN(new_n293_));
  AOI211_X1 g092(.A(new_n267_), .B(new_n271_), .C1(new_n285_), .C2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n266_), .A2(KEYINPUT1), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(G155gat), .A3(G162gat), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n295_), .B(new_n297_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n280_), .A3(new_n273_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n265_), .B1(new_n294_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n285_), .A2(new_n293_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n271_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n266_), .A3(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(KEYINPUT87), .A3(new_n299_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n264_), .B1(new_n301_), .B2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n271_), .B1(new_n285_), .B2(new_n293_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n300_), .B1(new_n307_), .B2(new_n266_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n208_), .B(KEYINPUT92), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT4), .B1(new_n306_), .B2(new_n311_), .ZN(new_n312_));
  AOI211_X1 g111(.A(new_n265_), .B(new_n300_), .C1(new_n307_), .C2(new_n266_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT87), .B1(new_n304_), .B2(new_n299_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n208_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT4), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n263_), .B1(new_n312_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n263_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n306_), .A2(new_n319_), .A3(new_n311_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n262_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n316_), .B1(new_n315_), .B2(new_n310_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n306_), .A2(KEYINPUT4), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n319_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n320_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(new_n261_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT27), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT20), .ZN(new_n328_));
  INV_X1    g127(.A(G197gat), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(G204gat), .ZN(new_n330_));
  INV_X1    g129(.A(G204gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(G197gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT21), .B1(new_n330_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(G197gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(G204gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT21), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G211gat), .B(G218gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n333_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G211gat), .B(G218gat), .Z(new_n340_));
  OAI211_X1 g139(.A(new_n340_), .B(KEYINPUT21), .C1(new_n330_), .C2(new_n332_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n328_), .B1(new_n251_), .B2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n234_), .A2(new_n236_), .A3(new_n241_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n233_), .A2(new_n243_), .A3(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n342_), .A2(new_n250_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT91), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT91), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n342_), .A2(new_n349_), .A3(new_n250_), .A4(new_n346_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n344_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT19), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n246_), .A2(new_n342_), .A3(new_n250_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT20), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT90), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n346_), .A2(new_n250_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n343_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n356_), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n359_), .A2(new_n353_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364_));
  INV_X1    g163(.A(G92gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT18), .B(G64gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  AND3_X1   g167(.A1(new_n355_), .A2(new_n363_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n355_), .B2(new_n363_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n327_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n355_), .A2(new_n363_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n368_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n359_), .A2(new_n354_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n344_), .A2(new_n347_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n353_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n368_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n379_), .A3(KEYINPUT27), .ZN(new_n380_));
  AND4_X1   g179(.A1(new_n321_), .A2(new_n326_), .A3(new_n371_), .A4(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT94), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT88), .B1(new_n308_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT88), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n385_), .B(KEYINPUT29), .C1(new_n294_), .C2(new_n300_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n343_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT29), .B1(new_n313_), .B2(new_n314_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(new_n343_), .A3(new_n388_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G78gat), .B(G106gat), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n390_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G22gat), .B(G50gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT28), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n313_), .A2(new_n314_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(new_n383_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n301_), .A2(new_n383_), .A3(new_n305_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(KEYINPUT28), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n400_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n402_), .A2(new_n401_), .A3(new_n383_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(KEYINPUT28), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n399_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n390_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n398_), .A2(new_n410_), .B1(KEYINPUT89), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n406_), .A2(new_n409_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT89), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(new_n396_), .A4(new_n397_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n381_), .A2(new_n382_), .A3(new_n412_), .A4(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n394_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n409_), .B(new_n406_), .C1(new_n411_), .C2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n411_), .A2(KEYINPUT89), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n415_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n321_), .A2(new_n326_), .A3(new_n371_), .A4(new_n380_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT94), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n416_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n420_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425_));
  NOR4_X1   g224(.A1(new_n318_), .A2(new_n425_), .A3(new_n320_), .A4(new_n262_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n369_), .A2(new_n370_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n326_), .A2(new_n425_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n319_), .B1(new_n312_), .B2(new_n317_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n315_), .A2(new_n319_), .A3(new_n310_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n262_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .A4(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n321_), .A2(new_n326_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n373_), .A2(KEYINPUT32), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n436_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n372_), .A2(new_n436_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n424_), .B1(new_n434_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n256_), .B1(new_n423_), .B2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n435_), .A2(new_n256_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n371_), .A2(new_n380_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n420_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT12), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G99gat), .A2(G106gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT6), .ZN(new_n450_));
  INV_X1    g249(.A(G99gat), .ZN(new_n451_));
  INV_X1    g250(.A(G106gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n452_), .A3(KEYINPUT64), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT7), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n451_), .A2(new_n452_), .A3(KEYINPUT64), .A4(KEYINPUT7), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n450_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G85gat), .B(G92gat), .Z(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT8), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT10), .B(G99gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(G106gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n449_), .B(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G85gat), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n466_), .A2(new_n365_), .A3(KEYINPUT9), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n463_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n459_), .A2(KEYINPUT9), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n460_), .A2(new_n461_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT65), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n471_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n453_), .A2(new_n454_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(KEYINPUT65), .A3(new_n456_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n450_), .A3(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(KEYINPUT8), .A3(new_n459_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n470_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT66), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT66), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n470_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G57gat), .B(G64gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT11), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G71gat), .B(G78gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n482_), .B(KEYINPUT11), .Z(new_n486_));
  OAI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(new_n484_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n448_), .B1(new_n481_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G230gat), .A2(G233gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n481_), .A2(new_n488_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n477_), .A2(KEYINPUT12), .A3(new_n487_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .A4(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n481_), .A2(new_n488_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n487_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n495_));
  OAI211_X1 g294(.A(G230gat), .B(G233gat), .C1(new_n494_), .C2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT5), .B(G176gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(G204gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G120gat), .B(G148gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n493_), .A2(new_n496_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT67), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT67), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n493_), .A2(new_n496_), .A3(new_n504_), .A4(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT13), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n493_), .A2(new_n496_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n500_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n506_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n507_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G43gat), .B(G50gat), .ZN(new_n514_));
  INV_X1    g313(.A(G36gat), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n515_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT71), .B(G29gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT15), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT15), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n524_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527_));
  INV_X1    g326(.A(G1gat), .ZN(new_n528_));
  INV_X1    g327(.A(G8gat), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT14), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G1gat), .B(G8gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n526_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n533_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n522_), .A2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT76), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n522_), .B(new_n535_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(G229gat), .A3(G233gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT77), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G169gat), .B(G197gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  AND3_X1   g346(.A1(new_n543_), .A2(KEYINPUT78), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n547_), .B1(new_n543_), .B2(KEYINPUT78), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n513_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n447_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n480_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n479_), .B1(new_n470_), .B2(new_n476_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n522_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n526_), .A2(new_n477_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT69), .ZN(new_n559_));
  XOR2_X1   g358(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n561_), .A2(KEYINPUT35), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n557_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(KEYINPUT35), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT70), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n566_), .B1(new_n557_), .B2(KEYINPUT72), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n523_), .A2(new_n525_), .B1(new_n470_), .B2(new_n476_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT72), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n565_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n571_), .A2(new_n556_), .A3(new_n557_), .A4(new_n562_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT74), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT36), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n568_), .A2(KEYINPUT74), .A3(new_n572_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n575_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n578_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(KEYINPUT36), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n568_), .A2(new_n583_), .A3(new_n572_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n581_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n579_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n568_), .B2(new_n572_), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT37), .B1(new_n584_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT73), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT73), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n592_), .B(KEYINPUT37), .C1(new_n584_), .C2(new_n589_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n587_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n533_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(new_n487_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(G211gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT16), .B(G183gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT17), .Z(new_n602_));
  NOR2_X1   g401(.A1(new_n597_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(KEYINPUT17), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n604_), .B2(new_n597_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT75), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n606_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n594_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n553_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(new_n528_), .A3(new_n435_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT38), .ZN(new_n614_));
  INV_X1    g413(.A(new_n446_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n312_), .A2(new_n317_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n320_), .B1(new_n616_), .B2(new_n319_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT33), .B1(new_n617_), .B2(new_n261_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n369_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n619_), .B(new_n374_), .C1(new_n432_), .C2(new_n430_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n618_), .A2(new_n426_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n439_), .ZN(new_n622_));
  AOI211_X1 g421(.A(new_n437_), .B(new_n622_), .C1(new_n321_), .C2(new_n326_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n420_), .B1(new_n621_), .B2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(new_n422_), .A3(new_n416_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n615_), .B1(new_n625_), .B2(new_n256_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n581_), .A2(new_n585_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT95), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT96), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n631_), .A2(new_n610_), .A3(new_n552_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n632_), .A2(new_n435_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n614_), .B1(new_n633_), .B2(new_n528_), .ZN(G1324gat));
  NAND3_X1  g433(.A1(new_n612_), .A2(new_n529_), .A3(new_n444_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n631_), .A2(new_n610_), .A3(new_n552_), .A4(new_n444_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n636_), .A2(new_n637_), .A3(G8gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n636_), .B2(G8gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(KEYINPUT40), .B(new_n635_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n256_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n612_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n632_), .A2(new_n646_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n648_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT41), .B1(new_n648_), .B2(G15gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n647_), .B1(new_n649_), .B2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n612_), .A2(new_n652_), .A3(new_n424_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n631_), .A2(new_n610_), .A3(new_n552_), .A4(new_n424_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT42), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n654_), .A2(new_n655_), .A3(G22gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n654_), .B2(G22gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT97), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT97), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n660_), .B(new_n653_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(G1327gat));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n594_), .B(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT43), .B1(new_n626_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n587_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n416_), .A2(new_n422_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n646_), .B1(new_n668_), .B2(new_n624_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n666_), .B(new_n667_), .C1(new_n669_), .C2(new_n615_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n665_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n552_), .A2(new_n609_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n671_), .A2(KEYINPUT44), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n435_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n672_), .B1(new_n665_), .B2(new_n670_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(KEYINPUT44), .ZN(new_n677_));
  OAI21_X1  g476(.A(G29gat), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT99), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n610_), .A2(new_n627_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT100), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n553_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n435_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n683_), .A2(G29gat), .A3(new_n684_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n679_), .A2(new_n685_), .ZN(G1328gat));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(KEYINPUT46), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n444_), .B1(new_n676_), .B2(KEYINPUT44), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  AOI211_X1 g489(.A(new_n690_), .B(new_n672_), .C1(new_n665_), .C2(new_n670_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G36gat), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  OAI211_X1 g493(.A(KEYINPUT101), .B(G36gat), .C1(new_n689_), .C2(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n682_), .A2(new_n515_), .A3(new_n444_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n688_), .B1(new_n696_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n688_), .ZN(new_n702_));
  AOI211_X1 g501(.A(new_n702_), .B(new_n699_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1329gat));
  INV_X1    g503(.A(G43gat), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n691_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n676_), .A2(KEYINPUT44), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n646_), .A4(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n674_), .A2(G43gat), .A3(new_n646_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT103), .B1(new_n710_), .B2(new_n677_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n705_), .B1(new_n683_), .B2(new_n256_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT47), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n712_), .A2(new_n716_), .A3(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1330gat));
  AOI21_X1  g517(.A(G50gat), .B1(new_n682_), .B2(new_n424_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n677_), .A2(new_n420_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n674_), .A2(G50gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n719_), .B1(new_n720_), .B2(new_n721_), .ZN(G1331gat));
  INV_X1    g521(.A(new_n512_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n510_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(new_n550_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n726_), .A2(new_n626_), .A3(new_n611_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT104), .ZN(new_n728_));
  AOI21_X1  g527(.A(G57gat), .B1(new_n728_), .B2(new_n435_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n631_), .A2(new_n610_), .A3(new_n725_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n731_));
  OAI21_X1  g530(.A(G57gat), .B1(new_n684_), .B2(new_n731_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n731_), .A2(G57gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n729_), .B1(new_n733_), .B2(new_n734_), .ZN(G1332gat));
  NOR2_X1   g534(.A1(new_n445_), .A2(G64gat), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT106), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n728_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n730_), .A2(new_n444_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G64gat), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(KEYINPUT48), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(KEYINPUT48), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(G1333gat));
  NOR2_X1   g542(.A1(new_n256_), .A2(G71gat), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT107), .Z(new_n745_));
  NAND2_X1  g544(.A1(new_n728_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n730_), .A2(new_n646_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G71gat), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(G1334gat));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n728_), .A2(new_n752_), .A3(new_n424_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n730_), .A2(new_n424_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G78gat), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(KEYINPUT50), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(KEYINPUT50), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(G1335gat));
  NOR3_X1   g557(.A1(new_n726_), .A2(new_n626_), .A3(new_n681_), .ZN(new_n759_));
  AOI21_X1  g558(.A(G85gat), .B1(new_n759_), .B2(new_n435_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n725_), .A2(new_n609_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT108), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(new_n671_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n763_), .A2(new_n435_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n760_), .B1(new_n764_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g564(.A(G92gat), .B1(new_n759_), .B2(new_n444_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n763_), .A2(new_n444_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(G92gat), .ZN(G1337gat));
  AOI21_X1  g567(.A(new_n451_), .B1(new_n763_), .B2(new_n646_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n256_), .A2(new_n462_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n759_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(G1338gat));
  NAND3_X1  g572(.A1(new_n759_), .A2(new_n452_), .A3(new_n424_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n763_), .A2(new_n424_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(G106gat), .ZN(new_n777_));
  AOI211_X1 g576(.A(KEYINPUT52), .B(new_n452_), .C1(new_n763_), .C2(new_n424_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT53), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(new_n774_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1339gat));
  INV_X1    g582(.A(G113gat), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n503_), .A2(new_n505_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n490_), .A2(KEYINPUT112), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT55), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n493_), .A2(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n489_), .A2(KEYINPUT55), .A3(new_n491_), .A4(new_n492_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n790_), .A2(new_n787_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n500_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT56), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n501_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n792_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n786_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n506_), .A2(new_n509_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n540_), .A2(new_n542_), .A3(new_n547_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n547_), .B1(new_n541_), .B2(new_n539_), .ZN(new_n801_));
  XOR2_X1   g600(.A(new_n801_), .B(KEYINPUT113), .Z(new_n802_));
  INV_X1    g601(.A(new_n537_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n803_), .A2(new_n539_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n800_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n798_), .A2(new_n550_), .B1(new_n799_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n627_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n785_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n799_), .A2(new_n805_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n793_), .A2(new_n794_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT56), .B1(new_n796_), .B2(new_n792_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n506_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n809_), .B1(new_n812_), .B2(new_n551_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(KEYINPUT57), .A3(new_n627_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n808_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n506_), .B(new_n805_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n816_), .A2(KEYINPUT114), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n816_), .B2(KEYINPUT114), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n594_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n609_), .B1(new_n815_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n611_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n550_), .B1(new_n723_), .B2(new_n510_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT110), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n551_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT54), .B1(new_n827_), .B2(new_n611_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT110), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n822_), .A2(new_n823_), .A3(new_n831_), .A4(new_n824_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT111), .B(KEYINPUT54), .C1(new_n827_), .C2(new_n611_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n826_), .A2(new_n830_), .A3(new_n832_), .A4(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n821_), .A2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n684_), .A2(new_n444_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n835_), .A2(new_n646_), .A3(new_n420_), .A4(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n784_), .B1(new_n837_), .B2(new_n551_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n839_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n837_), .A2(KEYINPUT59), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n424_), .B1(new_n821_), .B2(new_n834_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n646_), .A4(new_n836_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n842_), .A2(G113gat), .A3(new_n550_), .A4(new_n845_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n840_), .A2(new_n841_), .A3(new_n846_), .ZN(G1340gat));
  NAND3_X1  g646(.A1(new_n842_), .A2(new_n513_), .A3(new_n845_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G120gat), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT60), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n837_), .B1(new_n850_), .B2(G120gat), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n724_), .A2(KEYINPUT60), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(G120gat), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n853_), .ZN(G1341gat));
  NAND2_X1  g653(.A1(new_n610_), .A2(G127gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT116), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n842_), .A2(new_n845_), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(G127gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n837_), .B2(new_n609_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT117), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n857_), .A2(new_n862_), .A3(new_n859_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(G1342gat));
  INV_X1    g663(.A(G134gat), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n594_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n842_), .A2(new_n845_), .A3(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n865_), .B1(new_n837_), .B2(new_n628_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n867_), .A2(KEYINPUT118), .A3(new_n868_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1343gat));
  NAND3_X1  g672(.A1(new_n836_), .A2(new_n256_), .A3(new_n424_), .ZN(new_n874_));
  XOR2_X1   g673(.A(new_n874_), .B(KEYINPUT119), .Z(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n821_), .B2(new_n834_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n550_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT120), .B(G141gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1344gat));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n513_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g680(.A1(new_n876_), .A2(new_n610_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G155gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n883_), .B(new_n885_), .ZN(G1346gat));
  AOI21_X1  g685(.A(G162gat), .B1(new_n876_), .B2(new_n629_), .ZN(new_n887_));
  INV_X1    g686(.A(G162gat), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n664_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n887_), .B1(new_n876_), .B2(new_n889_), .ZN(G1347gat));
  NAND4_X1  g689(.A1(new_n835_), .A2(new_n420_), .A3(new_n444_), .A4(new_n443_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT122), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n843_), .A2(new_n893_), .A3(new_n444_), .A4(new_n443_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n892_), .A2(new_n550_), .A3(new_n247_), .A4(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896_));
  INV_X1    g695(.A(new_n891_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n550_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n896_), .B1(new_n898_), .B2(G169gat), .ZN(new_n899_));
  AOI211_X1 g698(.A(KEYINPUT62), .B(new_n219_), .C1(new_n897_), .C2(new_n550_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n895_), .B1(new_n899_), .B2(new_n900_), .ZN(G1348gat));
  OAI21_X1  g700(.A(G176gat), .B1(new_n891_), .B2(new_n724_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n892_), .A2(new_n220_), .A3(new_n894_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n724_), .ZN(G1349gat));
  AOI21_X1  g703(.A(new_n609_), .B1(new_n236_), .B2(new_n241_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n892_), .A2(new_n894_), .A3(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n240_), .B1(new_n891_), .B2(new_n609_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT123), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n906_), .A2(new_n910_), .A3(new_n907_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1350gat));
  NAND3_X1  g711(.A1(new_n892_), .A2(new_n667_), .A3(new_n894_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G190gat), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n892_), .A2(new_n629_), .A3(new_n234_), .A4(new_n894_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1351gat));
  NOR3_X1   g715(.A1(new_n420_), .A2(new_n646_), .A3(new_n435_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(KEYINPUT124), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n821_), .B2(new_n834_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n445_), .B1(new_n917_), .B2(KEYINPUT124), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n551_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(new_n329_), .ZN(G1352gat));
  INV_X1    g722(.A(new_n921_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n513_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n331_), .A2(KEYINPUT125), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n331_), .A2(KEYINPUT125), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n925_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n928_), .B1(new_n925_), .B2(new_n926_), .ZN(G1353gat));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n930_));
  INV_X1    g729(.A(G211gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n610_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT126), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n924_), .A2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n930_), .A2(new_n931_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1354gat));
  AND3_X1   g735(.A1(new_n924_), .A2(G218gat), .A3(new_n667_), .ZN(new_n937_));
  AOI21_X1  g736(.A(G218gat), .B1(new_n924_), .B2(new_n629_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1355gat));
endmodule


