//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n965_, new_n966_,
    new_n968_, new_n969_, new_n970_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_, new_n982_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT94), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT4), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT85), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(KEYINPUT84), .B2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT84), .B(KEYINPUT3), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(new_n209_), .B2(new_n206_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n205_), .B1(new_n210_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n206_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n207_), .A2(KEYINPUT84), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n207_), .A2(KEYINPUT84), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n211_), .B(KEYINPUT2), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT85), .A4(new_n208_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n214_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G155gat), .ZN(new_n222_));
  INV_X1    g021(.A(G162gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(KEYINPUT83), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT83), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n225_), .B1(G155gat), .B2(G162gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT86), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n224_), .A2(new_n226_), .A3(KEYINPUT86), .A4(new_n227_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n221_), .A2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n215_), .A2(KEYINPUT82), .ZN(new_n235_));
  AND3_X1   g034(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n224_), .B(new_n226_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n211_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n239_), .B1(new_n215_), .B2(KEYINPUT82), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n235_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G127gat), .B(G134gat), .Z(new_n242_));
  XOR2_X1   g041(.A(G113gat), .B(G120gat), .Z(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G113gat), .B(G120gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n234_), .A2(new_n241_), .A3(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT79), .B1(new_n245_), .B2(new_n246_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(new_n244_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n232_), .B1(new_n214_), .B2(new_n220_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n241_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n251_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n204_), .B1(new_n249_), .B2(new_n254_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n254_), .A2(new_n204_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n203_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n203_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n249_), .A2(new_n258_), .A3(new_n254_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G57gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(G85gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(G1gat), .B(G29gat), .Z(new_n263_));
  XOR2_X1   g062(.A(new_n262_), .B(new_n263_), .Z(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n264_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n257_), .A2(new_n259_), .A3(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n265_), .A2(KEYINPUT98), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT98), .B1(new_n265_), .B2(new_n267_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G15gat), .B(G43gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G227gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G71gat), .B(G99gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT78), .ZN(new_n276_));
  OR2_X1    g075(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(G176gat), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n276_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n278_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(KEYINPUT78), .A3(new_n280_), .ZN(new_n287_));
  INV_X1    g086(.A(G183gat), .ZN(new_n288_));
  INV_X1    g087(.A(G190gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT23), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(G183gat), .A3(G190gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n289_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n282_), .A2(new_n287_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT30), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT25), .B(G183gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT76), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT26), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n299_), .B1(new_n300_), .B2(G190gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT26), .B(G190gat), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n298_), .B(new_n301_), .C1(new_n302_), .C2(new_n299_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n292_), .A2(KEYINPUT77), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n305_), .A2(new_n291_), .A3(G183gat), .A4(G190gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n290_), .A3(new_n306_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n280_), .A2(KEYINPUT24), .ZN(new_n309_));
  INV_X1    g108(.A(G169gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n283_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n308_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n303_), .A2(new_n307_), .A3(new_n312_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n296_), .A2(new_n297_), .A3(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n297_), .B1(new_n296_), .B2(new_n313_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n275_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n296_), .A2(new_n313_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT30), .ZN(new_n318_));
  INV_X1    g117(.A(new_n274_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n273_), .B(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n296_), .A2(new_n297_), .A3(new_n313_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT80), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n316_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n251_), .B(KEYINPUT31), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n323_), .B1(new_n316_), .B2(new_n322_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AOI211_X1 g127(.A(new_n323_), .B(new_n325_), .C1(new_n322_), .C2(new_n316_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT81), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n326_), .A2(new_n327_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n316_), .A2(new_n322_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT80), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT81), .B1(new_n332_), .B2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n331_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT91), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n339_), .B1(new_n234_), .B2(new_n241_), .ZN(new_n340_));
  INV_X1    g139(.A(G197gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n341_), .A2(G204gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT87), .ZN(new_n343_));
  INV_X1    g142(.A(G204gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n343_), .B1(new_n344_), .B2(G197gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n342_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT21), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  AND2_X1   g148(.A1(G211gat), .A2(G218gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(G211gat), .A2(G218gat), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT88), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(G211gat), .ZN(new_n353_));
  INV_X1    g152(.A(G218gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT88), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G211gat), .A2(G218gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n352_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n344_), .A2(G197gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT21), .B1(new_n342_), .B2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n349_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n347_), .A2(new_n348_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n352_), .A2(new_n358_), .A3(KEYINPUT89), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT89), .B1(new_n352_), .B2(new_n358_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT90), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  OAI211_X1 g168(.A(KEYINPUT90), .B(new_n364_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n363_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n340_), .A2(new_n371_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT89), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n359_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n352_), .A2(new_n358_), .A3(KEYINPUT89), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT90), .B1(new_n378_), .B2(new_n364_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n370_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n362_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT29), .B1(new_n252_), .B2(new_n253_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n372_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n338_), .B1(new_n374_), .B2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n373_), .B1(new_n340_), .B2(new_n371_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n372_), .A3(new_n382_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(KEYINPUT91), .A3(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(G22gat), .B(G50gat), .Z(new_n388_));
  INV_X1    g187(.A(KEYINPUT28), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n253_), .B1(new_n221_), .B2(new_n233_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n390_), .B2(new_n339_), .ZN(new_n391_));
  NOR4_X1   g190(.A1(new_n252_), .A2(new_n253_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n388_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n234_), .A2(new_n339_), .A3(new_n241_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT28), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n390_), .A2(new_n389_), .A3(new_n339_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n388_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n384_), .A2(new_n387_), .B1(new_n393_), .B2(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n385_), .A2(KEYINPUT91), .A3(new_n386_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n393_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G78gat), .B(G106gat), .Z(new_n403_));
  NOR3_X1   g202(.A1(new_n399_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT91), .B1(new_n385_), .B2(new_n386_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n401_), .B1(new_n400_), .B2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n387_), .A2(new_n393_), .A3(new_n398_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n405_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n337_), .B1(new_n404_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n403_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n328_), .A2(new_n329_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n407_), .A2(new_n405_), .A3(new_n408_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n270_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G8gat), .B(G36gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n418_), .B(new_n419_), .Z(new_n420_));
  INV_X1    g219(.A(new_n317_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n421_), .B(new_n362_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n293_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n302_), .A2(KEYINPUT92), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT92), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n300_), .A2(G190gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n289_), .A2(KEYINPUT26), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n424_), .A2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n423_), .B1(new_n429_), .B2(new_n298_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n279_), .A2(new_n281_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n307_), .A2(new_n294_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n430_), .A2(new_n312_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n422_), .B(KEYINPUT20), .C1(new_n371_), .C2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G226gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT19), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n381_), .A2(new_n317_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n436_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n433_), .B(new_n362_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n438_), .A2(KEYINPUT20), .A3(new_n439_), .A4(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n420_), .B1(new_n437_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n437_), .A2(new_n441_), .A3(new_n420_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT27), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT99), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT96), .B(KEYINPUT20), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n371_), .B2(new_n433_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n438_), .B1(new_n448_), .B2(KEYINPUT97), .ZN(new_n449_));
  INV_X1    g248(.A(new_n447_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n440_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT97), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n436_), .B1(new_n449_), .B2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n434_), .A2(new_n436_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n420_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n444_), .A2(KEYINPUT27), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n446_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n420_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n451_), .A2(new_n452_), .B1(new_n381_), .B2(new_n317_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n448_), .A2(KEYINPUT97), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n439_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n460_), .B1(new_n463_), .B2(new_n455_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT27), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n440_), .A2(KEYINPUT20), .A3(new_n439_), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n438_), .A2(new_n466_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n467_), .B2(new_n420_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(KEYINPUT99), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n445_), .B1(new_n459_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n330_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n332_), .A2(new_n335_), .A3(KEYINPUT81), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n444_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n474_), .A2(new_n442_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n258_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n249_), .A2(new_n203_), .A3(new_n254_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n477_), .A2(new_n264_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n476_), .A2(new_n478_), .A3(KEYINPUT95), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT95), .B1(new_n476_), .B2(new_n478_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT33), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n267_), .A2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n257_), .A2(KEYINPUT33), .A3(new_n259_), .A4(new_n266_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n475_), .A2(new_n481_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n420_), .A2(KEYINPUT32), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n265_), .A2(new_n267_), .B1(new_n467_), .B2(new_n486_), .ZN(new_n487_));
  OAI211_X1 g286(.A(KEYINPUT32), .B(new_n420_), .C1(new_n463_), .C2(new_n455_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n473_), .B1(new_n485_), .B2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n404_), .A2(new_n409_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n415_), .A2(new_n470_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT74), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT16), .B(G183gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(G211gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G127gat), .B(G155gat), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n496_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n493_), .B1(new_n499_), .B2(KEYINPUT17), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G231gat), .A2(G233gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G15gat), .B(G22gat), .ZN(new_n503_));
  INV_X1    g302(.A(G1gat), .ZN(new_n504_));
  INV_X1    g303(.A(G8gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G1gat), .B(G8gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n501_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n510_), .B1(new_n512_), .B2(new_n493_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n502_), .A2(new_n509_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n509_), .B1(new_n502_), .B2(new_n513_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G57gat), .B(G64gat), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n517_), .A2(KEYINPUT11), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(KEYINPUT11), .ZN(new_n519_));
  XOR2_X1   g318(.A(G71gat), .B(G78gat), .Z(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n519_), .A2(new_n520_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n515_), .A2(new_n516_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n523_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n502_), .A2(new_n513_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n509_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n525_), .B1(new_n528_), .B2(new_n514_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n524_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n497_), .A2(new_n511_), .A3(new_n498_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT69), .B(KEYINPUT35), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(G50gat), .ZN(new_n536_));
  INV_X1    g335(.A(G29gat), .ZN(new_n537_));
  INV_X1    g336(.A(G36gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(G43gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G29gat), .A2(G36gat), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n536_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(G50gat), .A3(new_n542_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT6), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT66), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT66), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT6), .ZN(new_n553_));
  AND2_X1   g352(.A1(G99gat), .A2(G106gat), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n551_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT10), .B(G99gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT64), .B(G106gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT65), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(G85gat), .ZN(new_n563_));
  INV_X1    g362(.A(G92gat), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n563_), .A2(new_n564_), .A3(KEYINPUT9), .ZN(new_n565_));
  XOR2_X1   g364(.A(G85gat), .B(G92gat), .Z(new_n566_));
  AOI21_X1  g365(.A(new_n565_), .B1(new_n566_), .B2(KEYINPUT9), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n558_), .A2(KEYINPUT65), .A3(new_n559_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n557_), .A2(new_n562_), .A3(new_n567_), .A4(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n570_));
  OR3_X1    g369(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n570_), .B(new_n571_), .C1(new_n555_), .C2(new_n556_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT8), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n572_), .A2(new_n573_), .A3(new_n566_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n572_), .B2(new_n566_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n549_), .B(new_n569_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n535_), .B1(new_n576_), .B2(KEYINPUT70), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT68), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT34), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n545_), .A2(new_n547_), .A3(KEYINPUT15), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT15), .B1(new_n545_), .B2(new_n547_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n569_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n580_), .A2(new_n534_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n576_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n581_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n586_), .A2(new_n576_), .A3(new_n587_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n580_), .A3(new_n577_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(G134gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(new_n223_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT36), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n595_), .A2(new_n596_), .ZN(new_n598_));
  OR3_X1    g397(.A1(new_n597_), .A2(new_n598_), .A3(KEYINPUT71), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT71), .B1(new_n597_), .B2(new_n598_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT73), .B1(new_n592_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT73), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n589_), .A2(new_n591_), .A3(new_n597_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n602_), .A2(new_n603_), .A3(new_n606_), .A4(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n607_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT37), .B1(new_n609_), .B2(new_n604_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT72), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT72), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n612_), .B(KEYINPUT37), .C1(new_n609_), .C2(new_n604_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n608_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n492_), .A2(new_n533_), .A3(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT67), .B(KEYINPUT13), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(new_n344_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT5), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(new_n283_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n585_), .A2(new_n525_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n569_), .B(new_n523_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(KEYINPUT12), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT12), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n585_), .A2(new_n626_), .A3(new_n525_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n622_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n629_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n622_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n635_), .A2(new_n631_), .A3(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n618_), .B1(new_n633_), .B2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n630_), .A2(new_n632_), .A3(new_n622_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n636_), .B1(new_n635_), .B2(new_n631_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT13), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n639_), .B(new_n640_), .C1(KEYINPUT67), .C2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n638_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(G229gat), .A2(G233gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n549_), .A2(new_n527_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n548_), .A2(new_n509_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G113gat), .B(G141gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(new_n310_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(new_n341_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n584_), .A2(new_n509_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n654_), .B1(new_n548_), .B2(new_n509_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n649_), .B(new_n653_), .C1(new_n655_), .C2(new_n646_), .ZN(new_n656_));
  AOI211_X1 g455(.A(new_n646_), .B(new_n648_), .C1(new_n584_), .C2(new_n509_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n649_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n652_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n656_), .A2(KEYINPUT75), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT75), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n661_), .B(new_n652_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n644_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n616_), .A2(new_n664_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n268_), .A2(new_n269_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n665_), .A2(G1gat), .A3(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n602_), .A2(new_n607_), .A3(new_n606_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n485_), .A2(new_n489_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n337_), .A3(new_n491_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n473_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n666_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n459_), .A2(new_n469_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n445_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n673_), .B1(new_n676_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n663_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT101), .B1(new_n643_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n683_));
  AOI211_X1 g482(.A(new_n683_), .B(new_n663_), .C1(new_n638_), .C2(new_n642_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  AND4_X1   g484(.A1(new_n671_), .A2(new_n680_), .A3(new_n685_), .A4(new_n532_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n504_), .B1(new_n686_), .B2(new_n270_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT102), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n669_), .A2(new_n688_), .ZN(G1324gat));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n679_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G8gat), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT39), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(KEYINPUT103), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n665_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(new_n505_), .A3(new_n679_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(KEYINPUT103), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n692_), .A2(KEYINPUT103), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n690_), .A2(G8gat), .A3(new_n696_), .A4(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n693_), .A2(new_n695_), .A3(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g499(.A(G15gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n686_), .B2(new_n473_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT41), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n694_), .A2(new_n701_), .A3(new_n473_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1326gat));
  INV_X1    g504(.A(G22gat), .ZN(new_n706_));
  INV_X1    g505(.A(new_n491_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n686_), .B2(new_n707_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT42), .Z(new_n709_));
  NAND3_X1  g508(.A1(new_n694_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1327gat));
  NAND3_X1  g510(.A1(new_n680_), .A2(new_n670_), .A3(new_n533_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n712_), .A2(new_n663_), .A3(new_n644_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G29gat), .B1(new_n713_), .B2(new_n270_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT43), .B1(new_n492_), .B2(new_n614_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n680_), .A2(new_n716_), .A3(new_n615_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n533_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT104), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n720_), .B(new_n533_), .C1(new_n682_), .C2(new_n684_), .ZN(new_n721_));
  AOI22_X1  g520(.A1(new_n715_), .A2(new_n717_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n722_), .A2(KEYINPUT44), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n723_), .A2(new_n537_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n666_), .B1(new_n722_), .B2(KEYINPUT44), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n714_), .B1(new_n724_), .B2(new_n725_), .ZN(G1328gat));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n470_), .B1(new_n722_), .B2(KEYINPUT44), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n719_), .A2(new_n721_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n716_), .B1(new_n680_), .B2(new_n615_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n410_), .A2(new_n414_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n731_), .A2(new_n666_), .A3(new_n470_), .ZN(new_n732_));
  AOI211_X1 g531(.A(KEYINPUT43), .B(new_n614_), .C1(new_n732_), .C2(new_n673_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n730_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n538_), .B1(new_n728_), .B2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n713_), .A2(KEYINPUT45), .A3(new_n538_), .A4(new_n679_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n492_), .A2(new_n671_), .A3(new_n532_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(new_n538_), .A3(new_n664_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n741_), .B2(new_n470_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n727_), .B1(new_n737_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n743_), .ZN(new_n745_));
  OAI211_X1 g544(.A(KEYINPUT44), .B(new_n729_), .C1(new_n730_), .C2(new_n733_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n679_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G36gat), .B1(new_n747_), .B2(new_n723_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(KEYINPUT105), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT46), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n744_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT106), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n745_), .A2(KEYINPUT46), .A3(new_n748_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n744_), .A2(new_n749_), .A3(new_n754_), .A4(new_n750_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(new_n753_), .A3(new_n755_), .ZN(G1329gat));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n412_), .B1(new_n722_), .B2(KEYINPUT44), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n746_), .A2(G43gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT107), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n412_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n540_), .B1(new_n722_), .B2(KEYINPUT44), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n763_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(G43gat), .B1(new_n713_), .B2(new_n473_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n758_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  AOI211_X1 g569(.A(KEYINPUT108), .B(new_n768_), .C1(new_n761_), .C2(new_n766_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n757_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n759_), .A2(new_n760_), .A3(KEYINPUT107), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n765_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n769_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT108), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n767_), .A2(new_n758_), .A3(new_n769_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(KEYINPUT47), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n772_), .A2(new_n778_), .ZN(G1330gat));
  NAND2_X1  g578(.A1(new_n707_), .A2(new_n536_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT109), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n713_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n746_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n783_), .A2(new_n723_), .A3(new_n491_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n782_), .B1(new_n784_), .B2(new_n536_), .ZN(G1331gat));
  NOR2_X1   g584(.A1(new_n643_), .A2(new_n681_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n616_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(G57gat), .B1(new_n788_), .B2(new_n270_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n786_), .ZN(new_n790_));
  NOR4_X1   g589(.A1(new_n492_), .A2(new_n670_), .A3(new_n533_), .A4(new_n790_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n270_), .A2(G57gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n789_), .B1(new_n791_), .B2(new_n792_), .ZN(G1332gat));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n679_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(G64gat), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT110), .Z(new_n796_));
  AND2_X1   g595(.A1(new_n796_), .A2(KEYINPUT48), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(KEYINPUT48), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n470_), .A2(G64gat), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n799_), .B(KEYINPUT111), .Z(new_n800_));
  OAI22_X1  g599(.A1(new_n797_), .A2(new_n798_), .B1(new_n787_), .B2(new_n800_), .ZN(G1333gat));
  INV_X1    g600(.A(G71gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n791_), .B2(new_n473_), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n803_), .B(KEYINPUT49), .Z(new_n804_));
  NAND3_X1  g603(.A1(new_n788_), .A2(new_n802_), .A3(new_n473_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1334gat));
  INV_X1    g605(.A(G78gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n791_), .B2(new_n707_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT112), .B(KEYINPUT113), .Z(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT50), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n808_), .B(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n788_), .A2(new_n807_), .A3(new_n707_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(G1335gat));
  AOI211_X1 g612(.A(new_n532_), .B(new_n790_), .C1(new_n715_), .C2(new_n717_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(G85gat), .A3(new_n270_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n712_), .A2(new_n790_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n563_), .B1(new_n817_), .B2(new_n666_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n815_), .A2(new_n818_), .ZN(G1336gat));
  NAND3_X1  g618(.A1(new_n814_), .A2(G92gat), .A3(new_n679_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n564_), .B1(new_n817_), .B2(new_n470_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1337gat));
  AND3_X1   g621(.A1(new_n816_), .A2(new_n558_), .A3(new_n412_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n814_), .A2(new_n473_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(G99gat), .ZN(new_n825_));
  XOR2_X1   g624(.A(new_n825_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g625(.A1(new_n816_), .A2(new_n559_), .A3(new_n707_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n715_), .A2(new_n717_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(new_n707_), .A3(new_n533_), .A4(new_n786_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n829_), .A2(new_n830_), .A3(G106gat), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n829_), .B2(G106gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n827_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT114), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n835_), .B(new_n827_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n834_), .A2(KEYINPUT53), .A3(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT53), .B1(new_n834_), .B2(new_n836_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(G1339gat));
  NOR2_X1   g638(.A1(new_n679_), .A2(new_n666_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n628_), .A2(new_n629_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n630_), .A2(KEYINPUT55), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n635_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n843_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT56), .B1(new_n847_), .B2(new_n622_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n635_), .A2(new_n845_), .ZN(new_n849_));
  AOI211_X1 g648(.A(KEYINPUT55), .B(new_n634_), .C1(new_n625_), .C2(new_n627_), .ZN(new_n850_));
  OAI22_X1  g649(.A1(new_n849_), .A2(new_n850_), .B1(new_n629_), .B2(new_n628_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n636_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n848_), .A2(new_n681_), .A3(new_n639_), .A4(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n645_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n855_), .A2(new_n652_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n856_), .A2(KEYINPUT116), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(KEYINPUT116), .A3(new_n652_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n857_), .B(new_n858_), .C1(new_n645_), .C2(new_n655_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n859_), .A2(new_n656_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n633_), .B2(new_n637_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n854_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n842_), .B1(new_n862_), .B2(new_n671_), .ZN(new_n863_));
  AOI211_X1 g662(.A(new_n670_), .B(new_n841_), .C1(new_n854_), .C2(new_n861_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n847_), .A2(KEYINPUT56), .A3(new_n622_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n852_), .B1(new_n851_), .B2(new_n636_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n868_), .A2(KEYINPUT58), .A3(new_n639_), .A4(new_n860_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n848_), .A2(new_n860_), .A3(new_n639_), .A4(new_n853_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n869_), .A2(new_n615_), .A3(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n532_), .B1(new_n865_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n532_), .A2(new_n663_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT115), .B1(new_n644_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n643_), .A2(new_n877_), .A3(new_n532_), .A4(new_n663_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n878_), .A3(new_n614_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n876_), .A2(new_n878_), .A3(new_n614_), .A4(KEYINPUT54), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n674_), .B(new_n840_), .C1(new_n874_), .C2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(G113gat), .B1(new_n885_), .B2(new_n681_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n884_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n862_), .A2(new_n671_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n841_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n862_), .A2(new_n671_), .A3(new_n842_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(new_n891_), .A3(new_n873_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n533_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n883_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n895_), .A2(KEYINPUT59), .A3(new_n674_), .A4(new_n840_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n888_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n681_), .A2(G113gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT118), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n886_), .B1(new_n897_), .B2(new_n899_), .ZN(G1340gat));
  INV_X1    g699(.A(G120gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n901_), .B1(new_n643_), .B2(KEYINPUT60), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT119), .B1(new_n901_), .B2(KEYINPUT60), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n884_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n902_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n643_), .B1(new_n888_), .B2(new_n896_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n901_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(KEYINPUT120), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n907_), .B(new_n911_), .C1(new_n908_), .C2(new_n901_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(G1341gat));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n914_));
  INV_X1    g713(.A(new_n840_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n915_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n916_));
  AOI21_X1  g715(.A(KEYINPUT59), .B1(new_n916_), .B2(new_n674_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n883_), .B1(new_n892_), .B2(new_n533_), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n918_), .A2(new_n887_), .A3(new_n414_), .A4(new_n915_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n532_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(G127gat), .ZN(new_n921_));
  INV_X1    g720(.A(G127gat), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n885_), .A2(new_n922_), .A3(new_n532_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n914_), .B1(new_n921_), .B2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n533_), .B1(new_n888_), .B2(new_n896_), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n914_), .B(new_n923_), .C1(new_n925_), .C2(new_n922_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n924_), .A2(new_n927_), .ZN(G1342gat));
  AOI21_X1  g727(.A(G134gat), .B1(new_n885_), .B2(new_n670_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n614_), .B1(new_n888_), .B2(new_n896_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n930_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g730(.A1(new_n916_), .A2(new_n675_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n663_), .ZN(new_n933_));
  XOR2_X1   g732(.A(new_n933_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g733(.A1(new_n932_), .A2(new_n643_), .ZN(new_n935_));
  XOR2_X1   g734(.A(KEYINPUT122), .B(G148gat), .Z(new_n936_));
  XNOR2_X1  g735(.A(new_n935_), .B(new_n936_), .ZN(G1345gat));
  NAND3_X1  g736(.A1(new_n916_), .A2(new_n675_), .A3(new_n532_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(KEYINPUT123), .B(KEYINPUT124), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n938_), .A2(new_n939_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(KEYINPUT61), .B(G155gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1346gat));
  NOR3_X1   g743(.A1(new_n932_), .A2(new_n223_), .A3(new_n614_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n916_), .A2(new_n670_), .A3(new_n675_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n223_), .B2(new_n946_), .ZN(G1347gat));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n918_), .A2(new_n707_), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n470_), .A2(new_n270_), .A3(new_n337_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n951_), .A2(new_n663_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n948_), .B1(new_n952_), .B2(new_n310_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n285_), .B2(new_n284_), .ZN(new_n954_));
  OAI211_X1 g753(.A(KEYINPUT62), .B(G169gat), .C1(new_n951_), .C2(new_n663_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n953_), .A2(new_n954_), .A3(new_n955_), .ZN(G1348gat));
  NOR2_X1   g755(.A1(new_n951_), .A2(new_n643_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(new_n283_), .ZN(G1349gat));
  OR3_X1    g757(.A1(new_n951_), .A2(new_n298_), .A3(new_n533_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n959_), .A2(new_n960_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n288_), .B1(new_n951_), .B2(new_n533_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(KEYINPUT125), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n961_), .B1(new_n959_), .B2(new_n963_), .ZN(G1350gat));
  OAI21_X1  g763(.A(G190gat), .B1(new_n951_), .B2(new_n614_), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n949_), .A2(new_n429_), .A3(new_n950_), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n965_), .B1(new_n671_), .B2(new_n966_), .ZN(G1351gat));
  NOR3_X1   g766(.A1(new_n470_), .A2(new_n270_), .A3(new_n410_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n895_), .A2(new_n968_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n969_), .A2(new_n663_), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n970_), .B(new_n341_), .ZN(G1352gat));
  NOR2_X1   g770(.A1(new_n969_), .A2(new_n643_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(new_n344_), .ZN(G1353gat));
  INV_X1    g772(.A(new_n969_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n974_), .A2(new_n532_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n976_));
  AND2_X1   g775(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n975_), .A2(new_n976_), .A3(new_n977_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n978_), .B1(new_n975_), .B2(new_n976_), .ZN(G1354gat));
  AOI21_X1  g778(.A(G218gat), .B1(new_n974_), .B2(new_n670_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n615_), .A2(G218gat), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n981_), .B(KEYINPUT126), .ZN(new_n982_));
  AOI21_X1  g781(.A(new_n980_), .B1(new_n974_), .B2(new_n982_), .ZN(G1355gat));
endmodule


