//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_;
  OAI21_X1  g000(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n202_));
  AOI21_X1  g001(.A(new_n202_), .B1(G169gat), .B2(G176gat), .ZN(new_n203_));
  NOR3_X1   g002(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT25), .B(G183gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT79), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT26), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n207_), .B1(new_n208_), .B2(G190gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT26), .B(G190gat), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n206_), .B(new_n209_), .C1(new_n210_), .C2(new_n207_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT81), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n214_));
  NOR2_X1   g013(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n212_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT80), .B(KEYINPUT23), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT81), .B1(new_n220_), .B2(new_n213_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n205_), .B(new_n211_), .C1(new_n219_), .C2(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(G183gat), .B(G190gat), .C1(new_n214_), .C2(new_n215_), .ZN(new_n223_));
  OR2_X1    g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n213_), .A2(new_n217_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(G169gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n222_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT82), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n222_), .A2(KEYINPUT82), .A3(new_n229_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G15gat), .B(G43gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT84), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n234_), .B(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT31), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n234_), .A2(new_n236_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n234_), .A2(new_n236_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT31), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G227gat), .A2(G233gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n243_), .B(G71gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G99gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G127gat), .B(G134gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G113gat), .B(G120gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n247_), .B(new_n250_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n238_), .A2(new_n242_), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n251_), .B1(new_n238_), .B2(new_n242_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT92), .ZN(new_n255_));
  INV_X1    g054(.A(G218gat), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n256_), .A2(G211gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(G211gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n255_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G211gat), .B(G218gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT92), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n261_), .A3(KEYINPUT21), .ZN(new_n262_));
  INV_X1    g061(.A(G204gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT89), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT89), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G204gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n266_), .A3(G197gat), .ZN(new_n267_));
  INV_X1    g066(.A(G197gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT90), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(new_n263_), .B2(G197gat), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n267_), .A2(new_n269_), .A3(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n262_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT21), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n267_), .A2(new_n274_), .A3(new_n269_), .A4(new_n271_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT91), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n271_), .A2(new_n269_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n278_), .A2(KEYINPUT91), .A3(new_n274_), .A4(new_n267_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n264_), .A2(new_n266_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n268_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n274_), .B1(G197gat), .B2(G204gat), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n282_), .A2(new_n283_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n273_), .B1(new_n280_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT3), .ZN(new_n287_));
  INV_X1    g086(.A(G141gat), .ZN(new_n288_));
  INV_X1    g087(.A(G148gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT2), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n290_), .A2(new_n293_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT86), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT85), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT85), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT86), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n299_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n302_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n296_), .B(new_n297_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n297_), .A2(KEYINPUT1), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT1), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(G155gat), .A3(G162gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n302_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n300_), .A2(KEYINPUT86), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n298_), .A2(KEYINPUT85), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n299_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n309_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n288_), .A2(new_n289_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n291_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n305_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT88), .B1(new_n318_), .B2(KEYINPUT29), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G228gat), .A2(G233gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n320_), .B(G78gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G106gat), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n286_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(new_n286_), .B2(new_n319_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT93), .ZN(new_n326_));
  XOR2_X1   g125(.A(G22gat), .B(G50gat), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT28), .B1(new_n318_), .B2(KEYINPUT29), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n303_), .A2(new_n304_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n291_), .B(new_n316_), .C1(new_n330_), .C2(new_n309_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .A4(new_n305_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT87), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n329_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n335_), .B1(new_n329_), .B2(new_n334_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n328_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n329_), .A2(new_n334_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT87), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n329_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n327_), .A3(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n325_), .A2(new_n326_), .A3(new_n338_), .A4(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n338_), .A2(new_n342_), .A3(new_n326_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n325_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n326_), .B1(new_n338_), .B2(new_n342_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n343_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT19), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n232_), .A2(new_n285_), .A3(new_n233_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT20), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT94), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n216_), .A2(new_n212_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n213_), .A2(KEYINPUT23), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n220_), .B2(new_n213_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n354_), .B1(new_n356_), .B2(new_n212_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n353_), .B1(new_n357_), .B2(new_n224_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n353_), .B(new_n224_), .C1(new_n219_), .C2(new_n221_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n228_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n223_), .A2(new_n225_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n210_), .A2(new_n206_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n205_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n285_), .B1(new_n361_), .B2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n350_), .B1(new_n352_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT97), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n361_), .A2(new_n285_), .A3(new_n364_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT82), .B1(new_n222_), .B2(new_n229_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n222_), .A2(KEYINPUT82), .A3(new_n229_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n280_), .A2(new_n284_), .ZN(new_n371_));
  OAI22_X1  g170(.A1(new_n369_), .A2(new_n370_), .B1(new_n371_), .B2(new_n273_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n350_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n368_), .A2(new_n372_), .A3(KEYINPUT20), .A4(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n366_), .A2(new_n367_), .A3(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G8gat), .B(G36gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT18), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n375_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n366_), .A2(KEYINPUT97), .A3(new_n374_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n372_), .A2(KEYINPUT20), .ZN(new_n385_));
  INV_X1    g184(.A(new_n368_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n350_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n365_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n388_), .A2(KEYINPUT20), .A3(new_n373_), .A4(new_n351_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n384_), .A2(new_n381_), .A3(new_n387_), .A4(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n250_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n318_), .A2(new_n391_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n250_), .B(new_n305_), .C1(new_n315_), .C2(new_n317_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(KEYINPUT95), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT95), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n331_), .A2(new_n395_), .A3(new_n305_), .A4(new_n250_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(KEYINPUT4), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n392_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n401_), .B(KEYINPUT96), .Z(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G85gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT0), .B(G57gat), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n405_), .B(new_n406_), .Z(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n394_), .A2(new_n396_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n402_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n403_), .A2(KEYINPUT98), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT98), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n410_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n407_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n410_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n413_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n412_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n403_), .A2(new_n414_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n408_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n383_), .A2(new_n390_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n366_), .A2(new_n374_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n379_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n366_), .A2(new_n380_), .A3(new_n374_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n403_), .A2(KEYINPUT33), .A3(new_n411_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n400_), .A2(new_n410_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n407_), .B1(new_n409_), .B2(new_n402_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n426_), .A2(new_n428_), .A3(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n425_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n348_), .B1(new_n421_), .B2(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n418_), .A2(new_n420_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n348_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT27), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n366_), .A2(new_n380_), .A3(new_n374_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n380_), .B1(new_n366_), .B2(new_n374_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n352_), .A2(new_n365_), .A3(new_n350_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT20), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n234_), .B2(new_n286_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n373_), .B1(new_n443_), .B2(new_n368_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n379_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(KEYINPUT27), .A3(new_n424_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n435_), .A2(new_n436_), .A3(new_n440_), .A4(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n254_), .B1(new_n434_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n435_), .A2(new_n254_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n440_), .A2(new_n348_), .A3(new_n446_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT99), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n348_), .A2(new_n440_), .A3(new_n446_), .A4(KEYINPUT99), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n449_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT13), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G230gat), .A2(G233gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G99gat), .A2(G106gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT6), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n461_), .A2(KEYINPUT65), .ZN(new_n462_));
  OR3_X1    g261(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(KEYINPUT65), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n460_), .A2(new_n462_), .A3(new_n463_), .A4(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G85gat), .B(G92gat), .Z(new_n466_));
  INV_X1    g265(.A(KEYINPUT66), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT8), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT66), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G57gat), .B(G64gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT11), .ZN(new_n476_));
  XOR2_X1   g275(.A(G71gat), .B(G78gat), .Z(new_n477_));
  OR2_X1    g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n477_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n475_), .A2(KEYINPUT11), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G85gat), .ZN(new_n482_));
  INV_X1    g281(.A(G92gat), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n482_), .A2(new_n483_), .A3(KEYINPUT9), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(new_n466_), .B2(KEYINPUT9), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT64), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT10), .B(G99gat), .Z(new_n487_));
  INV_X1    g286(.A(G106gat), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n486_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT10), .B(G99gat), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n490_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n460_), .B(new_n485_), .C1(new_n489_), .C2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n465_), .A2(new_n472_), .A3(new_n469_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n474_), .A2(new_n481_), .A3(new_n492_), .A4(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT68), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n474_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(new_n481_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n458_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n494_), .A2(new_n457_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n481_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT12), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n492_), .A2(new_n493_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n472_), .B1(new_n465_), .B2(new_n469_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n502_), .B(new_n503_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n503_), .B1(new_n497_), .B2(new_n502_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n501_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G120gat), .B(G148gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G176gat), .B(G204gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n500_), .A2(new_n509_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n515_), .B1(new_n500_), .B2(new_n509_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n456_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n518_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(KEYINPUT13), .A3(new_n516_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G113gat), .B(G141gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G169gat), .B(G197gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526_));
  INV_X1    g325(.A(G1gat), .ZN(new_n527_));
  INV_X1    g326(.A(G8gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G1gat), .B(G8gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G29gat), .B(G36gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT77), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n532_), .A2(new_n536_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n532_), .A2(new_n536_), .A3(KEYINPUT77), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G229gat), .A2(G233gat), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n535_), .B(KEYINPUT15), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n532_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(new_n543_), .A3(new_n537_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT78), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n525_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n525_), .ZN(new_n551_));
  AOI211_X1 g350(.A(KEYINPUT78), .B(new_n551_), .C1(new_n544_), .C2(new_n547_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n522_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n455_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n497_), .A2(new_n545_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n497_), .A2(new_n536_), .ZN(new_n562_));
  OAI211_X1 g361(.A(KEYINPUT35), .B(new_n559_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G190gat), .B(G218gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT71), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT36), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT72), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n498_), .A2(new_n535_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n560_), .A4(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n563_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n563_), .A2(new_n575_), .A3(KEYINPUT73), .A4(new_n571_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n567_), .A2(new_n568_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n569_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n563_), .B2(new_n575_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT74), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n586_), .A3(KEYINPUT37), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n583_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT37), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT74), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n584_), .A2(KEYINPUT75), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT75), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n583_), .A2(new_n592_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n580_), .A2(new_n591_), .A3(new_n589_), .A4(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n587_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n532_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(new_n502_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(G127gat), .B(G155gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT16), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT17), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n605_), .A2(KEYINPUT76), .ZN(new_n606_));
  OR3_X1    g405(.A1(new_n600_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n605_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n600_), .B(new_n608_), .C1(new_n604_), .C2(new_n606_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n596_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n556_), .A2(new_n612_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n613_), .A2(G1gat), .A3(new_n435_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n614_), .A2(KEYINPUT38), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(KEYINPUT38), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n452_), .A2(new_n453_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n449_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n254_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n384_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n387_), .A2(new_n389_), .A3(new_n381_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n383_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n418_), .A2(new_n420_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n438_), .A2(new_n439_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n626_), .A2(new_n426_), .A3(new_n431_), .A4(new_n428_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n436_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n440_), .A2(new_n446_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n338_), .A2(new_n342_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT93), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n632_), .A2(new_n418_), .A3(new_n343_), .A4(new_n420_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n629_), .A2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n620_), .B1(new_n628_), .B2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n619_), .A2(new_n635_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n580_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n555_), .A2(new_n611_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n636_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G1gat), .B1(new_n640_), .B2(new_n435_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n615_), .A2(new_n616_), .A3(new_n641_), .ZN(G1324gat));
  NOR2_X1   g441(.A1(new_n455_), .A2(new_n637_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n629_), .A3(new_n639_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .A4(G8gat), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n528_), .B1(KEYINPUT100), .B2(KEYINPUT39), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n644_), .A2(new_n649_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n629_), .A2(new_n528_), .ZN(new_n651_));
  OAI22_X1  g450(.A1(new_n648_), .A2(new_n650_), .B1(new_n613_), .B2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g452(.A(G15gat), .B1(new_n640_), .B2(new_n620_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(KEYINPUT102), .B(G15gat), .C1(new_n640_), .C2(new_n620_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  OR3_X1    g460(.A1(new_n613_), .A2(G15gat), .A3(new_n620_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n656_), .A2(new_n659_), .A3(new_n657_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT103), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n661_), .A2(new_n666_), .A3(new_n662_), .A4(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1326gat));
  OAI21_X1  g467(.A(G22gat), .B1(new_n640_), .B2(new_n348_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT42), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n348_), .A2(G22gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n613_), .B2(new_n671_), .ZN(G1327gat));
  NOR2_X1   g471(.A1(new_n555_), .A2(new_n610_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n636_), .B2(new_n596_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n674_), .B(new_n596_), .C1(new_n448_), .C2(new_n454_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  OAI211_X1 g476(.A(KEYINPUT44), .B(new_n673_), .C1(new_n675_), .C2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n673_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT43), .B1(new_n455_), .B2(new_n595_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n680_), .B2(new_n676_), .ZN(new_n681_));
  XOR2_X1   g480(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(G29gat), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n683_), .A2(new_n684_), .A3(new_n435_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n638_), .A2(new_n610_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n636_), .A2(new_n554_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G29gat), .B1(new_n688_), .B2(new_n624_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n685_), .A2(new_n689_), .ZN(G1328gat));
  XNOR2_X1  g489(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n691_));
  INV_X1    g490(.A(new_n629_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n692_), .A2(G36gat), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n687_), .A2(new_n691_), .A3(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n691_), .B1(new_n687_), .B2(new_n693_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n678_), .B(new_n629_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(G36gat), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n699_), .A2(new_n700_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n698_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n701_), .A2(new_n704_), .ZN(G1329gat));
  NAND2_X1  g504(.A1(new_n254_), .A2(G43gat), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n687_), .A2(new_n620_), .ZN(new_n707_));
  OAI22_X1  g506(.A1(new_n683_), .A2(new_n706_), .B1(G43gat), .B2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g508(.A(G50gat), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n683_), .A2(new_n710_), .A3(new_n348_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G50gat), .B1(new_n688_), .B2(new_n436_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1331gat));
  INV_X1    g512(.A(new_n522_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n550_), .A2(new_n552_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n643_), .A2(new_n610_), .A3(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n435_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n636_), .A2(new_n716_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n612_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n435_), .A2(G57gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n720_), .B2(new_n721_), .ZN(G1332gat));
  OR3_X1    g521(.A1(new_n720_), .A2(G64gat), .A3(new_n692_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n717_), .A2(new_n692_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(G64gat), .ZN(new_n726_));
  OAI211_X1 g525(.A(G64gat), .B(new_n724_), .C1(new_n717_), .C2(new_n692_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n723_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT108), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n731_), .B(new_n723_), .C1(new_n726_), .C2(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1333gat));
  OAI21_X1  g532(.A(G71gat), .B1(new_n717_), .B2(new_n620_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT49), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n736_), .B(G71gat), .C1(new_n717_), .C2(new_n620_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  OR3_X1    g537(.A1(new_n720_), .A2(G71gat), .A3(new_n620_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n738_), .A2(KEYINPUT109), .A3(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1334gat));
  OAI21_X1  g543(.A(G78gat), .B1(new_n717_), .B2(new_n348_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT50), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n348_), .A2(G78gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n720_), .B2(new_n747_), .ZN(G1335gat));
  NAND2_X1  g547(.A1(new_n719_), .A2(new_n686_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n482_), .B1(new_n749_), .B2(new_n435_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT110), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n716_), .A2(new_n611_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n680_), .B2(new_n676_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n435_), .A2(new_n482_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n751_), .B1(new_n753_), .B2(new_n754_), .ZN(G1336gat));
  AND2_X1   g554(.A1(new_n753_), .A2(new_n629_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n629_), .A2(new_n483_), .ZN(new_n757_));
  OAI22_X1  g556(.A1(new_n756_), .A2(new_n483_), .B1(new_n749_), .B2(new_n757_), .ZN(G1337gat));
  AND4_X1   g557(.A1(new_n487_), .A2(new_n719_), .A3(new_n254_), .A4(new_n686_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n753_), .A2(new_n254_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(G99gat), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT111), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT51), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n761_), .B2(KEYINPUT111), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n763_), .B2(new_n766_), .ZN(G1338gat));
  INV_X1    g566(.A(new_n752_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n436_), .B(new_n768_), .C1(new_n675_), .C2(new_n677_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G106gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G106gat), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n436_), .A2(new_n488_), .ZN(new_n773_));
  OAI22_X1  g572(.A1(new_n771_), .A2(new_n772_), .B1(new_n749_), .B2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g574(.A(G113gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n617_), .A2(new_n624_), .A3(new_n254_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n507_), .A2(new_n508_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n458_), .B1(new_n778_), .B2(new_n496_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT55), .B(new_n501_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n509_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(new_n780_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n514_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT56), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(new_n786_), .A3(new_n514_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n785_), .A2(new_n516_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n543_), .B1(new_n546_), .B2(new_n537_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n790_));
  MUX2_X1   g589(.A(new_n790_), .B(new_n548_), .S(new_n525_), .Z(new_n791_));
  NAND4_X1  g590(.A1(new_n788_), .A2(KEYINPUT115), .A3(KEYINPUT58), .A4(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n785_), .A2(new_n791_), .A3(new_n516_), .A4(new_n787_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT114), .B(KEYINPUT58), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n792_), .A2(new_n596_), .A3(new_n796_), .A4(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n785_), .A2(new_n715_), .A3(new_n516_), .A4(new_n787_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n791_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT57), .B1(new_n802_), .B2(new_n638_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  AOI211_X1 g604(.A(new_n805_), .B(new_n637_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n799_), .A2(new_n804_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n611_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n522_), .A2(new_n715_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n595_), .A2(new_n811_), .A3(new_n610_), .ZN(new_n812_));
  XOR2_X1   g611(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n812_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n809_), .A2(new_n810_), .A3(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n803_), .A2(new_n806_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n610_), .B1(new_n819_), .B2(new_n799_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT116), .B1(new_n820_), .B2(new_n816_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n777_), .B1(new_n818_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT117), .B(new_n776_), .C1(new_n823_), .C2(new_n553_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n553_), .B(new_n777_), .C1(new_n818_), .C2(new_n821_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(G113gat), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n809_), .A2(new_n817_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n777_), .ZN(new_n829_));
  XOR2_X1   g628(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n830_));
  NAND3_X1  g629(.A1(new_n828_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n822_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n553_), .A2(new_n776_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n824_), .A2(new_n827_), .B1(new_n834_), .B2(new_n835_), .ZN(G1340gat));
  OAI21_X1  g635(.A(G120gat), .B1(new_n833_), .B2(new_n714_), .ZN(new_n837_));
  INV_X1    g636(.A(G120gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n714_), .B2(KEYINPUT60), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n822_), .B(new_n839_), .C1(KEYINPUT60), .C2(new_n838_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(G1341gat));
  OAI21_X1  g640(.A(G127gat), .B1(new_n833_), .B2(new_n611_), .ZN(new_n842_));
  OR3_X1    g641(.A1(new_n823_), .A2(G127gat), .A3(new_n611_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1342gat));
  OAI21_X1  g643(.A(G134gat), .B1(new_n833_), .B2(new_n595_), .ZN(new_n845_));
  OR3_X1    g644(.A1(new_n823_), .A2(G134gat), .A3(new_n638_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1343gat));
  NAND3_X1  g646(.A1(new_n620_), .A2(new_n436_), .A3(new_n624_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n629_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n818_), .B2(new_n821_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n715_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT119), .B(G141gat), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1344gat));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n522_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g655(.A(KEYINPUT61), .B(G155gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n851_), .A2(new_n859_), .A3(new_n610_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n851_), .B2(new_n610_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n858_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n818_), .A2(new_n821_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(new_n610_), .A3(new_n849_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT120), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n851_), .A2(new_n859_), .A3(new_n610_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n857_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n862_), .A2(new_n867_), .ZN(G1346gat));
  AOI211_X1 g667(.A(new_n638_), .B(new_n850_), .C1(new_n818_), .C2(new_n821_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT121), .B1(new_n869_), .B2(G162gat), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n851_), .A2(new_n637_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872_));
  INV_X1    g671(.A(G162gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n595_), .A2(new_n873_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT122), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n870_), .A2(new_n874_), .B1(new_n851_), .B2(new_n876_), .ZN(G1347gat));
  NAND2_X1  g676(.A1(new_n618_), .A2(new_n629_), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(KEYINPUT123), .Z(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n436_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n828_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n715_), .ZN(new_n883_));
  XOR2_X1   g682(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n884_));
  AND3_X1   g683(.A1(new_n883_), .A2(G169gat), .A3(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n883_), .B2(G169gat), .ZN(new_n886_));
  INV_X1    g685(.A(new_n882_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT22), .B(G169gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n715_), .A2(new_n888_), .ZN(new_n889_));
  XOR2_X1   g688(.A(new_n889_), .B(KEYINPUT125), .Z(new_n890_));
  OAI22_X1  g689(.A1(new_n885_), .A2(new_n886_), .B1(new_n887_), .B2(new_n890_), .ZN(G1348gat));
  AOI21_X1  g690(.A(G176gat), .B1(new_n882_), .B2(new_n522_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n436_), .B1(new_n818_), .B2(new_n821_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n879_), .A2(G176gat), .A3(new_n522_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1349gat));
  NOR3_X1   g694(.A1(new_n887_), .A2(new_n611_), .A3(new_n206_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n893_), .A2(new_n610_), .A3(new_n879_), .ZN(new_n897_));
  INV_X1    g696(.A(G183gat), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n896_), .B1(new_n897_), .B2(new_n898_), .ZN(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n887_), .B2(new_n595_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n882_), .A2(new_n637_), .A3(new_n210_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1351gat));
  NOR3_X1   g701(.A1(new_n692_), .A2(new_n254_), .A3(new_n633_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n863_), .A2(new_n715_), .A3(new_n903_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g704(.A1(new_n863_), .A2(new_n522_), .A3(new_n903_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n281_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n263_), .B2(new_n906_), .ZN(G1353gat));
  AND2_X1   g707(.A1(new_n863_), .A2(new_n903_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n611_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT126), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n911_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n909_), .A2(new_n910_), .A3(new_n913_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1354gat));
  AOI21_X1  g716(.A(G218gat), .B1(new_n909_), .B2(new_n637_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n596_), .A2(G218gat), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(KEYINPUT127), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n909_), .B2(new_n920_), .ZN(G1355gat));
endmodule


