//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n814_;
  INV_X1    g000(.A(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT26), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT77), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT25), .B(G183gat), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n202_), .A2(KEYINPUT26), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(KEYINPUT77), .ZN(new_n207_));
  NAND4_X1  g006(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .A4(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT78), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT23), .ZN(new_n216_));
  OR3_X1    g015(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n208_), .A2(new_n214_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n216_), .B1(G183gat), .B2(G190gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT79), .B(G176gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT22), .B(G169gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n224_), .A2(new_n211_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n219_), .A2(new_n220_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n218_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT30), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  INV_X1    g030(.A(G15gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(G43gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G71gat), .B(G99gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n234_), .B(new_n235_), .Z(new_n236_));
  NAND3_X1  g035(.A1(new_n229_), .A2(new_n230_), .A3(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n230_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n237_), .B(KEYINPUT83), .C1(new_n229_), .C2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n241_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(KEYINPUT82), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT82), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n240_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n247_), .B(KEYINPUT31), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n239_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n225_), .A2(new_n219_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT92), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n206_), .A2(new_n203_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n205_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n213_), .A2(new_n209_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G211gat), .B(G218gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(G197gat), .B(G204gat), .Z(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(KEYINPUT90), .ZN(new_n259_));
  INV_X1    g058(.A(G197gat), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n260_), .A2(G204gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT90), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT21), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  OAI221_X1 g062(.A(new_n257_), .B1(KEYINPUT21), .B2(new_n258_), .C1(new_n259_), .C2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n258_), .A2(KEYINPUT21), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(new_n257_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n256_), .A2(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n228_), .A2(new_n266_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(KEYINPUT20), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT19), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n228_), .A2(new_n266_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n273_), .A2(new_n274_), .A3(new_n271_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(new_n266_), .B2(new_n256_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G64gat), .B(G92gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT94), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G8gat), .B(G36gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n277_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n272_), .A2(new_n276_), .A3(new_n283_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT27), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n255_), .A2(new_n250_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT20), .B1(new_n266_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n271_), .B1(new_n273_), .B2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n284_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(KEYINPUT27), .A3(new_n286_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n289_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT86), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT3), .ZN(new_n300_));
  AND2_X1   g099(.A1(G141gat), .A2(G148gat), .ZN(new_n301_));
  OR2_X1    g100(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n302_));
  NAND2_X1  g101(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n298_), .B(new_n300_), .C1(new_n301_), .C2(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT84), .ZN(new_n309_));
  OR3_X1    g108(.A1(new_n307_), .A2(new_n309_), .A3(KEYINPUT1), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n309_), .B1(new_n307_), .B2(KEYINPUT1), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(KEYINPUT1), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .A4(new_n306_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G141gat), .B(G148gat), .Z(new_n314_));
  AOI22_X1  g113(.A1(new_n305_), .A2(new_n308_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(G22gat), .B(G50gat), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT89), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n266_), .B(new_n322_), .C1(new_n316_), .C2(new_n315_), .ZN(new_n323_));
  INV_X1    g122(.A(G233gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT88), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(G228gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(G228gat), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n324_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n323_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT91), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n321_), .A2(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G78gat), .B(G106gat), .Z(new_n333_));
  AND2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n332_), .A2(new_n333_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n330_), .A2(KEYINPUT91), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  OR3_X1    g136(.A1(new_n334_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n337_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n296_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT96), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n249_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n247_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(new_n315_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n344_), .A2(KEYINPUT4), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n242_), .A2(new_n243_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n315_), .A2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n343_), .B2(new_n315_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n345_), .B1(new_n348_), .B2(KEYINPUT4), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT95), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n351_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G85gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT0), .B(G57gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n357_), .B(new_n358_), .Z(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n359_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n352_), .A2(new_n361_), .A3(new_n354_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n338_), .A2(new_n339_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(KEYINPUT96), .A3(new_n296_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n342_), .A2(new_n364_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT97), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n342_), .A2(KEYINPUT97), .A3(new_n367_), .A4(new_n364_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n365_), .A2(new_n364_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n296_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n360_), .B(KEYINPUT33), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n361_), .B1(new_n348_), .B2(new_n353_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n349_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(new_n353_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n287_), .A2(new_n377_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n283_), .A2(KEYINPUT32), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n277_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n293_), .B2(new_n379_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n374_), .A2(new_n378_), .B1(new_n381_), .B2(new_n363_), .ZN(new_n382_));
  OAI22_X1  g181(.A1(new_n372_), .A2(new_n373_), .B1(new_n382_), .B2(new_n365_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n370_), .A2(new_n371_), .B1(new_n383_), .B2(new_n249_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G29gat), .B(G36gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G43gat), .B(G50gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT75), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G15gat), .B(G22gat), .ZN(new_n389_));
  INV_X1    g188(.A(G1gat), .ZN(new_n390_));
  INV_X1    g189(.A(G8gat), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT14), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G1gat), .B(G8gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n388_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT76), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n388_), .A2(new_n395_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n387_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n397_), .B1(new_n395_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G229gat), .A2(G233gat), .ZN(new_n404_));
  MUX2_X1   g203(.A(new_n399_), .B(new_n403_), .S(new_n404_), .Z(new_n405_));
  XOR2_X1   g204(.A(G113gat), .B(G141gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(G169gat), .B(G197gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n408_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n384_), .A2(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(G230gat), .A2(G233gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(G85gat), .B(G92gat), .Z(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT9), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G99gat), .A2(G106gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT6), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(G99gat), .A3(G106gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G85gat), .ZN(new_n422_));
  INV_X1    g221(.A(G92gat), .ZN(new_n423_));
  OR3_X1    g222(.A1(new_n422_), .A2(new_n423_), .A3(KEYINPUT9), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n416_), .A2(new_n421_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G106gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT10), .B(G99gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT64), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n425_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n430_));
  INV_X1    g229(.A(G99gat), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n426_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT7), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT7), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n430_), .A2(new_n434_), .A3(new_n431_), .A4(new_n426_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n421_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n415_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT8), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT8), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(new_n439_), .A3(new_n415_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n429_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G57gat), .B(G64gat), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n442_), .A2(KEYINPUT11), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(KEYINPUT11), .ZN(new_n444_));
  XOR2_X1   g243(.A(G71gat), .B(G78gat), .Z(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n441_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT66), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n449_), .A2(KEYINPUT66), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n441_), .A2(new_n447_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n414_), .B(new_n450_), .C1(new_n451_), .C2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT12), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n447_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n436_), .A2(new_n439_), .A3(new_n415_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n439_), .B1(new_n436_), .B2(new_n415_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n458_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n438_), .A2(KEYINPUT67), .A3(new_n440_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n429_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT68), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT68), .ZN(new_n466_));
  AOI211_X1 g265(.A(new_n466_), .B(new_n429_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n457_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n448_), .A2(new_n455_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n414_), .B1(new_n441_), .B2(new_n447_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n454_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G120gat), .B(G148gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT5), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G176gat), .B(G204gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n476_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n454_), .A2(new_n471_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT13), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n477_), .A2(KEYINPUT13), .A3(new_n479_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT69), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n447_), .B(new_n395_), .Z(new_n487_));
  NAND2_X1  g286(.A1(G231gat), .A2(G233gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G127gat), .B(G155gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G183gat), .B(G211gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT17), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n489_), .A2(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n494_), .A2(KEYINPUT17), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n489_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n401_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT35), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G232gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT34), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n441_), .A2(new_n387_), .B1(new_n502_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n501_), .A2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n505_), .A2(new_n502_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n507_), .A2(new_n508_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G190gat), .B(G218gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT71), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G134gat), .B(G162gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n512_), .B(new_n513_), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  OR4_X1    g314(.A1(KEYINPUT36), .A2(new_n509_), .A3(new_n510_), .A4(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n514_), .B(KEYINPUT36), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(KEYINPUT72), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT72), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n523_), .B1(new_n519_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n413_), .A2(new_n486_), .A3(new_n500_), .A4(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n528_), .B(KEYINPUT98), .Z(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(new_n390_), .A3(new_n363_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT38), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n484_), .A2(new_n412_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NOR4_X1   g333(.A1(new_n384_), .A2(new_n499_), .A3(new_n520_), .A4(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n390_), .B1(new_n535_), .B2(new_n363_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n531_), .B2(new_n530_), .ZN(G1324gat));
  NAND3_X1  g337(.A1(new_n529_), .A2(new_n391_), .A3(new_n373_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n535_), .A2(new_n373_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT99), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(KEYINPUT39), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n391_), .B1(new_n541_), .B2(KEYINPUT39), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n540_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n542_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n539_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g346(.A(new_n249_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n232_), .B1(new_n535_), .B2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT41), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n232_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n550_), .B1(new_n528_), .B2(new_n551_), .ZN(G1326gat));
  INV_X1    g351(.A(G22gat), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n535_), .B2(new_n365_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n554_), .B(KEYINPUT42), .Z(new_n555_));
  NAND2_X1  g354(.A1(new_n365_), .A2(new_n553_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n555_), .B1(new_n528_), .B2(new_n556_), .ZN(G1327gat));
  NOR2_X1   g356(.A1(new_n519_), .A2(new_n500_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(new_n484_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n413_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(G29gat), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n563_), .A3(new_n363_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT101), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n370_), .A2(new_n371_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n383_), .A2(new_n249_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT43), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n526_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT43), .B1(new_n384_), .B2(new_n527_), .ZN(new_n571_));
  AOI211_X1 g370(.A(new_n500_), .B(new_n534_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT100), .B(KEYINPUT44), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n571_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n575_), .A2(KEYINPUT44), .A3(new_n499_), .A4(new_n533_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n363_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n565_), .B1(new_n578_), .B2(G29gat), .ZN(new_n579_));
  AOI211_X1 g378(.A(KEYINPUT101), .B(new_n563_), .C1(new_n577_), .C2(new_n363_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n564_), .B1(new_n579_), .B2(new_n580_), .ZN(G1328gat));
  INV_X1    g380(.A(KEYINPUT104), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n296_), .A2(G36gat), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n413_), .A2(new_n560_), .A3(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n576_), .B(new_n373_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n586_), .B1(new_n587_), .B2(G36gat), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT103), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT46), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n582_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n587_), .A2(G36gat), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT103), .B1(new_n595_), .B2(new_n586_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n596_), .A2(KEYINPUT104), .A3(new_n592_), .A4(new_n590_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n588_), .A2(KEYINPUT46), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n594_), .A2(new_n597_), .A3(new_n598_), .ZN(G1329gat));
  NAND4_X1  g398(.A1(new_n574_), .A2(G43gat), .A3(new_n548_), .A4(new_n576_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n561_), .A2(new_n249_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n600_), .B1(G43gat), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g402(.A(G50gat), .B1(new_n562_), .B2(new_n365_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n365_), .A2(G50gat), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n577_), .B2(new_n605_), .ZN(G1331gat));
  NOR2_X1   g405(.A1(new_n411_), .A2(new_n499_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n568_), .A2(new_n485_), .A3(new_n519_), .A4(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G57gat), .B1(new_n608_), .B2(new_n364_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n527_), .A2(new_n484_), .A3(new_n500_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n384_), .A2(new_n411_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(G57gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n363_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(new_n613_), .ZN(G1332gat));
  OAI21_X1  g413(.A(G64gat), .B1(new_n608_), .B2(new_n296_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT105), .B(KEYINPUT48), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(G64gat), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n611_), .A2(new_n618_), .A3(new_n373_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(G1333gat));
  OAI21_X1  g419(.A(G71gat), .B1(new_n608_), .B2(new_n249_), .ZN(new_n621_));
  XOR2_X1   g420(.A(KEYINPUT106), .B(KEYINPUT49), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(G71gat), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n611_), .A2(new_n624_), .A3(new_n548_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(G1334gat));
  OAI21_X1  g425(.A(G78gat), .B1(new_n608_), .B2(new_n366_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT50), .ZN(new_n628_));
  INV_X1    g427(.A(G78gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n611_), .A2(new_n629_), .A3(new_n365_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(G1335gat));
  NOR2_X1   g430(.A1(new_n486_), .A2(new_n559_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n568_), .A2(new_n412_), .A3(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n422_), .B1(new_n633_), .B2(new_n364_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT107), .Z(new_n635_));
  INV_X1    g434(.A(new_n484_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n636_), .A2(new_n411_), .A3(new_n500_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n575_), .A2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(new_n422_), .A3(new_n364_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n635_), .A2(new_n639_), .ZN(G1336gat));
  OAI21_X1  g439(.A(new_n423_), .B1(new_n633_), .B2(new_n296_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT108), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n638_), .A2(new_n423_), .A3(new_n296_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1337gat));
  INV_X1    g443(.A(new_n633_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n548_), .A3(new_n428_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n575_), .A2(new_n548_), .A3(new_n637_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G99gat), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT109), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(KEYINPUT109), .A3(G99gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n647_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n654_), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT111), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT51), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n653_), .B2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT110), .B1(new_n654_), .B2(KEYINPUT51), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT110), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n653_), .A2(new_n660_), .A3(new_n657_), .ZN(new_n661_));
  OAI22_X1  g460(.A1(new_n655_), .A2(new_n658_), .B1(new_n659_), .B2(new_n661_), .ZN(G1338gat));
  NAND3_X1  g461(.A1(new_n645_), .A2(new_n426_), .A3(new_n365_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G106gat), .B1(new_n638_), .B2(new_n366_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(KEYINPUT52), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(KEYINPUT52), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n663_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT53), .ZN(G1339gat));
  AND2_X1   g467(.A1(new_n342_), .A2(new_n367_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n363_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n468_), .A2(new_n469_), .A3(new_n452_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n471_), .A2(KEYINPUT55), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT55), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n468_), .A2(new_n673_), .A3(new_n469_), .A4(new_n470_), .ZN(new_n674_));
  AOI221_X4 g473(.A(KEYINPUT113), .B1(new_n671_), .B2(new_n414_), .C1(new_n672_), .C2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT113), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n672_), .A2(new_n674_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n671_), .A2(new_n414_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n676_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n476_), .B1(new_n675_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT114), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT56), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n680_), .A2(KEYINPUT114), .A3(KEYINPUT56), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n683_), .A2(new_n411_), .A3(new_n479_), .A4(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n397_), .A2(new_n398_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n408_), .B1(new_n686_), .B2(new_n404_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n687_), .B1(new_n404_), .B2(new_n403_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n410_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n480_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT115), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n520_), .B1(new_n685_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT57), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n680_), .A2(new_n682_), .ZN(new_n695_));
  OAI211_X1 g494(.A(KEYINPUT56), .B(new_n476_), .C1(new_n675_), .C2(new_n679_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n695_), .A2(KEYINPUT116), .A3(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n689_), .A2(new_n479_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT116), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n680_), .A2(new_n699_), .A3(new_n682_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT117), .B1(new_n697_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT58), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n695_), .A2(KEYINPUT116), .A3(new_n696_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT117), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n700_), .A4(new_n698_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n702_), .A2(new_n703_), .A3(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(KEYINPUT118), .A3(new_n526_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n704_), .A2(KEYINPUT58), .A3(new_n700_), .A4(new_n698_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT118), .B1(new_n707_), .B2(new_n526_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n694_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT119), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT119), .B(new_n694_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n499_), .A3(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n527_), .A2(new_n636_), .A3(new_n607_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n670_), .B1(new_n716_), .B2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G113gat), .B1(new_n721_), .B2(new_n411_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n721_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT59), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n670_), .A2(KEYINPUT59), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n712_), .A2(new_n499_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(new_n719_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(G113gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n411_), .B2(KEYINPUT120), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(KEYINPUT120), .B2(new_n729_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n722_), .B1(new_n728_), .B2(new_n731_), .ZN(G1340gat));
  NAND3_X1  g531(.A1(new_n724_), .A2(new_n485_), .A3(new_n727_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(G120gat), .ZN(new_n734_));
  INV_X1    g533(.A(G120gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n735_), .B1(new_n636_), .B2(KEYINPUT60), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(KEYINPUT60), .B2(new_n735_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n734_), .B1(new_n723_), .B2(new_n737_), .ZN(G1341gat));
  NAND3_X1  g537(.A1(new_n724_), .A2(new_n500_), .A3(new_n727_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G127gat), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n499_), .A2(G127gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n740_), .B1(new_n723_), .B2(new_n741_), .ZN(G1342gat));
  INV_X1    g541(.A(KEYINPUT59), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n526_), .B(new_n727_), .C1(new_n721_), .C2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G134gat), .ZN(new_n745_));
  INV_X1    g544(.A(G134gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n721_), .A2(new_n746_), .A3(new_n520_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT121), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT121), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n745_), .A2(new_n750_), .A3(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1343gat));
  NAND3_X1  g551(.A1(new_n365_), .A2(new_n363_), .A3(new_n249_), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n373_), .B(new_n753_), .C1(new_n716_), .C2(new_n720_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n411_), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT122), .B(G141gat), .Z(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(G1344gat));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n485_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(KEYINPUT123), .B(G148gat), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(G1345gat));
  NAND2_X1  g559(.A1(new_n754_), .A2(new_n500_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT61), .B(G155gat), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(G1346gat));
  INV_X1    g562(.A(G162gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n754_), .A2(new_n764_), .A3(new_n520_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n754_), .A2(new_n526_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n764_), .ZN(G1347gat));
  INV_X1    g566(.A(KEYINPUT62), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n373_), .A2(new_n364_), .A3(new_n548_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n366_), .B(new_n770_), .C1(new_n726_), .C2(new_n719_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n412_), .ZN(new_n772_));
  INV_X1    g571(.A(G169gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n768_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n223_), .ZN(new_n775_));
  OAI211_X1 g574(.A(KEYINPUT62), .B(G169gat), .C1(new_n771_), .C2(new_n412_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(new_n775_), .A3(new_n776_), .ZN(G1348gat));
  OAI21_X1  g576(.A(new_n222_), .B1(new_n771_), .B2(new_n636_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n716_), .A2(new_n720_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n366_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n485_), .A2(G176gat), .A3(new_n770_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT124), .ZN(G1349gat));
  NOR3_X1   g582(.A1(new_n771_), .A2(new_n205_), .A3(new_n499_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n779_), .A2(new_n366_), .A3(new_n500_), .A4(new_n770_), .ZN(new_n785_));
  INV_X1    g584(.A(G183gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(G1350gat));
  OAI21_X1  g586(.A(G190gat), .B1(new_n771_), .B2(new_n527_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT125), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n788_), .A2(new_n789_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n520_), .A2(new_n252_), .ZN(new_n792_));
  OAI22_X1  g591(.A1(new_n790_), .A2(new_n791_), .B1(new_n771_), .B2(new_n792_), .ZN(G1351gat));
  NOR3_X1   g592(.A1(new_n372_), .A2(new_n296_), .A3(new_n548_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n779_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT126), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n779_), .A2(KEYINPUT126), .A3(new_n794_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n412_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(new_n260_), .ZN(G1352gat));
  AOI21_X1  g599(.A(new_n486_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n801_));
  AND2_X1   g600(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n802_));
  NOR2_X1   g601(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n801_), .B2(new_n803_), .ZN(G1353gat));
  AOI21_X1  g604(.A(new_n499_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n807_));
  AND2_X1   g606(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n806_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n806_), .B2(new_n807_), .ZN(G1354gat));
  NAND2_X1  g609(.A1(new_n797_), .A2(new_n798_), .ZN(new_n811_));
  INV_X1    g610(.A(G218gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n520_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n527_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n812_), .B2(new_n814_), .ZN(G1355gat));
endmodule


