//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_;
  XNOR2_X1  g000(.A(KEYINPUT71), .B(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G8gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G36gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G29gat), .ZN(new_n213_));
  INV_X1    g012(.A(G29gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G36gat), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n213_), .A2(new_n215_), .A3(KEYINPUT67), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT67), .B1(new_n213_), .B2(new_n215_), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n216_), .A2(new_n217_), .A3(KEYINPUT68), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n214_), .A2(G36gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n212_), .A2(G29gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n213_), .A2(new_n215_), .A3(KEYINPUT67), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n219_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n211_), .B1(new_n218_), .B2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT68), .B1(new_n216_), .B2(new_n217_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n223_), .A2(new_n219_), .A3(new_n224_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n210_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT15), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n226_), .A2(KEYINPUT15), .A3(new_n229_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n209_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n230_), .A2(new_n208_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n234_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n230_), .B(new_n208_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n238_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G113gat), .B(G141gat), .Z(new_n241_));
  XNOR2_X1  g040(.A(G169gat), .B(G197gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n240_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G99gat), .A2(G106gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT6), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT6), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(G99gat), .A3(G106gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT10), .B(G99gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G85gat), .A2(G92gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT9), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(KEYINPUT64), .A3(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(G85gat), .A2(G92gat), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n254_), .B(new_n255_), .C1(new_n253_), .C2(new_n252_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT64), .B1(new_n252_), .B2(new_n253_), .ZN(new_n257_));
  OAI221_X1 g056(.A(new_n250_), .B1(G106gat), .B2(new_n251_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(G99gat), .ZN(new_n259_));
  INV_X1    g058(.A(G106gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(new_n260_), .A3(KEYINPUT65), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT7), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT7), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n263_), .A2(new_n259_), .A3(new_n260_), .A4(KEYINPUT65), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n250_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT8), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n255_), .A2(new_n252_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n266_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n258_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G57gat), .B(G64gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G71gat), .B(G78gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT11), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(KEYINPUT11), .ZN(new_n274_));
  INV_X1    g073(.A(new_n272_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n271_), .A2(KEYINPUT11), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n273_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n270_), .A2(new_n279_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n278_), .B(new_n258_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G230gat), .A2(G233gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n265_), .A2(new_n267_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT8), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n278_), .B1(new_n289_), .B2(new_n258_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n281_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT12), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT12), .B1(new_n270_), .B2(new_n279_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n285_), .B1(new_n295_), .B2(new_n284_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G120gat), .B(G148gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT5), .ZN(new_n298_));
  XOR2_X1   g097(.A(G176gat), .B(G204gat), .Z(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n296_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT13), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n302_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G15gat), .B(G43gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT78), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT30), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT31), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT76), .ZN(new_n311_));
  INV_X1    g110(.A(G169gat), .ZN(new_n312_));
  INV_X1    g111(.A(G176gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT76), .B1(G169gat), .B2(G176gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n314_), .A2(KEYINPUT24), .A3(new_n315_), .A4(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT26), .B(G190gat), .ZN(new_n318_));
  INV_X1    g117(.A(G183gat), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT25), .B1(new_n319_), .B2(KEYINPUT75), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n319_), .A2(KEYINPUT25), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n318_), .B(new_n320_), .C1(new_n321_), .C2(KEYINPUT75), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n314_), .A2(new_n315_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT24), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT23), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n325_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n326_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n317_), .B(new_n322_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n334_));
  OR3_X1    g133(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G227gat), .A2(G233gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n338_), .B(G71gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(new_n259_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n340_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G127gat), .B(G134gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G113gat), .B(G120gat), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n344_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n343_), .B(new_n346_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n350_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n343_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(new_n348_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n341_), .A2(new_n342_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n355_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n310_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n358_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(new_n309_), .A3(new_n356_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G1gat), .B(G29gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(G85gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT0), .B(G57gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G141gat), .A2(G148gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT2), .B1(new_n369_), .B2(KEYINPUT82), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT2), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n368_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(G141gat), .A2(G148gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n370_), .A2(new_n373_), .A3(new_n376_), .A4(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n369_), .A2(new_n374_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n381_), .B1(new_n379_), .B2(KEYINPUT1), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n387_), .A2(KEYINPUT81), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n381_), .A2(KEYINPUT1), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n387_), .B2(KEYINPUT81), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n386_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n351_), .B(new_n354_), .C1(new_n384_), .C2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n344_), .A2(new_n345_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n346_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT86), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n388_), .A2(new_n390_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n385_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT86), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n346_), .A2(new_n398_), .A3(new_n393_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n395_), .A2(new_n397_), .A3(new_n383_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n392_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n392_), .A2(new_n400_), .A3(KEYINPUT4), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n397_), .A2(new_n383_), .ZN(new_n405_));
  XOR2_X1   g204(.A(KEYINPUT87), .B(KEYINPUT4), .Z(new_n406_));
  NAND4_X1  g205(.A1(new_n405_), .A2(new_n351_), .A3(new_n354_), .A4(new_n406_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n367_), .B(new_n403_), .C1(new_n408_), .C2(new_n402_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n367_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n402_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n401_), .A2(new_n402_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n410_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G78gat), .B(G106gat), .Z(new_n415_));
  NAND2_X1  g214(.A1(new_n405_), .A2(KEYINPUT29), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G228gat), .A2(G233gat), .ZN(new_n417_));
  OR2_X1    g216(.A1(G197gat), .A2(G204gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G197gat), .A2(G204gat), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(KEYINPUT21), .A4(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G211gat), .B(G218gat), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n418_), .A2(new_n420_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n421_), .B(new_n422_), .C1(new_n423_), .C2(KEYINPUT21), .ZN(new_n424_));
  XOR2_X1   g223(.A(G211gat), .B(G218gat), .Z(new_n425_));
  NAND4_X1  g224(.A1(new_n423_), .A2(new_n425_), .A3(new_n419_), .A4(KEYINPUT21), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n424_), .A2(new_n426_), .A3(KEYINPUT84), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT84), .B1(new_n424_), .B2(new_n426_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n416_), .A2(new_n417_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n424_), .A2(new_n426_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n417_), .B1(new_n416_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n415_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n415_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(new_n430_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G22gat), .B(G50gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT28), .B1(new_n405_), .B2(KEYINPUT29), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n405_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n439_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n442_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n439_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n440_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n438_), .A2(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n434_), .A2(new_n437_), .A3(new_n446_), .A4(new_n443_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n414_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT27), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT22), .B(G169gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n313_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n316_), .B(KEYINPUT85), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n333_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT25), .B(G183gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n318_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n325_), .A2(new_n328_), .A3(new_n458_), .A4(new_n317_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n452_), .B1(new_n460_), .B2(new_n432_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n337_), .B2(new_n429_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT19), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n427_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n428_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n322_), .A2(new_n317_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n325_), .A2(new_n328_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT77), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n325_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n468_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n336_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n466_), .B(new_n467_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n464_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT20), .B1(new_n460_), .B2(new_n432_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n475_), .A3(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT18), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G64gat), .B(G92gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n465_), .A2(new_n478_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n331_), .B(new_n336_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(new_n475_), .A3(new_n461_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n476_), .B1(new_n337_), .B2(new_n429_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n487_), .B1(new_n488_), .B2(new_n475_), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n484_), .A2(new_n485_), .B1(new_n489_), .B2(new_n482_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n474_), .A2(new_n475_), .A3(new_n477_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n475_), .B1(new_n486_), .B2(new_n461_), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n482_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT90), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n451_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n483_), .B1(new_n465_), .B2(new_n478_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n493_), .A2(new_n496_), .A3(KEYINPUT27), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n450_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n448_), .A2(new_n449_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n493_), .A2(new_n496_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT33), .B(new_n410_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT33), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n413_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n408_), .A2(new_n402_), .ZN(new_n504_));
  OAI211_X1 g303(.A(KEYINPUT88), .B(new_n367_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n367_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT88), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n504_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n500_), .A2(new_n501_), .A3(new_n503_), .A4(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n489_), .A2(KEYINPUT32), .A3(new_n483_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n483_), .A2(KEYINPUT32), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n465_), .A2(new_n478_), .A3(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n414_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n499_), .B1(new_n510_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT89), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n498_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  AOI211_X1 g316(.A(KEYINPUT89), .B(new_n499_), .C1(new_n510_), .C2(new_n514_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n363_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n497_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n490_), .A2(new_n494_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n521_), .B2(new_n451_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT91), .ZN(new_n523_));
  INV_X1    g322(.A(new_n499_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n414_), .B1(new_n361_), .B2(new_n359_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .A4(new_n525_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n524_), .B(new_n525_), .C1(new_n497_), .C2(new_n495_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT91), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  AOI211_X1 g328(.A(new_n245_), .B(new_n305_), .C1(new_n519_), .C2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT70), .ZN(new_n531_));
  INV_X1    g330(.A(new_n270_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT66), .B(KEYINPUT34), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G232gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT35), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n230_), .B2(new_n270_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n536_), .A2(new_n537_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n533_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n233_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT15), .B1(new_n226_), .B2(new_n229_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n270_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n539_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n542_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n531_), .B1(new_n541_), .B2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G190gat), .B(G218gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT69), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G134gat), .B(G162gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n552_), .A2(KEYINPUT36), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n553_), .B1(new_n541_), .B2(new_n547_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n552_), .A2(KEYINPUT36), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n548_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  OAI221_X1 g356(.A(new_n531_), .B1(new_n555_), .B2(new_n553_), .C1(new_n541_), .C2(new_n547_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT94), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT72), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n278_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n208_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G127gat), .B(G155gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G183gat), .B(G211gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OR3_X1    g371(.A1(new_n570_), .A2(KEYINPUT73), .A3(new_n571_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n565_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n565_), .A2(new_n573_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n561_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n530_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n414_), .ZN(new_n580_));
  OAI21_X1  g379(.A(G1gat), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n557_), .A2(KEYINPUT37), .A3(new_n558_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT37), .B1(new_n557_), .B2(new_n558_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(new_n577_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n530_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT92), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n587_), .A2(new_n202_), .A3(new_n414_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n587_), .A2(KEYINPUT38), .A3(new_n202_), .A4(new_n414_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n589_), .A2(KEYINPUT93), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(KEYINPUT93), .ZN(new_n591_));
  OAI221_X1 g390(.A(new_n581_), .B1(KEYINPUT38), .B2(new_n588_), .C1(new_n590_), .C2(new_n591_), .ZN(G1324gat));
  OAI21_X1  g391(.A(G8gat), .B1(new_n579_), .B2(new_n522_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT39), .ZN(new_n594_));
  INV_X1    g393(.A(new_n522_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n587_), .A2(new_n203_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g397(.A(G15gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n587_), .A2(new_n599_), .A3(new_n362_), .ZN(new_n600_));
  OAI21_X1  g399(.A(G15gat), .B1(new_n579_), .B2(new_n363_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT41), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(KEYINPUT41), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n600_), .A2(new_n602_), .A3(new_n603_), .ZN(G1326gat));
  OAI21_X1  g403(.A(G22gat), .B1(new_n579_), .B2(new_n524_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT42), .ZN(new_n606_));
  INV_X1    g405(.A(G22gat), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n587_), .A2(new_n607_), .A3(new_n499_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(G1327gat));
  INV_X1    g408(.A(new_n559_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n576_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n530_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(new_n214_), .A3(new_n414_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n305_), .A2(new_n576_), .A3(new_n245_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT43), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n519_), .A2(new_n529_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n616_), .B2(new_n584_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n584_), .ZN(new_n618_));
  AOI211_X1 g417(.A(KEYINPUT43), .B(new_n618_), .C1(new_n519_), .C2(new_n529_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n614_), .B1(new_n617_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT44), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  OAI211_X1 g421(.A(KEYINPUT44), .B(new_n614_), .C1(new_n617_), .C2(new_n619_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n414_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n624_), .A2(new_n625_), .A3(G29gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n624_), .B2(G29gat), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n613_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  OAI211_X1 g429(.A(KEYINPUT96), .B(new_n613_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1328gat));
  NAND3_X1  g431(.A1(new_n612_), .A2(new_n212_), .A3(new_n595_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT45), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n622_), .A2(new_n595_), .A3(new_n623_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(G36gat), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT46), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(G1329gat));
  NAND4_X1  g438(.A1(new_n622_), .A2(G43gat), .A3(new_n362_), .A4(new_n623_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n612_), .A2(new_n362_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n640_), .B1(G43gat), .B2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g442(.A1(new_n524_), .A2(G50gat), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT98), .Z(new_n645_));
  NAND2_X1  g444(.A1(new_n612_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n622_), .A2(new_n499_), .A3(new_n623_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n647_), .A2(new_n648_), .A3(G50gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n647_), .B2(G50gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(G1331gat));
  NAND2_X1  g450(.A1(new_n585_), .A2(new_n305_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT99), .Z(new_n653_));
  AOI21_X1  g452(.A(new_n244_), .B1(new_n519_), .B2(new_n529_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT100), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(G57gat), .B1(new_n657_), .B2(new_n414_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n654_), .A2(new_n305_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n659_), .A2(G57gat), .A3(new_n414_), .A4(new_n578_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT101), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n658_), .A2(new_n661_), .ZN(G1332gat));
  NAND2_X1  g461(.A1(new_n659_), .A2(new_n578_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G64gat), .B1(new_n663_), .B2(new_n522_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT48), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n522_), .A2(G64gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n656_), .B2(new_n666_), .ZN(G1333gat));
  OAI21_X1  g466(.A(G71gat), .B1(new_n663_), .B2(new_n363_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT102), .B(KEYINPUT49), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n363_), .A2(G71gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n656_), .B2(new_n671_), .ZN(G1334gat));
  OR3_X1    g471(.A1(new_n656_), .A2(G78gat), .A3(new_n524_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G78gat), .B1(new_n663_), .B2(new_n524_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT103), .B(KEYINPUT50), .Z(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n674_), .A2(new_n676_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n673_), .B1(new_n677_), .B2(new_n678_), .ZN(G1335gat));
  NAND2_X1  g478(.A1(new_n659_), .A2(new_n611_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n659_), .A2(KEYINPUT104), .A3(new_n611_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G85gat), .B1(new_n684_), .B2(new_n414_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n305_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n686_), .A2(new_n576_), .A3(new_n244_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n617_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n619_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n691_), .A2(KEYINPUT105), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(KEYINPUT105), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n414_), .A2(G85gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n685_), .B1(new_n694_), .B2(new_n695_), .ZN(G1336gat));
  AOI21_X1  g495(.A(G92gat), .B1(new_n684_), .B2(new_n595_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n595_), .A2(G92gat), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT106), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n694_), .B2(new_n699_), .ZN(G1337gat));
  INV_X1    g499(.A(new_n691_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G99gat), .B1(new_n701_), .B2(new_n363_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n363_), .A2(new_n251_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n684_), .A2(KEYINPUT107), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT107), .B1(new_n684_), .B2(new_n703_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n702_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT51), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT51), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n708_), .B(new_n702_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(G1338gat));
  OAI211_X1 g509(.A(new_n499_), .B(new_n687_), .C1(new_n617_), .C2(new_n619_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT108), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G106gat), .B1(new_n711_), .B2(KEYINPUT108), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT52), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n691_), .A2(new_n716_), .A3(new_n499_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(G106gat), .A4(new_n712_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n715_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n684_), .A2(new_n260_), .A3(new_n499_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n720_), .A2(new_n721_), .A3(new_n723_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1339gat));
  INV_X1    g526(.A(KEYINPUT116), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n240_), .A2(new_n243_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n296_), .A2(new_n300_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n243_), .B1(new_n239_), .B2(new_n235_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT114), .B1(new_n234_), .B2(new_n237_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n236_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n234_), .A2(KEYINPUT114), .A3(new_n237_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n731_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n729_), .A2(new_n730_), .A3(new_n735_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n292_), .A2(KEYINPUT55), .A3(new_n283_), .A4(new_n294_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT111), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n293_), .B1(new_n282_), .B2(KEYINPUT12), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(KEYINPUT55), .A4(new_n283_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT12), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n744_), .A2(new_n284_), .A3(new_n293_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n284_), .B1(new_n744_), .B2(new_n293_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(KEYINPUT55), .B2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n300_), .B1(new_n742_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT56), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT56), .B(new_n300_), .C1(new_n742_), .C2(new_n747_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n736_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n584_), .B1(new_n752_), .B2(KEYINPUT58), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT58), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n754_), .B(new_n736_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n728_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n751_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n295_), .B2(new_n284_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n738_), .B(new_n741_), .C1(new_n759_), .C2(new_n745_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT56), .B1(new_n760_), .B2(new_n300_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n757_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n754_), .B1(new_n762_), .B2(new_n736_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n752_), .A2(KEYINPUT58), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(KEYINPUT116), .A4(new_n584_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n756_), .A2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n301_), .A2(new_n729_), .A3(new_n735_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n750_), .A2(KEYINPUT112), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n761_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n751_), .A2(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n760_), .A2(KEYINPUT113), .A3(KEYINPUT56), .A4(new_n300_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n769_), .A2(new_n771_), .A3(new_n773_), .A4(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n244_), .A2(new_n730_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n768_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n767_), .B1(new_n778_), .B2(new_n559_), .ZN(new_n779_));
  AOI211_X1 g578(.A(KEYINPUT112), .B(KEYINPUT56), .C1(new_n760_), .C2(new_n300_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n770_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n773_), .A2(new_n774_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n776_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT57), .B(new_n610_), .C1(new_n784_), .C2(new_n768_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n766_), .A2(new_n779_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n577_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n305_), .A2(new_n244_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n585_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n788_), .A2(new_n585_), .A3(new_n790_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n787_), .A2(new_n795_), .ZN(new_n796_));
  NOR4_X1   g595(.A1(new_n595_), .A2(new_n363_), .A3(new_n499_), .A4(new_n580_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT59), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n779_), .B(new_n785_), .C1(new_n755_), .C2(new_n753_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n577_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n795_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n797_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n799_), .A2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(G113gat), .B1(new_n805_), .B2(new_n245_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n245_), .A2(G113gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n798_), .B2(new_n807_), .ZN(G1340gat));
  INV_X1    g607(.A(new_n798_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT60), .ZN(new_n810_));
  AOI21_X1  g609(.A(G120gat), .B1(new_n305_), .B2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n810_), .B2(G120gat), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT117), .ZN(new_n814_));
  OAI21_X1  g613(.A(G120gat), .B1(new_n805_), .B2(new_n686_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(G1341gat));
  INV_X1    g615(.A(G127gat), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n805_), .A2(new_n817_), .A3(new_n577_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n809_), .A2(new_n576_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT118), .B1(new_n819_), .B2(new_n817_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n821_), .B(G127gat), .C1(new_n809_), .C2(new_n576_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n818_), .A2(new_n820_), .A3(new_n822_), .ZN(G1342gat));
  OAI21_X1  g622(.A(G134gat), .B1(new_n805_), .B2(new_n618_), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n560_), .A2(G134gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n798_), .B2(new_n825_), .ZN(G1343gat));
  NOR2_X1   g625(.A1(new_n524_), .A2(new_n362_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n522_), .A3(new_n414_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n796_), .A2(KEYINPUT119), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n794_), .B1(new_n786_), .B2(new_n577_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n828_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n244_), .ZN(new_n835_));
  XOR2_X1   g634(.A(KEYINPUT120), .B(G141gat), .Z(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1344gat));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n305_), .ZN(new_n838_));
  XOR2_X1   g637(.A(KEYINPUT121), .B(G148gat), .Z(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(G1345gat));
  XNOR2_X1  g639(.A(KEYINPUT61), .B(G155gat), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n834_), .B2(new_n576_), .ZN(new_n844_));
  AOI211_X1 g643(.A(KEYINPUT122), .B(new_n577_), .C1(new_n830_), .C2(new_n833_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n842_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT119), .B1(new_n796_), .B2(new_n829_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n832_), .A2(new_n831_), .A3(new_n828_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n576_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT122), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n834_), .A2(new_n843_), .A3(new_n576_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n851_), .A3(new_n841_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n846_), .A2(new_n852_), .ZN(G1346gat));
  INV_X1    g652(.A(G162gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n834_), .A2(new_n854_), .A3(new_n561_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n618_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n854_), .ZN(G1347gat));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n595_), .A2(new_n525_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n499_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n802_), .A2(new_n244_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(G169gat), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n861_), .B2(G169gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n858_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n861_), .A2(G169gat), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT123), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n868_), .A2(new_n863_), .A3(KEYINPUT62), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n802_), .A2(new_n244_), .A3(new_n453_), .A4(new_n860_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n866_), .A2(new_n869_), .A3(new_n870_), .ZN(G1348gat));
  OR3_X1    g670(.A1(new_n832_), .A2(KEYINPUT124), .A3(new_n499_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT124), .B1(new_n832_), .B2(new_n499_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n859_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n686_), .A2(new_n313_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .A4(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n802_), .A2(new_n860_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n313_), .B1(new_n877_), .B2(new_n686_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT125), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n876_), .A2(new_n881_), .A3(new_n878_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1349gat));
  NOR3_X1   g682(.A1(new_n877_), .A2(new_n577_), .A3(new_n457_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n872_), .A2(new_n576_), .A3(new_n874_), .A4(new_n873_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n319_), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n877_), .B2(new_n618_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n561_), .A2(new_n318_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n877_), .B2(new_n888_), .ZN(G1351gat));
  AND4_X1   g688(.A1(new_n580_), .A2(new_n796_), .A3(new_n595_), .A4(new_n827_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n244_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n305_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT63), .ZN(new_n896_));
  INV_X1    g695(.A(G211gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n897_), .A3(KEYINPUT126), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n890_), .A2(new_n576_), .A3(new_n895_), .A4(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(KEYINPUT126), .B1(new_n896_), .B2(new_n897_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1354gat));
  AOI21_X1  g700(.A(G218gat), .B1(new_n890_), .B2(new_n561_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n584_), .A2(G218gat), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT127), .Z(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n890_), .B2(new_n904_), .ZN(G1355gat));
endmodule


